module SRAMTemplate(
  input         clock,
  input         reset,
  output        io_r_req_ready, // @[src/main/scala/utils/SRAMTemplate.scala 70:14]
  input         io_r_req_valid, // @[src/main/scala/utils/SRAMTemplate.scala 70:14]
  input  [8:0]  io_r_req_bits_setIdx, // @[src/main/scala/utils/SRAMTemplate.scala 70:14]
  output [27:0] io_r_resp_data_0_tag, // @[src/main/scala/utils/SRAMTemplate.scala 70:14]
  output [1:0]  io_r_resp_data_0__type, // @[src/main/scala/utils/SRAMTemplate.scala 70:14]
  output [38:0] io_r_resp_data_0_target, // @[src/main/scala/utils/SRAMTemplate.scala 70:14]
  output [2:0]  io_r_resp_data_0_brIdx, // @[src/main/scala/utils/SRAMTemplate.scala 70:14]
  output        io_r_resp_data_0_valid, // @[src/main/scala/utils/SRAMTemplate.scala 70:14]
  input         io_w_req_valid, // @[src/main/scala/utils/SRAMTemplate.scala 70:14]
  input  [8:0]  io_w_req_bits_setIdx, // @[src/main/scala/utils/SRAMTemplate.scala 70:14]
  input  [27:0] io_w_req_bits_data_tag, // @[src/main/scala/utils/SRAMTemplate.scala 70:14]
  input  [1:0]  io_w_req_bits_data__type, // @[src/main/scala/utils/SRAMTemplate.scala 70:14]
  input  [38:0] io_w_req_bits_data_target, // @[src/main/scala/utils/SRAMTemplate.scala 70:14]
  input  [2:0]  io_w_req_bits_data_brIdx // @[src/main/scala/utils/SRAMTemplate.scala 70:14]
);
`ifdef RANDOMIZE_MEM_INIT
  reg [95:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [95:0] _RAND_6;
`endif // RANDOMIZE_REG_INIT
  reg [72:0] array_0 [0:511]; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
  wire  array_0_rdata_MPORT_en; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
  wire [8:0] array_0_rdata_MPORT_addr; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
  wire [72:0] array_0_rdata_MPORT_data; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
  wire [72:0] array_0_MPORT_data; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
  wire [8:0] array_0_MPORT_addr; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
  wire  array_0_MPORT_mask; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
  wire  array_0_MPORT_en; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
  reg  array_0_rdata_MPORT_en_pipe_0;
  reg [8:0] array_0_rdata_MPORT_addr_pipe_0;
  reg  resetState; // @[src/main/scala/utils/SRAMTemplate.scala 80:30]
  reg [8:0] resetSet; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
  wire  wrap_wrap = resetSet == 9'h1ff; // @[src/main/scala/chisel3/util/Counter.scala 73:24]
  wire [8:0] _wrap_value_T_1 = resetSet + 9'h1; // @[src/main/scala/chisel3/util/Counter.scala 77:24]
  wire  resetFinish = resetState & wrap_wrap; // @[src/main/scala/chisel3/util/Counter.scala 118:{16,23} 117:24]
  wire  _GEN_2 = resetFinish ? 1'h0 : resetState; // @[src/main/scala/utils/SRAMTemplate.scala 82:24 80:30 82:38]
  wire  wen = io_w_req_valid | resetState; // @[src/main/scala/utils/SRAMTemplate.scala 88:52]
  wire  _realRen_T = ~wen; // @[src/main/scala/utils/SRAMTemplate.scala 89:41]
  wire [72:0] _wdataword_T = {io_w_req_bits_data_tag,io_w_req_bits_data__type,io_w_req_bits_data_target,
    io_w_req_bits_data_brIdx,1'h1}; // @[src/main/scala/utils/SRAMTemplate.scala 92:78]
  reg  rdata_REG; // @[src/main/scala/utils/Hold.scala 28:106]
  reg [72:0] rdata_r_0; // @[src/main/scala/utils/Hold.scala 23:65]
  wire [72:0] _GEN_14 = rdata_REG ? array_0_rdata_MPORT_data : rdata_r_0; // @[src/main/scala/utils/Hold.scala 23:{65,65,65}]
  assign array_0_rdata_MPORT_en = array_0_rdata_MPORT_en_pipe_0;
  assign array_0_rdata_MPORT_addr = array_0_rdata_MPORT_addr_pipe_0;
  assign array_0_rdata_MPORT_data = array_0[array_0_rdata_MPORT_addr]; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
  assign array_0_MPORT_data = resetState ? 73'h0 : _wdataword_T;
  assign array_0_MPORT_addr = resetState ? resetSet : io_w_req_bits_setIdx;
  assign array_0_MPORT_mask = 1'h1;
  assign array_0_MPORT_en = io_w_req_valid | resetState;
  assign io_r_req_ready = ~resetState & _realRen_T; // @[src/main/scala/utils/SRAMTemplate.scala 101:33]
  assign io_r_resp_data_0_tag = _GEN_14[72:45]; // @[src/main/scala/utils/SRAMTemplate.scala 98:78]
  assign io_r_resp_data_0__type = _GEN_14[44:43]; // @[src/main/scala/utils/SRAMTemplate.scala 98:78]
  assign io_r_resp_data_0_target = _GEN_14[42:4]; // @[src/main/scala/utils/SRAMTemplate.scala 98:78]
  assign io_r_resp_data_0_brIdx = _GEN_14[3:1]; // @[src/main/scala/utils/SRAMTemplate.scala 98:78]
  assign io_r_resp_data_0_valid = _GEN_14[0]; // @[src/main/scala/utils/SRAMTemplate.scala 98:78]
  always @(posedge clock) begin
    if (array_0_MPORT_en & array_0_MPORT_mask) begin
      array_0[array_0_MPORT_addr] <= array_0_MPORT_data; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
    end
    array_0_rdata_MPORT_en_pipe_0 <= io_r_req_valid & _realRen_T;
    if (io_r_req_valid & _realRen_T) begin
      array_0_rdata_MPORT_addr_pipe_0 <= io_r_req_bits_setIdx;
    end
    resetState <= reset | _GEN_2; // @[src/main/scala/utils/SRAMTemplate.scala 80:{30,30}]
    if (reset) begin // @[src/main/scala/chisel3/util/Counter.scala 61:40]
      resetSet <= 9'h0; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end else if (resetState) begin // @[src/main/scala/chisel3/util/Counter.scala 118:16]
      resetSet <= _wrap_value_T_1; // @[src/main/scala/chisel3/util/Counter.scala 77:15]
    end
    rdata_REG <= io_r_req_valid & ~wen; // @[src/main/scala/utils/SRAMTemplate.scala 89:38]
    if (reset) begin // @[src/main/scala/utils/Hold.scala 23:65]
      rdata_r_0 <= 73'h0; // @[src/main/scala/utils/Hold.scala 23:65]
    end else if (rdata_REG) begin // @[src/main/scala/utils/Hold.scala 23:65]
      rdata_r_0 <= array_0_rdata_MPORT_data; // @[src/main/scala/utils/Hold.scala 23:65]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {3{`RANDOM}};
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    array_0[initvar] = _RAND_0[72:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  array_0_rdata_MPORT_en_pipe_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  array_0_rdata_MPORT_addr_pipe_0 = _RAND_2[8:0];
  _RAND_3 = {1{`RANDOM}};
  resetState = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  resetSet = _RAND_4[8:0];
  _RAND_5 = {1{`RANDOM}};
  rdata_REG = _RAND_5[0:0];
  _RAND_6 = {3{`RANDOM}};
  rdata_r_0 = _RAND_6[72:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module BPU_inorder(
  input         clock,
  input         reset,
  input         io_in_pc_valid, // @[src/main/scala/nutcore/frontend/BPU.scala 281:14]
  input  [38:0] io_in_pc_bits, // @[src/main/scala/nutcore/frontend/BPU.scala 281:14]
  output [38:0] io_out_target, // @[src/main/scala/nutcore/frontend/BPU.scala 281:14]
  output        io_out_valid, // @[src/main/scala/nutcore/frontend/BPU.scala 281:14]
  input         io_flush, // @[src/main/scala/nutcore/frontend/BPU.scala 281:14]
  output [2:0]  io_brIdx, // @[src/main/scala/nutcore/frontend/BPU.scala 281:14]
  output        io_crosslineJump, // @[src/main/scala/nutcore/frontend/BPU.scala 281:14]
  input         bpuUpdateReq_valid,
  input  [38:0] bpuUpdateReq_pc,
  input         bpuUpdateReq_isMissPredict,
  input  [38:0] bpuUpdateReq_actualTarget,
  input         bpuUpdateReq_actualTaken,
  input  [6:0]  bpuUpdateReq_fuOpType,
  input  [1:0]  bpuUpdateReq_btbType,
  input         bpuUpdateReq_isRVC,
  input         DISPLAY_ENABLE,
  input         MOUFlushICache,
  input         MOUFlushTLB
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [63:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [63:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
`endif // RANDOMIZE_REG_INIT
  wire  btb_clock; // @[src/main/scala/nutcore/frontend/BPU.scala 302:19]
  wire  btb_reset; // @[src/main/scala/nutcore/frontend/BPU.scala 302:19]
  wire  btb_io_r_req_ready; // @[src/main/scala/nutcore/frontend/BPU.scala 302:19]
  wire  btb_io_r_req_valid; // @[src/main/scala/nutcore/frontend/BPU.scala 302:19]
  wire [8:0] btb_io_r_req_bits_setIdx; // @[src/main/scala/nutcore/frontend/BPU.scala 302:19]
  wire [27:0] btb_io_r_resp_data_0_tag; // @[src/main/scala/nutcore/frontend/BPU.scala 302:19]
  wire [1:0] btb_io_r_resp_data_0__type; // @[src/main/scala/nutcore/frontend/BPU.scala 302:19]
  wire [38:0] btb_io_r_resp_data_0_target; // @[src/main/scala/nutcore/frontend/BPU.scala 302:19]
  wire [2:0] btb_io_r_resp_data_0_brIdx; // @[src/main/scala/nutcore/frontend/BPU.scala 302:19]
  wire  btb_io_r_resp_data_0_valid; // @[src/main/scala/nutcore/frontend/BPU.scala 302:19]
  wire  btb_io_w_req_valid; // @[src/main/scala/nutcore/frontend/BPU.scala 302:19]
  wire [8:0] btb_io_w_req_bits_setIdx; // @[src/main/scala/nutcore/frontend/BPU.scala 302:19]
  wire [27:0] btb_io_w_req_bits_data_tag; // @[src/main/scala/nutcore/frontend/BPU.scala 302:19]
  wire [1:0] btb_io_w_req_bits_data__type; // @[src/main/scala/nutcore/frontend/BPU.scala 302:19]
  wire [38:0] btb_io_w_req_bits_data_target; // @[src/main/scala/nutcore/frontend/BPU.scala 302:19]
  wire [2:0] btb_io_w_req_bits_data_brIdx; // @[src/main/scala/nutcore/frontend/BPU.scala 302:19]
  reg [1:0] pht [0:511]; // @[src/main/scala/nutcore/frontend/BPU.scala 339:16]
  wire  pht_phtTaken_MPORT_en; // @[src/main/scala/nutcore/frontend/BPU.scala 339:16]
  wire [8:0] pht_phtTaken_MPORT_addr; // @[src/main/scala/nutcore/frontend/BPU.scala 339:16]
  wire [1:0] pht_phtTaken_MPORT_data; // @[src/main/scala/nutcore/frontend/BPU.scala 339:16]
  wire  pht_cnt_MPORT_en; // @[src/main/scala/nutcore/frontend/BPU.scala 339:16]
  wire [8:0] pht_cnt_MPORT_addr; // @[src/main/scala/nutcore/frontend/BPU.scala 339:16]
  wire [1:0] pht_cnt_MPORT_data; // @[src/main/scala/nutcore/frontend/BPU.scala 339:16]
  wire [1:0] pht_MPORT_data; // @[src/main/scala/nutcore/frontend/BPU.scala 339:16]
  wire [8:0] pht_MPORT_addr; // @[src/main/scala/nutcore/frontend/BPU.scala 339:16]
  wire  pht_MPORT_mask; // @[src/main/scala/nutcore/frontend/BPU.scala 339:16]
  wire  pht_MPORT_en; // @[src/main/scala/nutcore/frontend/BPU.scala 339:16]
  reg [38:0] ras [0:15]; // @[src/main/scala/nutcore/frontend/BPU.scala 345:16]
  wire  ras_rasTarget_MPORT_en; // @[src/main/scala/nutcore/frontend/BPU.scala 345:16]
  wire [3:0] ras_rasTarget_MPORT_addr; // @[src/main/scala/nutcore/frontend/BPU.scala 345:16]
  wire [38:0] ras_rasTarget_MPORT_data; // @[src/main/scala/nutcore/frontend/BPU.scala 345:16]
  wire [38:0] ras_MPORT_1_data; // @[src/main/scala/nutcore/frontend/BPU.scala 345:16]
  wire [3:0] ras_MPORT_1_addr; // @[src/main/scala/nutcore/frontend/BPU.scala 345:16]
  wire  ras_MPORT_1_mask; // @[src/main/scala/nutcore/frontend/BPU.scala 345:16]
  wire  ras_MPORT_1_en; // @[src/main/scala/nutcore/frontend/BPU.scala 345:16]
  reg  flush; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  _GEN_0 = io_in_pc_valid ? 1'h0 : flush; // @[src/main/scala/utils/StopWatch.scala 26:19 24:20 26:23]
  wire  _GEN_1 = io_flush | _GEN_0; // @[src/main/scala/utils/StopWatch.scala 27:{20,24}]
  wire  _btb_reset_T_2 = reset | (MOUFlushICache | MOUFlushTLB); // @[src/main/scala/nutcore/frontend/BPU.scala 308:29]
  reg [63:0] c; // @[src/main/scala/utils/GTimer.scala 24:20]
  wire [63:0] _c_T_1 = c + 64'h1; // @[src/main/scala/utils/GTimer.scala 25:12]
  wire  _T_3 = _btb_reset_T_2 & DISPLAY_ENABLE; // @[src/main/scala/utils/Debug.scala 55:16]
  wire  _T_5 = ~reset; // @[src/main/scala/utils/Debug.scala 56:24]
  reg [38:0] pcLatch; // @[src/main/scala/nutcore/frontend/BPU.scala 319:26]
  wire [27:0] btbRead_tag = btb_io_r_resp_data_0_tag; // @[src/main/scala/nutcore/frontend/BPU.scala 315:21 316:11]
  wire  btbRead_valid = btb_io_r_resp_data_0_valid; // @[src/main/scala/nutcore/frontend/BPU.scala 315:21 316:11]
  reg  btbHit_REG; // @[src/main/scala/nutcore/frontend/BPU.scala 320:93]
  wire [2:0] btbRead_brIdx = btb_io_r_resp_data_0_brIdx; // @[src/main/scala/nutcore/frontend/BPU.scala 315:21 316:11]
  wire  btbHit = btbRead_valid & btbRead_tag == pcLatch[38:11] & ~flush & btbHit_REG & ~(pcLatch[1] & btbRead_brIdx[0]); // @[src/main/scala/nutcore/frontend/BPU.scala 320:130]
  wire  crosslineJump = btbRead_brIdx[2] & btbHit; // @[src/main/scala/nutcore/frontend/BPU.scala 330:40]
  reg [63:0] c_1; // @[src/main/scala/utils/GTimer.scala 24:20]
  wire [63:0] _c_T_3 = c_1 + 64'h1; // @[src/main/scala/utils/GTimer.scala 25:12]
  reg [63:0] c_2; // @[src/main/scala/utils/GTimer.scala 24:20]
  wire [63:0] _c_T_5 = c_2 + 64'h1; // @[src/main/scala/utils/GTimer.scala 25:12]
  wire  _T_14 = btbHit & DISPLAY_ENABLE; // @[src/main/scala/utils/Debug.scala 55:16]
  wire [1:0] _T_20 = io_out_valid ? 2'h3 : 2'h0; // @[src/main/scala/nutcore/frontend/BPU.scala 335:94]
  wire [2:0] _T_21 = {crosslineJump,_T_20}; // @[src/main/scala/nutcore/frontend/BPU.scala 335:74]
  reg [63:0] c_3; // @[src/main/scala/utils/GTimer.scala 24:20]
  wire [63:0] _c_T_7 = c_3 + 64'h1; // @[src/main/scala/utils/GTimer.scala 25:12]
  reg  phtTaken; // @[src/main/scala/nutcore/frontend/BPU.scala 340:27]
  reg [3:0] sp_value; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
  reg [38:0] rasTarget; // @[src/main/scala/nutcore/frontend/BPU.scala 348:28]
  wire  _T_35 = ~bpuUpdateReq_pc[1]; // @[src/main/scala/nutcore/frontend/BPU.scala 356:150]
  wire [1:0] _T_36 = {bpuUpdateReq_pc[1],_T_35}; // @[src/main/scala/nutcore/frontend/BPU.scala 356:138]
  reg [63:0] c_4; // @[src/main/scala/utils/GTimer.scala 24:20]
  wire [63:0] _c_T_9 = c_4 + 64'h1; // @[src/main/scala/utils/GTimer.scala 25:12]
  wire  _T_37 = bpuUpdateReq_valid & DISPLAY_ENABLE; // @[src/main/scala/utils/Debug.scala 55:16]
  wire  _btbWrite_brIdx_T_3 = bpuUpdateReq_pc[2:0] == 3'h6 & ~bpuUpdateReq_isRVC; // @[src/main/scala/nutcore/frontend/BPU.scala 370:46]
  wire [1:0] btbWrite_brIdx_hi = {_btbWrite_brIdx_T_3,bpuUpdateReq_pc[1]}; // @[src/main/scala/nutcore/frontend/BPU.scala 370:24]
  reg [1:0] cnt; // @[src/main/scala/nutcore/frontend/BPU.scala 392:20]
  reg  reqLatch_valid; // @[src/main/scala/nutcore/frontend/BPU.scala 393:25]
  reg [38:0] reqLatch_pc; // @[src/main/scala/nutcore/frontend/BPU.scala 393:25]
  reg  reqLatch_actualTaken; // @[src/main/scala/nutcore/frontend/BPU.scala 393:25]
  reg [6:0] reqLatch_fuOpType; // @[src/main/scala/nutcore/frontend/BPU.scala 393:25]
  wire  _T_43 = ~reqLatch_fuOpType[3]; // @[src/main/scala/nutcore/backend/fu/ALU.scala 63:30]
  wire  _T_44 = reqLatch_valid & _T_43; // @[src/main/scala/nutcore/frontend/BPU.scala 394:24]
  wire [1:0] _newCnt_T_1 = cnt + 2'h1; // @[src/main/scala/nutcore/frontend/BPU.scala 396:33]
  wire [1:0] _newCnt_T_3 = cnt - 2'h1; // @[src/main/scala/nutcore/frontend/BPU.scala 396:44]
  wire  wen = reqLatch_actualTaken & cnt != 2'h3 | ~reqLatch_actualTaken & cnt != 2'h0; // @[src/main/scala/nutcore/frontend/BPU.scala 397:44]
  wire  _T_48 = bpuUpdateReq_fuOpType == 7'h5c; // @[src/main/scala/nutcore/frontend/BPU.scala 406:24]
  wire [3:0] _T_50 = sp_value + 4'h1; // @[src/main/scala/nutcore/frontend/BPU.scala 407:26]
  wire [38:0] _T_52 = bpuUpdateReq_pc + 39'h2; // @[src/main/scala/nutcore/frontend/BPU.scala 407:55]
  wire [38:0] _T_54 = bpuUpdateReq_pc + 39'h4; // @[src/main/scala/nutcore/frontend/BPU.scala 407:69]
  wire  _T_57 = sp_value == 4'h0; // @[src/main/scala/nutcore/frontend/BPU.scala 412:21]
  wire [3:0] _value_T_4 = sp_value - 4'h1; // @[src/main/scala/nutcore/frontend/BPU.scala 415:53]
  wire [3:0] _value_T_5 = _T_57 ? 4'h0 : _value_T_4; // @[src/main/scala/nutcore/frontend/BPU.scala 415:22]
  wire [1:0] btbRead__type = btb_io_r_resp_data_0__type; // @[src/main/scala/nutcore/frontend/BPU.scala 315:21 316:11]
  wire [38:0] btbRead_target = btb_io_r_resp_data_0_target; // @[src/main/scala/nutcore/frontend/BPU.scala 315:21 316:11]
  wire [3:0] _io_brIdx_T_2 = {1'h1,crosslineJump,_T_20}; // @[src/main/scala/nutcore/frontend/BPU.scala 422:35]
  wire [3:0] _GEN_28 = {{1'd0}, btbRead_brIdx}; // @[src/main/scala/nutcore/frontend/BPU.scala 422:30]
  wire [3:0] _io_brIdx_T_3 = _GEN_28 & _io_brIdx_T_2; // @[src/main/scala/nutcore/frontend/BPU.scala 422:30]
  wire  _io_out_valid_T_3 = btbRead__type == 2'h0 ? phtTaken : rasTarget != 39'h0; // @[src/main/scala/nutcore/frontend/BPU.scala 423:32]
  SRAMTemplate btb ( // @[src/main/scala/nutcore/frontend/BPU.scala 302:19]
    .clock(btb_clock),
    .reset(btb_reset),
    .io_r_req_ready(btb_io_r_req_ready),
    .io_r_req_valid(btb_io_r_req_valid),
    .io_r_req_bits_setIdx(btb_io_r_req_bits_setIdx),
    .io_r_resp_data_0_tag(btb_io_r_resp_data_0_tag),
    .io_r_resp_data_0__type(btb_io_r_resp_data_0__type),
    .io_r_resp_data_0_target(btb_io_r_resp_data_0_target),
    .io_r_resp_data_0_brIdx(btb_io_r_resp_data_0_brIdx),
    .io_r_resp_data_0_valid(btb_io_r_resp_data_0_valid),
    .io_w_req_valid(btb_io_w_req_valid),
    .io_w_req_bits_setIdx(btb_io_w_req_bits_setIdx),
    .io_w_req_bits_data_tag(btb_io_w_req_bits_data_tag),
    .io_w_req_bits_data__type(btb_io_w_req_bits_data__type),
    .io_w_req_bits_data_target(btb_io_w_req_bits_data_target),
    .io_w_req_bits_data_brIdx(btb_io_w_req_bits_data_brIdx)
  );
  assign pht_phtTaken_MPORT_en = 1'h1;
  assign pht_phtTaken_MPORT_addr = io_in_pc_bits[10:2];
  assign pht_phtTaken_MPORT_data = pht[pht_phtTaken_MPORT_addr]; // @[src/main/scala/nutcore/frontend/BPU.scala 339:16]
  assign pht_cnt_MPORT_en = 1'h1;
  assign pht_cnt_MPORT_addr = bpuUpdateReq_pc[10:2];
  assign pht_cnt_MPORT_data = pht[pht_cnt_MPORT_addr]; // @[src/main/scala/nutcore/frontend/BPU.scala 339:16]
  assign pht_MPORT_data = reqLatch_actualTaken ? _newCnt_T_1 : _newCnt_T_3;
  assign pht_MPORT_addr = reqLatch_pc[10:2];
  assign pht_MPORT_mask = 1'h1;
  assign pht_MPORT_en = _T_44 & wen;
  assign ras_rasTarget_MPORT_en = 1'h1;
  assign ras_rasTarget_MPORT_addr = sp_value;
  assign ras_rasTarget_MPORT_data = ras[ras_rasTarget_MPORT_addr]; // @[src/main/scala/nutcore/frontend/BPU.scala 345:16]
  assign ras_MPORT_1_data = bpuUpdateReq_isRVC ? _T_52 : _T_54;
  assign ras_MPORT_1_addr = sp_value + 4'h1;
  assign ras_MPORT_1_mask = 1'h1;
  assign ras_MPORT_1_en = bpuUpdateReq_valid & _T_48;
  assign io_out_target = btbRead__type == 2'h3 ? rasTarget : btbRead_target; // @[src/main/scala/nutcore/frontend/BPU.scala 419:23]
  assign io_out_valid = btbHit & _io_out_valid_T_3; // @[src/main/scala/nutcore/frontend/BPU.scala 423:26]
  assign io_brIdx = _io_brIdx_T_3[2:0]; // @[src/main/scala/nutcore/frontend/BPU.scala 422:13]
  assign io_crosslineJump = btbRead_brIdx[2] & btbHit; // @[src/main/scala/nutcore/frontend/BPU.scala 330:40]
  assign btb_clock = clock;
  assign btb_reset = reset | (MOUFlushICache | MOUFlushTLB); // @[src/main/scala/nutcore/frontend/BPU.scala 308:29]
  assign btb_io_r_req_valid = io_in_pc_valid; // @[src/main/scala/nutcore/frontend/BPU.scala 311:22]
  assign btb_io_r_req_bits_setIdx = io_in_pc_bits[10:2]; // @[src/main/scala/nutcore/frontend/BPU.scala 35:65]
  assign btb_io_w_req_valid = bpuUpdateReq_isMissPredict & bpuUpdateReq_valid; // @[src/main/scala/nutcore/frontend/BPU.scala 378:43]
  assign btb_io_w_req_bits_setIdx = bpuUpdateReq_pc[10:2]; // @[src/main/scala/nutcore/frontend/BPU.scala 35:65]
  assign btb_io_w_req_bits_data_tag = bpuUpdateReq_pc[38:11]; // @[src/main/scala/nutcore/frontend/BPU.scala 35:65]
  assign btb_io_w_req_bits_data__type = bpuUpdateReq_btbType; // @[src/main/scala/nutcore/frontend/BPU.scala 352:21]
  assign btb_io_w_req_bits_data_target = bpuUpdateReq_actualTarget; // @[src/main/scala/nutcore/frontend/BPU.scala 352:21]
  assign btb_io_w_req_bits_data_brIdx = {btbWrite_brIdx_hi,_T_35}; // @[src/main/scala/nutcore/frontend/BPU.scala 370:24]
  always @(posedge clock) begin
    if (pht_MPORT_en & pht_MPORT_mask) begin
      pht[pht_MPORT_addr] <= pht_MPORT_data; // @[src/main/scala/nutcore/frontend/BPU.scala 339:16]
    end
    if (ras_MPORT_1_en & ras_MPORT_1_mask) begin
      ras[ras_MPORT_1_addr] <= ras_MPORT_1_data; // @[src/main/scala/nutcore/frontend/BPU.scala 345:16]
    end
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      flush <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else begin
      flush <= _GEN_1;
    end
    if (reset) begin // @[src/main/scala/utils/GTimer.scala 24:20]
      c <= 64'h0; // @[src/main/scala/utils/GTimer.scala 24:20]
    end else begin
      c <= _c_T_1; // @[src/main/scala/utils/GTimer.scala 25:7]
    end
    if (io_in_pc_valid) begin // @[src/main/scala/nutcore/frontend/BPU.scala 319:26]
      pcLatch <= io_in_pc_bits; // @[src/main/scala/nutcore/frontend/BPU.scala 319:26]
    end
    if (reset) begin // @[src/main/scala/nutcore/frontend/BPU.scala 320:93]
      btbHit_REG <= 1'h0; // @[src/main/scala/nutcore/frontend/BPU.scala 320:93]
    end else begin
      btbHit_REG <= btb_io_r_req_ready; // @[src/main/scala/nutcore/frontend/BPU.scala 320:93]
    end
    if (reset) begin // @[src/main/scala/utils/GTimer.scala 24:20]
      c_1 <= 64'h0; // @[src/main/scala/utils/GTimer.scala 24:20]
    end else begin
      c_1 <= _c_T_3; // @[src/main/scala/utils/GTimer.scala 25:7]
    end
    if (reset) begin // @[src/main/scala/utils/GTimer.scala 24:20]
      c_2 <= 64'h0; // @[src/main/scala/utils/GTimer.scala 24:20]
    end else begin
      c_2 <= _c_T_5; // @[src/main/scala/utils/GTimer.scala 25:7]
    end
    if (reset) begin // @[src/main/scala/utils/GTimer.scala 24:20]
      c_3 <= 64'h0; // @[src/main/scala/utils/GTimer.scala 24:20]
    end else begin
      c_3 <= _c_T_7; // @[src/main/scala/utils/GTimer.scala 25:7]
    end
    if (io_in_pc_valid) begin // @[src/main/scala/nutcore/frontend/BPU.scala 340:27]
      phtTaken <= pht_phtTaken_MPORT_data[1]; // @[src/main/scala/nutcore/frontend/BPU.scala 340:27]
    end
    if (reset) begin // @[src/main/scala/chisel3/util/Counter.scala 61:40]
      sp_value <= 4'h0; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end else if (bpuUpdateReq_valid) begin // @[src/main/scala/nutcore/frontend/BPU.scala 405:20]
      if (bpuUpdateReq_fuOpType == 7'h5c) begin // @[src/main/scala/nutcore/frontend/BPU.scala 406:45]
        sp_value <= _T_50; // @[src/main/scala/nutcore/frontend/BPU.scala 409:16]
      end else if (bpuUpdateReq_fuOpType == 7'h5e) begin // @[src/main/scala/nutcore/frontend/BPU.scala 411:48]
        sp_value <= _value_T_5; // @[src/main/scala/nutcore/frontend/BPU.scala 415:16]
      end
    end
    if (io_in_pc_valid) begin // @[src/main/scala/nutcore/frontend/BPU.scala 348:28]
      rasTarget <= ras_rasTarget_MPORT_data; // @[src/main/scala/nutcore/frontend/BPU.scala 348:28]
    end
    if (reset) begin // @[src/main/scala/utils/GTimer.scala 24:20]
      c_4 <= 64'h0; // @[src/main/scala/utils/GTimer.scala 24:20]
    end else begin
      c_4 <= _c_T_9; // @[src/main/scala/utils/GTimer.scala 25:7]
    end
    cnt <= pht_cnt_MPORT_data; // @[src/main/scala/nutcore/frontend/BPU.scala 392:20]
    reqLatch_valid <= bpuUpdateReq_valid; // @[src/main/scala/nutcore/frontend/BPU.scala 352:21]
    reqLatch_pc <= bpuUpdateReq_pc; // @[src/main/scala/nutcore/frontend/BPU.scala 352:21]
    reqLatch_actualTaken <= bpuUpdateReq_actualTaken; // @[src/main/scala/nutcore/frontend/BPU.scala 352:21]
    reqLatch_fuOpType <= bpuUpdateReq_fuOpType; // @[src/main/scala/nutcore/frontend/BPU.scala 352:21]
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3 & ~reset) begin
          $fwrite(32'h80000002,"[%d] BPU_inorder: ",c); // @[src/main/scala/utils/Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3 & _T_5) begin
          $fwrite(32'h80000002,"[BPU-RESET] bpu-reset flushBTB:%d flushTLB:%d\n",MOUFlushICache,MOUFlushTLB); // @[src/main/scala/utils/Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_14 & ~reset) begin
          $fwrite(32'h80000002,"[%d] BPU_inorder: ",c_2); // @[src/main/scala/utils/Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_14 & _T_5) begin
          $fwrite(32'h80000002,"[BTBHT1] %d pc=%x tag=%x,%x index=%x bridx=%x tgt=%x,%x flush %x type:%x\n",c_1,pcLatch,
            btbRead_tag,pcLatch[38:11],pcLatch[10:2],btbRead_brIdx,btbRead_target,io_out_target,flush,btbRead__type); // @[src/main/scala/utils/Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_14 & ~reset) begin
          $fwrite(32'h80000002,"[%d] BPU_inorder: ",c_3); // @[src/main/scala/utils/Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_14 & _T_5) begin
          $fwrite(32'h80000002,"[BTBHT2] btbRead.brIdx %x mask %x\n",btbRead_brIdx,_T_21); // @[src/main/scala/utils/Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_37 & ~reset) begin
          $fwrite(32'h80000002,"[%d] BPU_inorder: ",c_4); // @[src/main/scala/utils/Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_37 & _T_5) begin
          $fwrite(32'h80000002,"[BTBUP] pc=%x tag=%x index=%x bridx=%x tgt=%x type=%x\n",bpuUpdateReq_pc,bpuUpdateReq_pc
            [38:11],bpuUpdateReq_pc[10:2],_T_36,bpuUpdateReq_actualTarget,bpuUpdateReq_btbType); // @[src/main/scala/utils/Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    pht[initvar] = _RAND_0[1:0];
  _RAND_1 = {2{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    ras[initvar] = _RAND_1[38:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  flush = _RAND_2[0:0];
  _RAND_3 = {2{`RANDOM}};
  c = _RAND_3[63:0];
  _RAND_4 = {2{`RANDOM}};
  pcLatch = _RAND_4[38:0];
  _RAND_5 = {1{`RANDOM}};
  btbHit_REG = _RAND_5[0:0];
  _RAND_6 = {2{`RANDOM}};
  c_1 = _RAND_6[63:0];
  _RAND_7 = {2{`RANDOM}};
  c_2 = _RAND_7[63:0];
  _RAND_8 = {2{`RANDOM}};
  c_3 = _RAND_8[63:0];
  _RAND_9 = {1{`RANDOM}};
  phtTaken = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  sp_value = _RAND_10[3:0];
  _RAND_11 = {2{`RANDOM}};
  rasTarget = _RAND_11[38:0];
  _RAND_12 = {2{`RANDOM}};
  c_4 = _RAND_12[63:0];
  _RAND_13 = {1{`RANDOM}};
  cnt = _RAND_13[1:0];
  _RAND_14 = {1{`RANDOM}};
  reqLatch_valid = _RAND_14[0:0];
  _RAND_15 = {2{`RANDOM}};
  reqLatch_pc = _RAND_15[38:0];
  _RAND_16 = {1{`RANDOM}};
  reqLatch_actualTaken = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  reqLatch_fuOpType = _RAND_17[6:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module IFU_inorder(
  input         clock,
  input         reset,
  input         io_imem_req_ready, // @[src/main/scala/nutcore/frontend/IFU.scala 310:14]
  output        io_imem_req_valid, // @[src/main/scala/nutcore/frontend/IFU.scala 310:14]
  output [38:0] io_imem_req_bits_addr, // @[src/main/scala/nutcore/frontend/IFU.scala 310:14]
  output [81:0] io_imem_req_bits_user, // @[src/main/scala/nutcore/frontend/IFU.scala 310:14]
  output        io_imem_resp_ready, // @[src/main/scala/nutcore/frontend/IFU.scala 310:14]
  input         io_imem_resp_valid, // @[src/main/scala/nutcore/frontend/IFU.scala 310:14]
  input  [63:0] io_imem_resp_bits_rdata, // @[src/main/scala/nutcore/frontend/IFU.scala 310:14]
  input  [81:0] io_imem_resp_bits_user, // @[src/main/scala/nutcore/frontend/IFU.scala 310:14]
  input         io_out_ready, // @[src/main/scala/nutcore/frontend/IFU.scala 310:14]
  output        io_out_valid, // @[src/main/scala/nutcore/frontend/IFU.scala 310:14]
  output [63:0] io_out_bits_instr, // @[src/main/scala/nutcore/frontend/IFU.scala 310:14]
  output [38:0] io_out_bits_pc, // @[src/main/scala/nutcore/frontend/IFU.scala 310:14]
  output [38:0] io_out_bits_pnpc, // @[src/main/scala/nutcore/frontend/IFU.scala 310:14]
  output        io_out_bits_exceptionVec_12, // @[src/main/scala/nutcore/frontend/IFU.scala 310:14]
  output [3:0]  io_out_bits_brIdx, // @[src/main/scala/nutcore/frontend/IFU.scala 310:14]
  input  [38:0] io_redirect_target, // @[src/main/scala/nutcore/frontend/IFU.scala 310:14]
  input         io_redirect_valid, // @[src/main/scala/nutcore/frontend/IFU.scala 310:14]
  output [3:0]  io_flushVec, // @[src/main/scala/nutcore/frontend/IFU.scala 310:14]
  input         io_ipf, // @[src/main/scala/nutcore/frontend/IFU.scala 310:14]
  input         REG_valid,
  input  [38:0] REG_pc,
  input         REG_isMissPredict,
  input  [38:0] REG_actualTarget,
  input         REG_actualTaken,
  input  [6:0]  REG_fuOpType,
  input  [1:0]  REG_btbType,
  input         REG_isRVC,
  input         DISPLAY_ENABLE,
  output        _WIRE_7,
  input         _WIRE_11,
  input         _WIRE_1_4,
  output        r_2
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [31:0] _RAND_6;
`endif // RANDOMIZE_REG_INIT
  wire  bp1_clock; // @[src/main/scala/nutcore/frontend/IFU.scala 326:19]
  wire  bp1_reset; // @[src/main/scala/nutcore/frontend/IFU.scala 326:19]
  wire  bp1_io_in_pc_valid; // @[src/main/scala/nutcore/frontend/IFU.scala 326:19]
  wire [38:0] bp1_io_in_pc_bits; // @[src/main/scala/nutcore/frontend/IFU.scala 326:19]
  wire [38:0] bp1_io_out_target; // @[src/main/scala/nutcore/frontend/IFU.scala 326:19]
  wire  bp1_io_out_valid; // @[src/main/scala/nutcore/frontend/IFU.scala 326:19]
  wire  bp1_io_flush; // @[src/main/scala/nutcore/frontend/IFU.scala 326:19]
  wire [2:0] bp1_io_brIdx; // @[src/main/scala/nutcore/frontend/IFU.scala 326:19]
  wire  bp1_io_crosslineJump; // @[src/main/scala/nutcore/frontend/IFU.scala 326:19]
  wire  bp1_bpuUpdateReq_valid; // @[src/main/scala/nutcore/frontend/IFU.scala 326:19]
  wire [38:0] bp1_bpuUpdateReq_pc; // @[src/main/scala/nutcore/frontend/IFU.scala 326:19]
  wire  bp1_bpuUpdateReq_isMissPredict; // @[src/main/scala/nutcore/frontend/IFU.scala 326:19]
  wire [38:0] bp1_bpuUpdateReq_actualTarget; // @[src/main/scala/nutcore/frontend/IFU.scala 326:19]
  wire  bp1_bpuUpdateReq_actualTaken; // @[src/main/scala/nutcore/frontend/IFU.scala 326:19]
  wire [6:0] bp1_bpuUpdateReq_fuOpType; // @[src/main/scala/nutcore/frontend/IFU.scala 326:19]
  wire [1:0] bp1_bpuUpdateReq_btbType; // @[src/main/scala/nutcore/frontend/IFU.scala 326:19]
  wire  bp1_bpuUpdateReq_isRVC; // @[src/main/scala/nutcore/frontend/IFU.scala 326:19]
  wire  bp1_DISPLAY_ENABLE; // @[src/main/scala/nutcore/frontend/IFU.scala 326:19]
  wire  bp1_MOUFlushICache; // @[src/main/scala/nutcore/frontend/IFU.scala 326:19]
  wire  bp1_MOUFlushTLB; // @[src/main/scala/nutcore/frontend/IFU.scala 326:19]
  reg [38:0] pc; // @[src/main/scala/nutcore/frontend/IFU.scala 322:19]
  wire  _pcUpdate_T = io_imem_req_ready & io_imem_req_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  wire  pcUpdate = io_redirect_valid | _pcUpdate_T; // @[src/main/scala/nutcore/frontend/IFU.scala 323:36]
  wire [38:0] _snpc_T_2 = pc + 39'h2; // @[src/main/scala/nutcore/frontend/IFU.scala 324:28]
  wire [38:0] _snpc_T_4 = pc + 39'h4; // @[src/main/scala/nutcore/frontend/IFU.scala 324:38]
  wire [38:0] snpc = pc[1] ? _snpc_T_2 : _snpc_T_4; // @[src/main/scala/nutcore/frontend/IFU.scala 324:17]
  reg  crosslineJumpLatch; // @[src/main/scala/nutcore/frontend/IFU.scala 329:35]
  reg [38:0] crosslineJumpTarget; // @[src/main/scala/nutcore/frontend/IFU.scala 333:38]
  wire [38:0] pnpc = bp1_io_crosslineJump ? snpc : bp1_io_out_target; // @[src/main/scala/nutcore/frontend/IFU.scala 338:17]
  wire [38:0] _npc_T = bp1_io_out_valid ? pnpc : snpc; // @[src/main/scala/nutcore/frontend/IFU.scala 340:104]
  wire [38:0] _npc_T_1 = crosslineJumpLatch ? crosslineJumpTarget : _npc_T; // @[src/main/scala/nutcore/frontend/IFU.scala 340:59]
  wire [38:0] npc = io_redirect_valid ? io_redirect_target : _npc_T_1; // @[src/main/scala/nutcore/frontend/IFU.scala 340:16]
  wire  _npcIsSeq_T = bp1_io_out_valid ? 1'h0 : 1'h1; // @[src/main/scala/nutcore/frontend/IFU.scala 341:114]
  wire  _npcIsSeq_T_2 = crosslineJumpLatch ? 1'h0 : bp1_io_crosslineJump | _npcIsSeq_T; // @[src/main/scala/nutcore/frontend/IFU.scala 341:54]
  wire  npcIsSeq = io_redirect_valid ? 1'h0 : _npcIsSeq_T_2; // @[src/main/scala/nutcore/frontend/IFU.scala 341:21]
  wire [2:0] _brIdx_T = io_redirect_valid ? 3'h0 : bp1_io_brIdx; // @[src/main/scala/nutcore/frontend/IFU.scala 349:29]
  wire [3:0] brIdx = {npcIsSeq,_brIdx_T}; // @[src/main/scala/nutcore/frontend/IFU.scala 349:15]
  reg [63:0] c; // @[src/main/scala/utils/GTimer.scala 24:20]
  wire [63:0] _c_T_1 = c + 64'h1; // @[src/main/scala/utils/GTimer.scala 25:12]
  wire  _T_1 = pcUpdate & DISPLAY_ENABLE; // @[src/main/scala/utils/Debug.scala 55:16]
  wire  _T_3 = ~reset; // @[src/main/scala/utils/Debug.scala 56:24]
  wire [42:0] x6_hi = {npcIsSeq,_brIdx_T,npc}; // @[src/main/scala/nutcore/frontend/IFU.scala 371:82]
  reg [63:0] c_1; // @[src/main/scala/utils/GTimer.scala 24:20]
  wire [63:0] _c_T_3 = c_1 + 64'h1; // @[src/main/scala/utils/GTimer.scala 25:12]
  wire  _T_7 = _pcUpdate_T & DISPLAY_ENABLE; // @[src/main/scala/utils/Debug.scala 55:16]
  wire  _T_12 = io_out_ready & io_out_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  reg [63:0] c_2; // @[src/main/scala/utils/GTimer.scala 24:20]
  wire [63:0] _c_T_5 = c_2 + 64'h1; // @[src/main/scala/utils/GTimer.scala 25:12]
  wire  _T_13 = _T_12 & DISPLAY_ENABLE; // @[src/main/scala/utils/Debug.scala 55:16]
  wire  _T_18 = io_imem_resp_ready & io_imem_resp_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  reg  r; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  _GEN_3 = io_imem_req_valid | r; // @[src/main/scala/utils/StopWatch.scala 24:20 30:{20,24}]
  wire  _WIRE = |io_flushVec; // @[src/main/scala/nutcore/frontend/IFU.scala 394:46]
  BPU_inorder bp1 ( // @[src/main/scala/nutcore/frontend/IFU.scala 326:19]
    .clock(bp1_clock),
    .reset(bp1_reset),
    .io_in_pc_valid(bp1_io_in_pc_valid),
    .io_in_pc_bits(bp1_io_in_pc_bits),
    .io_out_target(bp1_io_out_target),
    .io_out_valid(bp1_io_out_valid),
    .io_flush(bp1_io_flush),
    .io_brIdx(bp1_io_brIdx),
    .io_crosslineJump(bp1_io_crosslineJump),
    .bpuUpdateReq_valid(bp1_bpuUpdateReq_valid),
    .bpuUpdateReq_pc(bp1_bpuUpdateReq_pc),
    .bpuUpdateReq_isMissPredict(bp1_bpuUpdateReq_isMissPredict),
    .bpuUpdateReq_actualTarget(bp1_bpuUpdateReq_actualTarget),
    .bpuUpdateReq_actualTaken(bp1_bpuUpdateReq_actualTaken),
    .bpuUpdateReq_fuOpType(bp1_bpuUpdateReq_fuOpType),
    .bpuUpdateReq_btbType(bp1_bpuUpdateReq_btbType),
    .bpuUpdateReq_isRVC(bp1_bpuUpdateReq_isRVC),
    .DISPLAY_ENABLE(bp1_DISPLAY_ENABLE),
    .MOUFlushICache(bp1_MOUFlushICache),
    .MOUFlushTLB(bp1_MOUFlushTLB)
  );
  assign io_imem_req_valid = io_out_ready; // @[src/main/scala/nutcore/frontend/IFU.scala 372:21]
  assign io_imem_req_bits_addr = {pc[38:1],1'h0}; // @[src/main/scala/nutcore/frontend/IFU.scala 370:36]
  assign io_imem_req_bits_user = {x6_hi,pc}; // @[src/main/scala/nutcore/frontend/IFU.scala 371:82]
  assign io_imem_resp_ready = io_out_ready | io_flushVec[0]; // @[src/main/scala/nutcore/frontend/IFU.scala 374:38]
  assign io_out_valid = io_imem_resp_valid & ~io_flushVec[0]; // @[src/main/scala/nutcore/frontend/IFU.scala 391:38]
  assign io_out_bits_instr = io_imem_resp_bits_rdata; // @[src/main/scala/nutcore/frontend/IFU.scala 384:21]
  assign io_out_bits_pc = io_imem_resp_bits_user[38:0]; // @[src/main/scala/nutcore/frontend/IFU.scala 386:24]
  assign io_out_bits_pnpc = io_imem_resp_bits_user[77:39]; // @[src/main/scala/nutcore/frontend/IFU.scala 387:26]
  assign io_out_bits_exceptionVec_12 = io_ipf; // @[src/main/scala/nutcore/frontend/IFU.scala 390:44]
  assign io_out_bits_brIdx = io_imem_resp_bits_user[81:78]; // @[src/main/scala/nutcore/frontend/IFU.scala 388:27]
  assign io_flushVec = io_redirect_valid ? 4'hf : 4'h0; // @[src/main/scala/nutcore/frontend/IFU.scala 367:21]
  assign _WIRE_7 = _WIRE;
  assign r_2 = r;
  assign bp1_clock = clock;
  assign bp1_reset = reset;
  assign bp1_io_in_pc_valid = io_imem_req_ready & io_imem_req_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  assign bp1_io_in_pc_bits = io_redirect_valid ? io_redirect_target : _npc_T_1; // @[src/main/scala/nutcore/frontend/IFU.scala 340:16]
  assign bp1_io_flush = io_redirect_valid; // @[src/main/scala/nutcore/frontend/IFU.scala 358:16]
  assign bp1_bpuUpdateReq_valid = REG_valid;
  assign bp1_bpuUpdateReq_pc = REG_pc;
  assign bp1_bpuUpdateReq_isMissPredict = REG_isMissPredict;
  assign bp1_bpuUpdateReq_actualTarget = REG_actualTarget;
  assign bp1_bpuUpdateReq_actualTaken = REG_actualTaken;
  assign bp1_bpuUpdateReq_fuOpType = REG_fuOpType;
  assign bp1_bpuUpdateReq_btbType = REG_btbType;
  assign bp1_bpuUpdateReq_isRVC = REG_isRVC;
  assign bp1_DISPLAY_ENABLE = DISPLAY_ENABLE;
  assign bp1_MOUFlushICache = _WIRE_11;
  assign bp1_MOUFlushTLB = _WIRE_1_4;
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/nutcore/frontend/IFU.scala 322:19]
      pc <= 39'h80000000; // @[src/main/scala/nutcore/frontend/IFU.scala 322:19]
    end else if (pcUpdate) begin // @[src/main/scala/nutcore/frontend/IFU.scala 360:19]
      if (io_redirect_valid) begin // @[src/main/scala/nutcore/frontend/IFU.scala 340:16]
        pc <= io_redirect_target;
      end else if (crosslineJumpLatch) begin // @[src/main/scala/nutcore/frontend/IFU.scala 340:59]
        pc <= crosslineJumpTarget;
      end else begin
        pc <= _npc_T;
      end
    end
    if (reset) begin // @[src/main/scala/nutcore/frontend/IFU.scala 329:35]
      crosslineJumpLatch <= 1'h0; // @[src/main/scala/nutcore/frontend/IFU.scala 329:35]
    end else if (pcUpdate | bp1_io_flush) begin // @[src/main/scala/nutcore/frontend/IFU.scala 330:34]
      if (bp1_io_flush) begin // @[src/main/scala/nutcore/frontend/IFU.scala 331:30]
        crosslineJumpLatch <= 1'h0;
      end else begin
        crosslineJumpLatch <= bp1_io_crosslineJump & ~crosslineJumpLatch;
      end
    end
    if (bp1_io_crosslineJump) begin // @[src/main/scala/nutcore/frontend/IFU.scala 333:38]
      crosslineJumpTarget <= bp1_io_out_target; // @[src/main/scala/nutcore/frontend/IFU.scala 333:38]
    end
    if (reset) begin // @[src/main/scala/utils/GTimer.scala 24:20]
      c <= 64'h0; // @[src/main/scala/utils/GTimer.scala 24:20]
    end else begin
      c <= _c_T_1; // @[src/main/scala/utils/GTimer.scala 25:7]
    end
    if (reset) begin // @[src/main/scala/utils/GTimer.scala 24:20]
      c_1 <= 64'h0; // @[src/main/scala/utils/GTimer.scala 24:20]
    end else begin
      c_1 <= _c_T_3; // @[src/main/scala/utils/GTimer.scala 25:7]
    end
    if (reset) begin // @[src/main/scala/utils/GTimer.scala 24:20]
      c_2 <= 64'h0; // @[src/main/scala/utils/GTimer.scala 24:20]
    end else begin
      c_2 <= _c_T_5; // @[src/main/scala/utils/GTimer.scala 25:7]
    end
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      r <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else if (_T_18) begin // @[src/main/scala/utils/StopWatch.scala 31:19]
      r <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 31:23]
    end else begin
      r <= _GEN_3;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1 & ~reset) begin
          $fwrite(32'h80000002,"[%d] IFU_inorder: ",c); // @[src/main/scala/utils/Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1 & _T_3) begin
          $fwrite(32'h80000002,
            "[IFUPC] pc:%x pcUpdate:%d npc:%x RedValid:%d RedTarget:%x LJL:%d LJTarget:%x LJ:%d snpc:%x bpValid:%d pnpn:%x \n"
            ,pc,pcUpdate,npc,io_redirect_valid,io_redirect_target,crosslineJumpLatch,crosslineJumpTarget,
            bp1_io_crosslineJump,snpc,bp1_io_out_valid,pnpc); // @[src/main/scala/utils/Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_7 & ~reset) begin
          $fwrite(32'h80000002,"[%d] IFU_inorder: ",c_1); // @[src/main/scala/utils/Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_7 & _T_3) begin
          $fwrite(32'h80000002,"[IFI] pc=%x user=%x %x %x %x \n",io_imem_req_bits_addr,io_imem_req_bits_user,
            io_redirect_valid,bp1_io_brIdx,brIdx); // @[src/main/scala/utils/Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_13 & ~reset) begin
          $fwrite(32'h80000002,"[%d] IFU_inorder: ",c_2); // @[src/main/scala/utils/Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_13 & _T_3) begin
          $fwrite(32'h80000002,"[IFO] pc=%x inst=%x\n",io_out_bits_pc,io_out_bits_instr); // @[src/main/scala/utils/Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  pc = _RAND_0[38:0];
  _RAND_1 = {1{`RANDOM}};
  crosslineJumpLatch = _RAND_1[0:0];
  _RAND_2 = {2{`RANDOM}};
  crosslineJumpTarget = _RAND_2[38:0];
  _RAND_3 = {2{`RANDOM}};
  c = _RAND_3[63:0];
  _RAND_4 = {2{`RANDOM}};
  c_1 = _RAND_4[63:0];
  _RAND_5 = {2{`RANDOM}};
  c_2 = _RAND_5[63:0];
  _RAND_6 = {1{`RANDOM}};
  r = _RAND_6[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module NaiveRVCAlignBuffer(
  input         clock,
  input         reset,
  output        io_in_ready, // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 27:14]
  input         io_in_valid, // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 27:14]
  input  [63:0] io_in_bits_instr, // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 27:14]
  input  [38:0] io_in_bits_pc, // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 27:14]
  input  [38:0] io_in_bits_pnpc, // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 27:14]
  input         io_in_bits_exceptionVec_12, // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 27:14]
  input  [3:0]  io_in_bits_brIdx, // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 27:14]
  input         io_out_ready, // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 27:14]
  output        io_out_valid, // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 27:14]
  output [63:0] io_out_bits_instr, // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 27:14]
  output [38:0] io_out_bits_pc, // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 27:14]
  output [38:0] io_out_bits_pnpc, // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 27:14]
  output        io_out_bits_exceptionVec_12, // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 27:14]
  output [3:0]  io_out_bits_brIdx, // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 27:14]
  output        io_out_bits_crossPageIPFFix, // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 27:14]
  input         io_flush, // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 27:14]
  input         DISPLAY_ENABLE
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [31:0] _RAND_6;
`endif // RANDOMIZE_REG_INIT
  reg [1:0] state; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 39:22]
  wire  _instr_T = state == 2'h2; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 90:23]
  wire  _instr_T_1 = state == 2'h3; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 90:47]
  wire [79:0] instIn = {16'h0,io_in_bits_instr}; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 42:19]
  reg [15:0] specialInstR; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 66:25]
  wire [31:0] _instr_T_4 = {instIn[15:0],specialInstR}; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 90:73]
  wire  _pcOffset_T = state == 2'h0; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 41:28]
  reg [2:0] pcOffsetR; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 40:26]
  wire [2:0] pcOffset = state == 2'h0 ? io_in_bits_pc[2:0] : pcOffsetR; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 41:21]
  wire  _instr_T_9 = 3'h0 == pcOffset; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [31:0] _instr_T_13 = _instr_T_9 ? instIn[31:0] : 32'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _instr_T_10 = 3'h2 == pcOffset; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [31:0] _instr_T_14 = _instr_T_10 ? instIn[47:16] : 32'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] _instr_T_17 = _instr_T_13 | _instr_T_14; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _instr_T_11 = 3'h4 == pcOffset; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [31:0] _instr_T_15 = _instr_T_11 ? instIn[63:32] : 32'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] _instr_T_18 = _instr_T_17 | _instr_T_15; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _instr_T_12 = 3'h6 == pcOffset; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [31:0] _instr_T_16 = _instr_T_12 ? instIn[79:48] : 32'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] _instr_T_19 = _instr_T_18 | _instr_T_16; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] instr = state == 2'h2 | state == 2'h3 ? _instr_T_4 : _instr_T_19; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 90:15]
  wire  isRVC = instr[1:0] != 2'h3; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 34:26]
  wire  _rvcFinish_T = pcOffset == 3'h0; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 48:28]
  wire  _rvcFinish_T_1 = ~isRVC; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 48:40]
  wire  _rvcFinish_T_5 = pcOffset == 3'h4; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 48:72]
  wire  _rvcFinish_T_11 = pcOffset == 3'h2; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 48:116]
  wire  _rvcFinish_T_16 = pcOffset == 3'h6; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 48:159]
  wire  rvcFinish = pcOffset == 3'h0 & (~isRVC | io_in_bits_brIdx[0]) | pcOffset == 3'h4 & (~isRVC | io_in_bits_brIdx[0]
    ) | pcOffset == 3'h2 & (isRVC | io_in_bits_brIdx[1]) | pcOffset == 3'h6 & isRVC; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 48:147]
  wire  _rvcNext_T_13 = _rvcFinish_T_11 & _rvcFinish_T_1; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 51:122]
  wire  _rvcNext_T_15 = ~io_in_bits_brIdx[1]; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 51:135]
  wire  rvcNext = _rvcFinish_T & (isRVC & ~io_in_bits_brIdx[0]) | _rvcFinish_T_5 & (isRVC & ~io_in_bits_brIdx[0]) |
    _rvcFinish_T_11 & _rvcFinish_T_1 & ~io_in_bits_brIdx[1]; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 51:102]
  wire  _rvcSpecial_T_2 = _rvcFinish_T_16 & _rvcFinish_T_1; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 52:37]
  wire  rvcSpecial = _rvcFinish_T_16 & _rvcFinish_T_1 & ~io_in_bits_brIdx[2]; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 52:47]
  wire  rvcSpecialJump = _rvcSpecial_T_2 & io_in_bits_brIdx[2]; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 53:51]
  wire  pnpcIsSeq = io_in_bits_brIdx[3]; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 54:24]
  wire  _flushIFU_T_2 = _pcOffset_T | state == 2'h1; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 57:36]
  wire  flushIFU = (_pcOffset_T | state == 2'h1) & rvcSpecial & io_in_valid & ~pnpcIsSeq; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 57:87]
  reg [63:0] c; // @[src/main/scala/utils/GTimer.scala 24:20]
  wire [63:0] _c_T_1 = c + 64'h1; // @[src/main/scala/utils/GTimer.scala 25:12]
  wire  _T = flushIFU & DISPLAY_ENABLE; // @[src/main/scala/utils/Debug.scala 55:16]
  wire  _T_2 = ~reset; // @[src/main/scala/utils/Debug.scala 56:24]
  wire  loadNextInstline = _flushIFU_T_2 & (rvcSpecial | rvcSpecialJump) & io_in_valid & pnpcIsSeq; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 60:115]
  reg [38:0] specialPCR; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 64:23]
  reg [38:0] specialNPCR; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 65:24]
  reg  specialIPFR; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 67:28]
  wire  rvcForceLoadNext = _rvcNext_T_13 & io_in_bits_pnpc[2:0] == 3'h4 & _rvcNext_T_15; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 69:86]
  wire  _canGo_T = rvcFinish | rvcNext; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 100:28]
  wire  _canIn_T = rvcFinish | rvcForceLoadNext; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 101:28]
  wire [38:0] _pnpcOut_T_1 = io_in_bits_pc + 39'h2; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 103:76]
  wire [38:0] _pnpcOut_T_3 = io_in_bits_pc + 39'h4; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 103:95]
  wire [38:0] _pnpcOut_T_4 = isRVC ? _pnpcOut_T_1 : _pnpcOut_T_3; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 103:55]
  wire [38:0] _pnpcOut_T_5 = rvcFinish ? io_in_bits_pnpc : _pnpcOut_T_4; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 103:23]
  wire  _T_11 = io_out_ready & io_out_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  wire [1:0] _GEN_0 = _T_11 & rvcFinish ? 2'h0 : state; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 104:{39,46} 39:22]
  wire [2:0] _pcOffsetR_T = isRVC ? 3'h2 : 3'h4; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 107:38]
  wire [2:0] _pcOffsetR_T_2 = pcOffset + _pcOffsetR_T; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 107:33]
  wire [1:0] _GEN_1 = _T_11 & rvcNext ? 2'h1 : _GEN_0; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 105:37 106:17]
  wire [2:0] _GEN_2 = _T_11 & rvcNext ? _pcOffsetR_T_2 : pcOffsetR; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 105:37 107:21 40:26]
  wire [1:0] _GEN_3 = rvcSpecial & io_in_valid ? 2'h2 : _GEN_1; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 109:40 110:17]
  wire [38:0] _pcOut_T_2 = {io_in_bits_pc[38:3],pcOffsetR}; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 126:21]
  wire [38:0] _GEN_27 = 2'h3 == state ? specialPCR : 39'h0; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 161:15 98:18 62:23]
  wire [38:0] _GEN_32 = 2'h2 == state ? specialPCR : _GEN_27; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 149:15 98:18]
  wire [38:0] _GEN_40 = 2'h1 == state ? _pcOut_T_2 : _GEN_32; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 126:15 98:18]
  wire [38:0] pcOut = 2'h0 == state ? io_in_bits_pc : _GEN_40; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 102:15 98:18]
  wire [38:0] _GEN_4 = rvcSpecial & io_in_valid ? pcOut : specialPCR; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 109:40 111:22 64:23]
  wire [15:0] _GEN_5 = rvcSpecial & io_in_valid ? io_in_bits_instr[63:48] : specialInstR; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 109:40 112:24 66:25]
  wire  _GEN_6 = rvcSpecial & io_in_valid ? io_in_bits_exceptionVec_12 : specialIPFR; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 109:40 113:23 67:28]
  wire [1:0] _GEN_7 = rvcSpecialJump & io_in_valid ? 2'h3 : _GEN_3; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 115:44 116:17]
  wire [38:0] _GEN_8 = rvcSpecialJump & io_in_valid ? pcOut : _GEN_4; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 115:44 117:22]
  wire [38:0] _GEN_9 = rvcSpecialJump & io_in_valid ? io_in_bits_pnpc : specialNPCR; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 115:44 118:23 65:24]
  wire [15:0] _GEN_10 = rvcSpecialJump & io_in_valid ? io_in_bits_instr[63:48] : _GEN_5; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 115:44 119:24]
  wire  _GEN_11 = rvcSpecialJump & io_in_valid ? io_in_bits_exceptionVec_12 : _GEN_6; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 115:44 120:23]
  wire [38:0] _pnpcOut_T_7 = pcOut + 39'h2; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 127:68]
  wire [38:0] _pnpcOut_T_9 = pcOut + 39'h4; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 127:79]
  wire [38:0] _pnpcOut_T_10 = isRVC ? _pnpcOut_T_7 : _pnpcOut_T_9; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 127:55]
  wire [38:0] _pnpcOut_T_11 = rvcFinish ? io_in_bits_pnpc : _pnpcOut_T_10; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 127:23]
  wire [38:0] _pnpcOut_T_13 = specialPCR + 39'h4; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 150:31]
  wire [1:0] _GEN_24 = _T_11 ? 2'h1 : state; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 154:26 155:17 39:22]
  wire [2:0] _GEN_25 = _T_11 ? 3'h2 : pcOffsetR; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 154:26 156:21 40:26]
  wire [1:0] _GEN_26 = _T_11 ? 2'h0 : state; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 166:26 167:17 39:22]
  wire [38:0] _GEN_28 = 2'h3 == state ? specialNPCR : 39'h0; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 162:17 98:18 63:25]
  wire  _GEN_29 = 2'h3 == state & io_in_valid; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 164:15 98:18 44:23]
  wire [1:0] _GEN_31 = 2'h3 == state ? _GEN_26 : state; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 98:18 39:22]
  wire [38:0] _GEN_33 = 2'h2 == state ? _pnpcOut_T_13 : _GEN_28; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 150:17 98:18]
  wire  _GEN_34 = 2'h2 == state ? io_in_valid : _GEN_29; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 152:15 98:18]
  wire  _GEN_35 = 2'h2 == state ? 1'h0 : 2'h3 == state; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 153:15 98:18]
  wire [1:0] _GEN_36 = 2'h2 == state ? _GEN_24 : _GEN_31; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 98:18]
  wire [2:0] _GEN_37 = 2'h2 == state ? _GEN_25 : pcOffsetR; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 98:18 40:26]
  wire  _GEN_38 = 2'h1 == state ? _canGo_T : _GEN_34; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 124:15 98:18]
  wire  _GEN_39 = 2'h1 == state ? _canIn_T : _GEN_35; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 125:15 98:18]
  wire [38:0] _GEN_41 = 2'h1 == state ? _pnpcOut_T_11 : _GEN_33; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 127:17 98:18]
  wire  canGo = 2'h0 == state ? rvcFinish | rvcNext : _GEN_38; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 100:15 98:18]
  wire  canIn = 2'h0 == state ? rvcFinish | rvcForceLoadNext : _GEN_39; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 101:15 98:18]
  wire [38:0] pnpcOut = 2'h0 == state ? _pnpcOut_T_5 : _GEN_41; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 103:17 98:18]
  wire  _io_out_bits_brIdx_T_10 = pnpcOut == _pnpcOut_T_9 & _rvcFinish_T_1 | pnpcOut == _pnpcOut_T_7 & isRVC ? 1'h0 : 1'h1
    ; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 185:27]
  wire  _io_out_bits_exceptionVec_12_T_2 = _instr_T_1 | _instr_T; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 191:133]
  assign io_in_ready = ~io_in_valid | _T_11 & canIn | loadNextInstline; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 188:58]
  assign io_out_valid = io_in_valid & canGo; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 187:31]
  assign io_out_bits_instr = {{32'd0}, instr}; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 184:21]
  assign io_out_bits_pc = 2'h0 == state ? io_in_bits_pc : _GEN_40; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 102:15 98:18]
  assign io_out_bits_pnpc = 2'h0 == state ? _pnpcOut_T_5 : _GEN_41; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 103:17 98:18]
  assign io_out_bits_exceptionVec_12 = io_in_bits_exceptionVec_12 | specialIPFR & (_instr_T_1 | _instr_T); // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 191:87]
  assign io_out_bits_brIdx = {{3'd0}, _io_out_bits_brIdx_T_10}; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 185:21]
  assign io_out_bits_crossPageIPFFix = io_in_bits_exceptionVec_12 & _io_out_bits_exceptionVec_12_T_2 & ~specialIPFR; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 192:130]
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 39:22]
      state <= 2'h0; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 39:22]
    end else if (~io_flush) begin // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 97:18]
      if (2'h0 == state) begin // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 98:18]
        state <= _GEN_7;
      end else if (2'h1 == state) begin // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 98:18]
        state <= _GEN_7;
      end else begin
        state <= _GEN_36;
      end
    end else begin
      state <= 2'h0; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 172:11]
    end
    if (~io_flush) begin // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 97:18]
      if (2'h0 == state) begin // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 98:18]
        specialInstR <= _GEN_10;
      end else if (2'h1 == state) begin // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 98:18]
        specialInstR <= _GEN_10;
      end
    end
    if (reset) begin // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 40:26]
      pcOffsetR <= 3'h0; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 40:26]
    end else if (~io_flush) begin // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 97:18]
      if (2'h0 == state) begin // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 98:18]
        pcOffsetR <= _GEN_2;
      end else if (2'h1 == state) begin // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 98:18]
        pcOffsetR <= _GEN_2;
      end else begin
        pcOffsetR <= _GEN_37;
      end
    end
    if (reset) begin // @[src/main/scala/utils/GTimer.scala 24:20]
      c <= 64'h0; // @[src/main/scala/utils/GTimer.scala 24:20]
    end else begin
      c <= _c_T_1; // @[src/main/scala/utils/GTimer.scala 25:7]
    end
    if (~io_flush) begin // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 97:18]
      if (2'h0 == state) begin // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 98:18]
        specialPCR <= _GEN_8;
      end else if (2'h1 == state) begin // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 98:18]
        specialPCR <= _GEN_8;
      end
    end
    if (~io_flush) begin // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 97:18]
      if (2'h0 == state) begin // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 98:18]
        specialNPCR <= _GEN_9;
      end else if (2'h1 == state) begin // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 98:18]
        specialNPCR <= _GEN_9;
      end
    end
    if (reset) begin // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 67:28]
      specialIPFR <= 1'h0; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 67:28]
    end else if (~io_flush) begin // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 97:18]
      if (2'h0 == state) begin // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 98:18]
        specialIPFR <= _GEN_11;
      end else if (2'h1 == state) begin // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 98:18]
        specialIPFR <= _GEN_11;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T & ~reset) begin
          $fwrite(32'h80000002,"[%d] NaiveRVCAlignBuffer: ",c); // @[src/main/scala/utils/Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T & _T_2) begin
          $fwrite(32'h80000002,"flushIFU at pc %x offset %x\n",io_in_bits_pc,pcOffset); // @[src/main/scala/utils/Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2 & ~(~flushIFU)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at NaiveIBF.scala:59 assert(!flushIFU)\n"); // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 59:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~flushIFU) & _T_2) begin
          $fatal; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 59:9]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  specialInstR = _RAND_1[15:0];
  _RAND_2 = {1{`RANDOM}};
  pcOffsetR = _RAND_2[2:0];
  _RAND_3 = {2{`RANDOM}};
  c = _RAND_3[63:0];
  _RAND_4 = {2{`RANDOM}};
  specialPCR = _RAND_4[38:0];
  _RAND_5 = {2{`RANDOM}};
  specialNPCR = _RAND_5[38:0];
  _RAND_6 = {1{`RANDOM}};
  specialIPFR = _RAND_6[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Decoder(
  input         clock,
  input         reset,
  output        io_in_ready, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  input         io_in_valid, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  input  [63:0] io_in_bits_instr, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  input  [38:0] io_in_bits_pc, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  input  [38:0] io_in_bits_pnpc, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  input         io_in_bits_exceptionVec_12, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  input  [3:0]  io_in_bits_brIdx, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  input         io_in_bits_crossPageIPFFix, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  input         io_out_ready, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  output        io_out_valid, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  output [63:0] io_out_bits_cf_instr, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  output [38:0] io_out_bits_cf_pc, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  output [38:0] io_out_bits_cf_pnpc, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  output        io_out_bits_cf_exceptionVec_1, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  output        io_out_bits_cf_exceptionVec_2, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  output        io_out_bits_cf_exceptionVec_12, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  output        io_out_bits_cf_intrVec_0, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  output        io_out_bits_cf_intrVec_1, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  output        io_out_bits_cf_intrVec_2, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  output        io_out_bits_cf_intrVec_3, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  output        io_out_bits_cf_intrVec_4, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  output        io_out_bits_cf_intrVec_5, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  output        io_out_bits_cf_intrVec_6, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  output        io_out_bits_cf_intrVec_7, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  output        io_out_bits_cf_intrVec_8, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  output        io_out_bits_cf_intrVec_9, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  output        io_out_bits_cf_intrVec_10, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  output        io_out_bits_cf_intrVec_11, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  output [3:0]  io_out_bits_cf_brIdx, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  output        io_out_bits_cf_crossPageIPFFix, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  output        io_out_bits_ctrl_src1Type, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  output        io_out_bits_ctrl_src2Type, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  output [2:0]  io_out_bits_ctrl_fuType, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  output [6:0]  io_out_bits_ctrl_fuOpType, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  output [4:0]  io_out_bits_ctrl_rfSrc1, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  output [4:0]  io_out_bits_ctrl_rfSrc2, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  output        io_out_bits_ctrl_rfWen, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  output [4:0]  io_out_bits_ctrl_rfDest, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  output        io_out_bits_ctrl_isNutCoreTrap, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  output [63:0] io_out_bits_data_imm, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  output        io_isWFI, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  input         DISPLAY_ENABLE,
  input  [11:0] intrVecIDU,
  input         DTLBENABLE
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire [63:0] _decodeList_T = io_in_bits_instr & 64'h707f; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_1 = 64'h13 == _decodeList_T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire [63:0] _decodeList_T_2 = io_in_bits_instr & 64'hfc00707f; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_3 = 64'h1013 == _decodeList_T_2; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_5 = 64'h2013 == _decodeList_T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_7 = 64'h3013 == _decodeList_T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_9 = 64'h4013 == _decodeList_T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_11 = 64'h5013 == _decodeList_T_2; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_13 = 64'h6013 == _decodeList_T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_15 = 64'h7013 == _decodeList_T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_17 = 64'h40005013 == _decodeList_T_2; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire [63:0] _decodeList_T_18 = io_in_bits_instr & 64'hfe00707f; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_19 = 64'h33 == _decodeList_T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_21 = 64'h1033 == _decodeList_T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_23 = 64'h2033 == _decodeList_T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_25 = 64'h3033 == _decodeList_T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_27 = 64'h4033 == _decodeList_T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_29 = 64'h5033 == _decodeList_T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_31 = 64'h6033 == _decodeList_T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_33 = 64'h7033 == _decodeList_T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_35 = 64'h40000033 == _decodeList_T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_37 = 64'h40005033 == _decodeList_T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire [63:0] _decodeList_T_38 = io_in_bits_instr & 64'h7f; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_39 = 64'h17 == _decodeList_T_38; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_41 = 64'h37 == _decodeList_T_38; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_43 = 64'h6f == _decodeList_T_38; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_45 = 64'h67 == _decodeList_T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_47 = 64'h63 == _decodeList_T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_49 = 64'h1063 == _decodeList_T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_51 = 64'h4063 == _decodeList_T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_53 = 64'h5063 == _decodeList_T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_55 = 64'h6063 == _decodeList_T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_57 = 64'h7063 == _decodeList_T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_59 = 64'h3 == _decodeList_T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_61 = 64'h1003 == _decodeList_T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_63 = 64'h2003 == _decodeList_T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_65 = 64'h4003 == _decodeList_T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_67 = 64'h5003 == _decodeList_T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_69 = 64'h23 == _decodeList_T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_71 = 64'h1023 == _decodeList_T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_73 = 64'h2023 == _decodeList_T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_75 = 64'h1b == _decodeList_T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_77 = 64'h101b == _decodeList_T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_79 = 64'h501b == _decodeList_T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_81 = 64'h4000501b == _decodeList_T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_83 = 64'h103b == _decodeList_T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_85 = 64'h503b == _decodeList_T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_87 = 64'h4000503b == _decodeList_T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_89 = 64'h3b == _decodeList_T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_91 = 64'h4000003b == _decodeList_T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_93 = 64'h6003 == _decodeList_T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_95 = 64'h3003 == _decodeList_T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_97 = 64'h3023 == _decodeList_T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_99 = 64'h6b == _decodeList_T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_101 = 64'h2000033 == _decodeList_T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_103 = 64'h2001033 == _decodeList_T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_105 = 64'h2002033 == _decodeList_T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_107 = 64'h2003033 == _decodeList_T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_109 = 64'h2004033 == _decodeList_T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_111 = 64'h2005033 == _decodeList_T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_113 = 64'h2006033 == _decodeList_T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_115 = 64'h2007033 == _decodeList_T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_117 = 64'h200003b == _decodeList_T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_119 = 64'h200403b == _decodeList_T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_121 = 64'h200503b == _decodeList_T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_123 = 64'h200603b == _decodeList_T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_125 = 64'h200703b == _decodeList_T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire [63:0] _decodeList_T_126 = io_in_bits_instr & 64'hffffffff; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_127 = 64'h0 == _decodeList_T_126; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire [63:0] _decodeList_T_128 = io_in_bits_instr & 64'he003; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_129 = 64'h0 == _decodeList_T_128; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_131 = 64'h4000 == _decodeList_T_128; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_133 = 64'h6000 == _decodeList_T_128; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_135 = 64'hc000 == _decodeList_T_128; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_137 = 64'he000 == _decodeList_T_128; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire [63:0] _decodeList_T_138 = io_in_bits_instr & 64'hef83; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_139 = 64'h1 == _decodeList_T_138; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_141 = 64'h1 == _decodeList_T_128; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_143 = 64'h2001 == _decodeList_T_128; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_145 = 64'h4001 == _decodeList_T_128; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_147 = 64'h6101 == _decodeList_T_138; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_149 = 64'h6001 == _decodeList_T_128; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire [63:0] _decodeList_T_150 = io_in_bits_instr & 64'hec03; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_151 = 64'h8001 == _decodeList_T_150; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_153 = 64'h8401 == _decodeList_T_150; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_155 = 64'h8801 == _decodeList_T_150; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire [63:0] _decodeList_T_156 = io_in_bits_instr & 64'hfc63; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_157 = 64'h8c01 == _decodeList_T_156; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_159 = 64'h8c21 == _decodeList_T_156; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_161 = 64'h8c41 == _decodeList_T_156; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_163 = 64'h8c61 == _decodeList_T_156; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_165 = 64'h9c01 == _decodeList_T_156; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_167 = 64'h9c21 == _decodeList_T_156; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_169 = 64'ha001 == _decodeList_T_128; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_171 = 64'hc001 == _decodeList_T_128; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_173 = 64'he001 == _decodeList_T_128; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_175 = 64'h2 == _decodeList_T_128; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_177 = 64'h4002 == _decodeList_T_128; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_179 = 64'h6002 == _decodeList_T_128; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire [63:0] _decodeList_T_180 = io_in_bits_instr & 64'hf07f; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_181 = 64'h8002 == _decodeList_T_180; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire [63:0] _decodeList_T_182 = io_in_bits_instr & 64'hf003; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_183 = 64'h8002 == _decodeList_T_182; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire [63:0] _decodeList_T_184 = io_in_bits_instr & 64'hffff; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_185 = 64'h9002 == _decodeList_T_184; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_187 = 64'h9002 == _decodeList_T_180; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_189 = 64'h9002 == _decodeList_T_182; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_191 = 64'hc002 == _decodeList_T_128; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_193 = 64'he002 == _decodeList_T_128; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_195 = 64'h73 == _decodeList_T_126; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_197 = 64'h100073 == _decodeList_T_126; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_199 = 64'h30200073 == _decodeList_T_126; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_201 = 64'hf == _decodeList_T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_203 = 64'h10500073 == _decodeList_T_126; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_205 = 64'h10200073 == _decodeList_T_126; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire [63:0] _decodeList_T_206 = io_in_bits_instr & 64'hfe007fff; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_207 = 64'h12000073 == _decodeList_T_206; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire [63:0] _decodeList_T_208 = io_in_bits_instr & 64'hf9f0707f; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_209 = 64'h1000302f == _decodeList_T_208; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_211 = 64'h1000202f == _decodeList_T_208; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire [63:0] _decodeList_T_212 = io_in_bits_instr & 64'hf800707f; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_213 = 64'h1800302f == _decodeList_T_212; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_215 = 64'h1800202f == _decodeList_T_212; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire [63:0] _decodeList_T_216 = io_in_bits_instr & 64'hf800607f; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_217 = 64'h800202f == _decodeList_T_216; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_219 = 64'h202f == _decodeList_T_216; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_221 = 64'h2000202f == _decodeList_T_216; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_223 = 64'h6000202f == _decodeList_T_216; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_225 = 64'h4000202f == _decodeList_T_216; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_227 = 64'h8000202f == _decodeList_T_216; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_229 = 64'ha000202f == _decodeList_T_216; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_231 = 64'hc000202f == _decodeList_T_216; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_233 = 64'he000202f == _decodeList_T_216; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_235 = 64'h1073 == _decodeList_T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_237 = 64'h2073 == _decodeList_T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_239 = 64'h3073 == _decodeList_T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_241 = 64'h5073 == _decodeList_T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_243 = 64'h6073 == _decodeList_T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_245 = 64'h7073 == _decodeList_T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_247 = 64'h100f == _decodeList_T_126; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire [2:0] _decodeList_T_249 = _decodeList_T_245 ? 3'h4 : {{2'd0}, _decodeList_T_247}; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_250 = _decodeList_T_243 ? 3'h4 : _decodeList_T_249; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_251 = _decodeList_T_241 ? 3'h4 : _decodeList_T_250; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_252 = _decodeList_T_239 ? 3'h4 : _decodeList_T_251; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_253 = _decodeList_T_237 ? 3'h4 : _decodeList_T_252; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_254 = _decodeList_T_235 ? 3'h4 : _decodeList_T_253; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_255 = _decodeList_T_233 ? 3'h5 : _decodeList_T_254; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_256 = _decodeList_T_231 ? 3'h5 : _decodeList_T_255; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_257 = _decodeList_T_229 ? 3'h5 : _decodeList_T_256; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_258 = _decodeList_T_227 ? 3'h5 : _decodeList_T_257; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_259 = _decodeList_T_225 ? 3'h5 : _decodeList_T_258; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_260 = _decodeList_T_223 ? 3'h5 : _decodeList_T_259; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_261 = _decodeList_T_221 ? 3'h5 : _decodeList_T_260; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_262 = _decodeList_T_219 ? 3'h5 : _decodeList_T_261; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_263 = _decodeList_T_217 ? 3'h5 : _decodeList_T_262; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_264 = _decodeList_T_215 ? 4'hf : {{1'd0}, _decodeList_T_263}; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_265 = _decodeList_T_213 ? 4'hf : _decodeList_T_264; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_266 = _decodeList_T_211 ? 4'h4 : _decodeList_T_265; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_267 = _decodeList_T_209 ? 4'h4 : _decodeList_T_266; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_268 = _decodeList_T_207 ? 4'h5 : _decodeList_T_267; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_269 = _decodeList_T_205 ? 4'h4 : _decodeList_T_268; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_270 = _decodeList_T_203 ? 4'h4 : _decodeList_T_269; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_271 = _decodeList_T_201 ? 4'h2 : _decodeList_T_270; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_272 = _decodeList_T_199 ? 4'h4 : _decodeList_T_271; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_273 = _decodeList_T_197 ? 4'h4 : _decodeList_T_272; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_274 = _decodeList_T_195 ? 4'h4 : _decodeList_T_273; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_275 = _decodeList_T_193 ? 4'h2 : _decodeList_T_274; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_276 = _decodeList_T_191 ? 4'h2 : _decodeList_T_275; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_277 = _decodeList_T_189 ? 4'h5 : _decodeList_T_276; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_278 = _decodeList_T_187 ? 4'h4 : _decodeList_T_277; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_279 = _decodeList_T_185 ? 4'h4 : _decodeList_T_278; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_280 = _decodeList_T_183 ? 4'h5 : _decodeList_T_279; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_281 = _decodeList_T_181 ? 4'h4 : _decodeList_T_280; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_282 = _decodeList_T_179 ? 4'h4 : _decodeList_T_281; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_283 = _decodeList_T_177 ? 4'h4 : _decodeList_T_282; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_284 = _decodeList_T_175 ? 4'h4 : _decodeList_T_283; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_285 = _decodeList_T_173 ? 4'h1 : _decodeList_T_284; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_286 = _decodeList_T_171 ? 4'h1 : _decodeList_T_285; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_287 = _decodeList_T_169 ? 4'h7 : _decodeList_T_286; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_288 = _decodeList_T_167 ? 4'h5 : _decodeList_T_287; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_289 = _decodeList_T_165 ? 4'h5 : _decodeList_T_288; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_290 = _decodeList_T_163 ? 4'h5 : _decodeList_T_289; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_291 = _decodeList_T_161 ? 4'h5 : _decodeList_T_290; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_292 = _decodeList_T_159 ? 4'h5 : _decodeList_T_291; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_293 = _decodeList_T_157 ? 4'h5 : _decodeList_T_292; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_294 = _decodeList_T_155 ? 4'h4 : _decodeList_T_293; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_295 = _decodeList_T_153 ? 4'h4 : _decodeList_T_294; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_296 = _decodeList_T_151 ? 4'h4 : _decodeList_T_295; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_297 = _decodeList_T_149 ? 4'h4 : _decodeList_T_296; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_298 = _decodeList_T_147 ? 4'h4 : _decodeList_T_297; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_299 = _decodeList_T_145 ? 4'h4 : _decodeList_T_298; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_300 = _decodeList_T_143 ? 4'h4 : _decodeList_T_299; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_301 = _decodeList_T_141 ? 4'h4 : _decodeList_T_300; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_302 = _decodeList_T_139 ? 4'h4 : _decodeList_T_301; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_303 = _decodeList_T_137 ? 4'h2 : _decodeList_T_302; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_304 = _decodeList_T_135 ? 4'h2 : _decodeList_T_303; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_305 = _decodeList_T_133 ? 4'h4 : _decodeList_T_304; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_306 = _decodeList_T_131 ? 4'h4 : _decodeList_T_305; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_307 = _decodeList_T_129 ? 4'h4 : _decodeList_T_306; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_308 = _decodeList_T_127 ? 4'h0 : _decodeList_T_307; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_309 = _decodeList_T_125 ? 4'h5 : _decodeList_T_308; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_310 = _decodeList_T_123 ? 4'h5 : _decodeList_T_309; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_311 = _decodeList_T_121 ? 4'h5 : _decodeList_T_310; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_312 = _decodeList_T_119 ? 4'h5 : _decodeList_T_311; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_313 = _decodeList_T_117 ? 4'h5 : _decodeList_T_312; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_314 = _decodeList_T_115 ? 4'h5 : _decodeList_T_313; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_315 = _decodeList_T_113 ? 4'h5 : _decodeList_T_314; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_316 = _decodeList_T_111 ? 4'h5 : _decodeList_T_315; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_317 = _decodeList_T_109 ? 4'h5 : _decodeList_T_316; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_318 = _decodeList_T_107 ? 4'h5 : _decodeList_T_317; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_319 = _decodeList_T_105 ? 4'h5 : _decodeList_T_318; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_320 = _decodeList_T_103 ? 4'h5 : _decodeList_T_319; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_321 = _decodeList_T_101 ? 4'h5 : _decodeList_T_320; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_322 = _decodeList_T_99 ? 4'h4 : _decodeList_T_321; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_323 = _decodeList_T_97 ? 4'h2 : _decodeList_T_322; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_324 = _decodeList_T_95 ? 4'h4 : _decodeList_T_323; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_325 = _decodeList_T_93 ? 4'h4 : _decodeList_T_324; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_326 = _decodeList_T_91 ? 4'h5 : _decodeList_T_325; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_327 = _decodeList_T_89 ? 4'h5 : _decodeList_T_326; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_328 = _decodeList_T_87 ? 4'h5 : _decodeList_T_327; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_329 = _decodeList_T_85 ? 4'h5 : _decodeList_T_328; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_330 = _decodeList_T_83 ? 4'h5 : _decodeList_T_329; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_331 = _decodeList_T_81 ? 4'h4 : _decodeList_T_330; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_332 = _decodeList_T_79 ? 4'h4 : _decodeList_T_331; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_333 = _decodeList_T_77 ? 4'h4 : _decodeList_T_332; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_334 = _decodeList_T_75 ? 4'h4 : _decodeList_T_333; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_335 = _decodeList_T_73 ? 4'h2 : _decodeList_T_334; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_336 = _decodeList_T_71 ? 4'h2 : _decodeList_T_335; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_337 = _decodeList_T_69 ? 4'h2 : _decodeList_T_336; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_338 = _decodeList_T_67 ? 4'h4 : _decodeList_T_337; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_339 = _decodeList_T_65 ? 4'h4 : _decodeList_T_338; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_340 = _decodeList_T_63 ? 4'h4 : _decodeList_T_339; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_341 = _decodeList_T_61 ? 4'h4 : _decodeList_T_340; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_342 = _decodeList_T_59 ? 4'h4 : _decodeList_T_341; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_343 = _decodeList_T_57 ? 4'h1 : _decodeList_T_342; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_344 = _decodeList_T_55 ? 4'h1 : _decodeList_T_343; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_345 = _decodeList_T_53 ? 4'h1 : _decodeList_T_344; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_346 = _decodeList_T_51 ? 4'h1 : _decodeList_T_345; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_347 = _decodeList_T_49 ? 4'h1 : _decodeList_T_346; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_348 = _decodeList_T_47 ? 4'h1 : _decodeList_T_347; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_349 = _decodeList_T_45 ? 4'h4 : _decodeList_T_348; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_350 = _decodeList_T_43 ? 4'h7 : _decodeList_T_349; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_351 = _decodeList_T_41 ? 4'h6 : _decodeList_T_350; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_352 = _decodeList_T_39 ? 4'h6 : _decodeList_T_351; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_353 = _decodeList_T_37 ? 4'h5 : _decodeList_T_352; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_354 = _decodeList_T_35 ? 4'h5 : _decodeList_T_353; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_355 = _decodeList_T_33 ? 4'h5 : _decodeList_T_354; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_356 = _decodeList_T_31 ? 4'h5 : _decodeList_T_355; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_357 = _decodeList_T_29 ? 4'h5 : _decodeList_T_356; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_358 = _decodeList_T_27 ? 4'h5 : _decodeList_T_357; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_359 = _decodeList_T_25 ? 4'h5 : _decodeList_T_358; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_360 = _decodeList_T_23 ? 4'h5 : _decodeList_T_359; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_361 = _decodeList_T_21 ? 4'h5 : _decodeList_T_360; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_362 = _decodeList_T_19 ? 4'h5 : _decodeList_T_361; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_363 = _decodeList_T_17 ? 4'h4 : _decodeList_T_362; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_364 = _decodeList_T_15 ? 4'h4 : _decodeList_T_363; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_365 = _decodeList_T_13 ? 4'h4 : _decodeList_T_364; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_366 = _decodeList_T_11 ? 4'h4 : _decodeList_T_365; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_367 = _decodeList_T_9 ? 4'h4 : _decodeList_T_366; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_368 = _decodeList_T_7 ? 4'h4 : _decodeList_T_367; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_369 = _decodeList_T_5 ? 4'h4 : _decodeList_T_368; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_370 = _decodeList_T_3 ? 4'h4 : _decodeList_T_369; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] decodeList_0 = _decodeList_T_1 ? 4'h4 : _decodeList_T_370; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_371 = _decodeList_T_247 ? 3'h4 : 3'h3; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_372 = _decodeList_T_245 ? 3'h3 : _decodeList_T_371; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_373 = _decodeList_T_243 ? 3'h3 : _decodeList_T_372; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_374 = _decodeList_T_241 ? 3'h3 : _decodeList_T_373; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_375 = _decodeList_T_239 ? 3'h3 : _decodeList_T_374; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_376 = _decodeList_T_237 ? 3'h3 : _decodeList_T_375; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_377 = _decodeList_T_235 ? 3'h3 : _decodeList_T_376; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_378 = _decodeList_T_233 ? 3'h1 : _decodeList_T_377; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_379 = _decodeList_T_231 ? 3'h1 : _decodeList_T_378; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_380 = _decodeList_T_229 ? 3'h1 : _decodeList_T_379; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_381 = _decodeList_T_227 ? 3'h1 : _decodeList_T_380; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_382 = _decodeList_T_225 ? 3'h1 : _decodeList_T_381; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_383 = _decodeList_T_223 ? 3'h1 : _decodeList_T_382; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_384 = _decodeList_T_221 ? 3'h1 : _decodeList_T_383; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_385 = _decodeList_T_219 ? 3'h1 : _decodeList_T_384; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_386 = _decodeList_T_217 ? 3'h1 : _decodeList_T_385; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_387 = _decodeList_T_215 ? 3'h1 : _decodeList_T_386; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_388 = _decodeList_T_213 ? 3'h1 : _decodeList_T_387; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_389 = _decodeList_T_211 ? 3'h1 : _decodeList_T_388; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_390 = _decodeList_T_209 ? 3'h1 : _decodeList_T_389; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_391 = _decodeList_T_207 ? 3'h4 : _decodeList_T_390; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_392 = _decodeList_T_205 ? 3'h3 : _decodeList_T_391; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_393 = _decodeList_T_203 ? 3'h0 : _decodeList_T_392; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_394 = _decodeList_T_201 ? 3'h4 : _decodeList_T_393; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_395 = _decodeList_T_199 ? 3'h3 : _decodeList_T_394; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_396 = _decodeList_T_197 ? 3'h3 : _decodeList_T_395; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_397 = _decodeList_T_195 ? 3'h3 : _decodeList_T_396; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_398 = _decodeList_T_193 ? 3'h1 : _decodeList_T_397; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_399 = _decodeList_T_191 ? 3'h1 : _decodeList_T_398; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_400 = _decodeList_T_189 ? 3'h0 : _decodeList_T_399; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_401 = _decodeList_T_187 ? 3'h0 : _decodeList_T_400; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_402 = _decodeList_T_185 ? 3'h3 : _decodeList_T_401; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_403 = _decodeList_T_183 ? 3'h0 : _decodeList_T_402; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_404 = _decodeList_T_181 ? 3'h0 : _decodeList_T_403; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_405 = _decodeList_T_179 ? 3'h1 : _decodeList_T_404; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_406 = _decodeList_T_177 ? 3'h1 : _decodeList_T_405; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_407 = _decodeList_T_175 ? 3'h0 : _decodeList_T_406; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_408 = _decodeList_T_173 ? 3'h0 : _decodeList_T_407; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_409 = _decodeList_T_171 ? 3'h0 : _decodeList_T_408; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_410 = _decodeList_T_169 ? 3'h0 : _decodeList_T_409; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_411 = _decodeList_T_167 ? 3'h0 : _decodeList_T_410; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_412 = _decodeList_T_165 ? 3'h0 : _decodeList_T_411; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_413 = _decodeList_T_163 ? 3'h0 : _decodeList_T_412; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_414 = _decodeList_T_161 ? 3'h0 : _decodeList_T_413; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_415 = _decodeList_T_159 ? 3'h0 : _decodeList_T_414; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_416 = _decodeList_T_157 ? 3'h0 : _decodeList_T_415; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_417 = _decodeList_T_155 ? 3'h0 : _decodeList_T_416; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_418 = _decodeList_T_153 ? 3'h0 : _decodeList_T_417; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_419 = _decodeList_T_151 ? 3'h0 : _decodeList_T_418; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_420 = _decodeList_T_149 ? 3'h0 : _decodeList_T_419; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_421 = _decodeList_T_147 ? 3'h0 : _decodeList_T_420; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_422 = _decodeList_T_145 ? 3'h0 : _decodeList_T_421; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_423 = _decodeList_T_143 ? 3'h0 : _decodeList_T_422; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_424 = _decodeList_T_141 ? 3'h0 : _decodeList_T_423; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_425 = _decodeList_T_139 ? 3'h0 : _decodeList_T_424; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_426 = _decodeList_T_137 ? 3'h1 : _decodeList_T_425; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_427 = _decodeList_T_135 ? 3'h1 : _decodeList_T_426; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_428 = _decodeList_T_133 ? 3'h1 : _decodeList_T_427; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_429 = _decodeList_T_131 ? 3'h1 : _decodeList_T_428; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_430 = _decodeList_T_129 ? 3'h0 : _decodeList_T_429; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_431 = _decodeList_T_127 ? 3'h3 : _decodeList_T_430; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_432 = _decodeList_T_125 ? 3'h2 : _decodeList_T_431; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_433 = _decodeList_T_123 ? 3'h2 : _decodeList_T_432; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_434 = _decodeList_T_121 ? 3'h2 : _decodeList_T_433; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_435 = _decodeList_T_119 ? 3'h2 : _decodeList_T_434; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_436 = _decodeList_T_117 ? 3'h2 : _decodeList_T_435; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_437 = _decodeList_T_115 ? 3'h2 : _decodeList_T_436; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_438 = _decodeList_T_113 ? 3'h2 : _decodeList_T_437; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_439 = _decodeList_T_111 ? 3'h2 : _decodeList_T_438; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_440 = _decodeList_T_109 ? 3'h2 : _decodeList_T_439; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_441 = _decodeList_T_107 ? 3'h2 : _decodeList_T_440; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_442 = _decodeList_T_105 ? 3'h2 : _decodeList_T_441; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_443 = _decodeList_T_103 ? 3'h2 : _decodeList_T_442; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_444 = _decodeList_T_101 ? 3'h2 : _decodeList_T_443; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_445 = _decodeList_T_99 ? 3'h3 : _decodeList_T_444; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_446 = _decodeList_T_97 ? 3'h1 : _decodeList_T_445; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_447 = _decodeList_T_95 ? 3'h1 : _decodeList_T_446; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_448 = _decodeList_T_93 ? 3'h1 : _decodeList_T_447; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_449 = _decodeList_T_91 ? 3'h0 : _decodeList_T_448; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_450 = _decodeList_T_89 ? 3'h0 : _decodeList_T_449; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_451 = _decodeList_T_87 ? 3'h0 : _decodeList_T_450; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_452 = _decodeList_T_85 ? 3'h0 : _decodeList_T_451; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_453 = _decodeList_T_83 ? 3'h0 : _decodeList_T_452; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_454 = _decodeList_T_81 ? 3'h0 : _decodeList_T_453; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_455 = _decodeList_T_79 ? 3'h0 : _decodeList_T_454; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_456 = _decodeList_T_77 ? 3'h0 : _decodeList_T_455; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_457 = _decodeList_T_75 ? 3'h0 : _decodeList_T_456; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_458 = _decodeList_T_73 ? 3'h1 : _decodeList_T_457; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_459 = _decodeList_T_71 ? 3'h1 : _decodeList_T_458; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_460 = _decodeList_T_69 ? 3'h1 : _decodeList_T_459; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_461 = _decodeList_T_67 ? 3'h1 : _decodeList_T_460; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_462 = _decodeList_T_65 ? 3'h1 : _decodeList_T_461; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_463 = _decodeList_T_63 ? 3'h1 : _decodeList_T_462; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_464 = _decodeList_T_61 ? 3'h1 : _decodeList_T_463; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_465 = _decodeList_T_59 ? 3'h1 : _decodeList_T_464; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_466 = _decodeList_T_57 ? 3'h0 : _decodeList_T_465; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_467 = _decodeList_T_55 ? 3'h0 : _decodeList_T_466; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_468 = _decodeList_T_53 ? 3'h0 : _decodeList_T_467; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_469 = _decodeList_T_51 ? 3'h0 : _decodeList_T_468; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_470 = _decodeList_T_49 ? 3'h0 : _decodeList_T_469; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_471 = _decodeList_T_47 ? 3'h0 : _decodeList_T_470; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_472 = _decodeList_T_45 ? 3'h0 : _decodeList_T_471; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_473 = _decodeList_T_43 ? 3'h0 : _decodeList_T_472; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_474 = _decodeList_T_41 ? 3'h0 : _decodeList_T_473; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_475 = _decodeList_T_39 ? 3'h0 : _decodeList_T_474; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_476 = _decodeList_T_37 ? 3'h0 : _decodeList_T_475; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_477 = _decodeList_T_35 ? 3'h0 : _decodeList_T_476; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_478 = _decodeList_T_33 ? 3'h0 : _decodeList_T_477; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_479 = _decodeList_T_31 ? 3'h0 : _decodeList_T_478; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_480 = _decodeList_T_29 ? 3'h0 : _decodeList_T_479; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_481 = _decodeList_T_27 ? 3'h0 : _decodeList_T_480; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_482 = _decodeList_T_25 ? 3'h0 : _decodeList_T_481; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_483 = _decodeList_T_23 ? 3'h0 : _decodeList_T_482; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_484 = _decodeList_T_21 ? 3'h0 : _decodeList_T_483; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_485 = _decodeList_T_19 ? 3'h0 : _decodeList_T_484; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_486 = _decodeList_T_17 ? 3'h0 : _decodeList_T_485; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_487 = _decodeList_T_15 ? 3'h0 : _decodeList_T_486; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_488 = _decodeList_T_13 ? 3'h0 : _decodeList_T_487; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_489 = _decodeList_T_11 ? 3'h0 : _decodeList_T_488; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_490 = _decodeList_T_9 ? 3'h0 : _decodeList_T_489; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_491 = _decodeList_T_7 ? 3'h0 : _decodeList_T_490; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_492 = _decodeList_T_5 ? 3'h0 : _decodeList_T_491; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_493 = _decodeList_T_3 ? 3'h0 : _decodeList_T_492; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] decodeList_1 = _decodeList_T_1 ? 3'h0 : _decodeList_T_493; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_495 = _decodeList_T_245 ? 3'h7 : {{2'd0}, _decodeList_T_247}; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_496 = _decodeList_T_243 ? 3'h6 : _decodeList_T_495; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_497 = _decodeList_T_241 ? 3'h5 : _decodeList_T_496; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_498 = _decodeList_T_239 ? 3'h3 : _decodeList_T_497; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_499 = _decodeList_T_237 ? 3'h2 : _decodeList_T_498; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_500 = _decodeList_T_235 ? 3'h1 : _decodeList_T_499; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [5:0] _decodeList_T_501 = _decodeList_T_233 ? 6'h32 : {{3'd0}, _decodeList_T_500}; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [5:0] _decodeList_T_502 = _decodeList_T_231 ? 6'h31 : _decodeList_T_501; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [5:0] _decodeList_T_503 = _decodeList_T_229 ? 6'h30 : _decodeList_T_502; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [5:0] _decodeList_T_504 = _decodeList_T_227 ? 6'h37 : _decodeList_T_503; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [5:0] _decodeList_T_505 = _decodeList_T_225 ? 6'h26 : _decodeList_T_504; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [5:0] _decodeList_T_506 = _decodeList_T_223 ? 6'h25 : _decodeList_T_505; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [5:0] _decodeList_T_507 = _decodeList_T_221 ? 6'h24 : _decodeList_T_506; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_508 = _decodeList_T_219 ? 7'h63 : {{1'd0}, _decodeList_T_507}; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_509 = _decodeList_T_217 ? 7'h22 : _decodeList_T_508; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_510 = _decodeList_T_215 ? 7'h21 : _decodeList_T_509; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_511 = _decodeList_T_213 ? 7'h21 : _decodeList_T_510; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_512 = _decodeList_T_211 ? 7'h20 : _decodeList_T_511; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_513 = _decodeList_T_209 ? 7'h20 : _decodeList_T_512; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_514 = _decodeList_T_207 ? 7'h2 : _decodeList_T_513; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_515 = _decodeList_T_205 ? 7'h0 : _decodeList_T_514; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_516 = _decodeList_T_203 ? 7'h40 : _decodeList_T_515; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_517 = _decodeList_T_201 ? 7'h0 : _decodeList_T_516; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_518 = _decodeList_T_199 ? 7'h0 : _decodeList_T_517; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_519 = _decodeList_T_197 ? 7'h0 : _decodeList_T_518; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_520 = _decodeList_T_195 ? 7'h0 : _decodeList_T_519; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_521 = _decodeList_T_193 ? 7'hb : _decodeList_T_520; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_522 = _decodeList_T_191 ? 7'ha : _decodeList_T_521; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_523 = _decodeList_T_189 ? 7'h40 : _decodeList_T_522; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_524 = _decodeList_T_187 ? 7'h5a : _decodeList_T_523; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_525 = _decodeList_T_185 ? 7'h0 : _decodeList_T_524; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_526 = _decodeList_T_183 ? 7'h40 : _decodeList_T_525; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_527 = _decodeList_T_181 ? 7'h5a : _decodeList_T_526; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_528 = _decodeList_T_179 ? 7'h3 : _decodeList_T_527; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_529 = _decodeList_T_177 ? 7'h2 : _decodeList_T_528; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_530 = _decodeList_T_175 ? 7'h1 : _decodeList_T_529; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_531 = _decodeList_T_173 ? 7'h11 : _decodeList_T_530; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_532 = _decodeList_T_171 ? 7'h10 : _decodeList_T_531; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_533 = _decodeList_T_169 ? 7'h58 : _decodeList_T_532; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_534 = _decodeList_T_167 ? 7'h60 : _decodeList_T_533; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_535 = _decodeList_T_165 ? 7'h28 : _decodeList_T_534; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_536 = _decodeList_T_163 ? 7'h7 : _decodeList_T_535; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_537 = _decodeList_T_161 ? 7'h6 : _decodeList_T_536; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_538 = _decodeList_T_159 ? 7'h4 : _decodeList_T_537; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_539 = _decodeList_T_157 ? 7'h8 : _decodeList_T_538; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_540 = _decodeList_T_155 ? 7'h7 : _decodeList_T_539; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_541 = _decodeList_T_153 ? 7'hd : _decodeList_T_540; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_542 = _decodeList_T_151 ? 7'h5 : _decodeList_T_541; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_543 = _decodeList_T_149 ? 7'h40 : _decodeList_T_542; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_544 = _decodeList_T_147 ? 7'h40 : _decodeList_T_543; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_545 = _decodeList_T_145 ? 7'h40 : _decodeList_T_544; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_546 = _decodeList_T_143 ? 7'h60 : _decodeList_T_545; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_547 = _decodeList_T_141 ? 7'h40 : _decodeList_T_546; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_548 = _decodeList_T_139 ? 7'h40 : _decodeList_T_547; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_549 = _decodeList_T_137 ? 7'hb : _decodeList_T_548; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_550 = _decodeList_T_135 ? 7'ha : _decodeList_T_549; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_551 = _decodeList_T_133 ? 7'h3 : _decodeList_T_550; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_552 = _decodeList_T_131 ? 7'h2 : _decodeList_T_551; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_553 = _decodeList_T_129 ? 7'h40 : _decodeList_T_552; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_554 = _decodeList_T_127 ? 7'h0 : _decodeList_T_553; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_555 = _decodeList_T_125 ? 7'hf : _decodeList_T_554; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_556 = _decodeList_T_123 ? 7'he : _decodeList_T_555; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_557 = _decodeList_T_121 ? 7'hd : _decodeList_T_556; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_558 = _decodeList_T_119 ? 7'hc : _decodeList_T_557; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_559 = _decodeList_T_117 ? 7'h8 : _decodeList_T_558; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_560 = _decodeList_T_115 ? 7'h7 : _decodeList_T_559; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_561 = _decodeList_T_113 ? 7'h6 : _decodeList_T_560; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_562 = _decodeList_T_111 ? 7'h5 : _decodeList_T_561; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_563 = _decodeList_T_109 ? 7'h4 : _decodeList_T_562; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_564 = _decodeList_T_107 ? 7'h3 : _decodeList_T_563; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_565 = _decodeList_T_105 ? 7'h2 : _decodeList_T_564; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_566 = _decodeList_T_103 ? 7'h1 : _decodeList_T_565; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_567 = _decodeList_T_101 ? 7'h0 : _decodeList_T_566; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_568 = _decodeList_T_99 ? 7'h2 : _decodeList_T_567; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_569 = _decodeList_T_97 ? 7'hb : _decodeList_T_568; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_570 = _decodeList_T_95 ? 7'h3 : _decodeList_T_569; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_571 = _decodeList_T_93 ? 7'h6 : _decodeList_T_570; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_572 = _decodeList_T_91 ? 7'h28 : _decodeList_T_571; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_573 = _decodeList_T_89 ? 7'h60 : _decodeList_T_572; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_574 = _decodeList_T_87 ? 7'h2d : _decodeList_T_573; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_575 = _decodeList_T_85 ? 7'h25 : _decodeList_T_574; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_576 = _decodeList_T_83 ? 7'h21 : _decodeList_T_575; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_577 = _decodeList_T_81 ? 7'h2d : _decodeList_T_576; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_578 = _decodeList_T_79 ? 7'h25 : _decodeList_T_577; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_579 = _decodeList_T_77 ? 7'h21 : _decodeList_T_578; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_580 = _decodeList_T_75 ? 7'h60 : _decodeList_T_579; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_581 = _decodeList_T_73 ? 7'ha : _decodeList_T_580; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_582 = _decodeList_T_71 ? 7'h9 : _decodeList_T_581; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_583 = _decodeList_T_69 ? 7'h8 : _decodeList_T_582; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_584 = _decodeList_T_67 ? 7'h5 : _decodeList_T_583; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_585 = _decodeList_T_65 ? 7'h4 : _decodeList_T_584; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_586 = _decodeList_T_63 ? 7'h2 : _decodeList_T_585; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_587 = _decodeList_T_61 ? 7'h1 : _decodeList_T_586; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_588 = _decodeList_T_59 ? 7'h0 : _decodeList_T_587; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_589 = _decodeList_T_57 ? 7'h17 : _decodeList_T_588; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_590 = _decodeList_T_55 ? 7'h16 : _decodeList_T_589; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_591 = _decodeList_T_53 ? 7'h15 : _decodeList_T_590; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_592 = _decodeList_T_51 ? 7'h14 : _decodeList_T_591; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_593 = _decodeList_T_49 ? 7'h11 : _decodeList_T_592; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_594 = _decodeList_T_47 ? 7'h10 : _decodeList_T_593; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_595 = _decodeList_T_45 ? 7'h5a : _decodeList_T_594; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_596 = _decodeList_T_43 ? 7'h58 : _decodeList_T_595; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_597 = _decodeList_T_41 ? 7'h40 : _decodeList_T_596; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_598 = _decodeList_T_39 ? 7'h40 : _decodeList_T_597; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_599 = _decodeList_T_37 ? 7'hd : _decodeList_T_598; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_600 = _decodeList_T_35 ? 7'h8 : _decodeList_T_599; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_601 = _decodeList_T_33 ? 7'h7 : _decodeList_T_600; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_602 = _decodeList_T_31 ? 7'h6 : _decodeList_T_601; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_603 = _decodeList_T_29 ? 7'h5 : _decodeList_T_602; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_604 = _decodeList_T_27 ? 7'h4 : _decodeList_T_603; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_605 = _decodeList_T_25 ? 7'h3 : _decodeList_T_604; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_606 = _decodeList_T_23 ? 7'h2 : _decodeList_T_605; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_607 = _decodeList_T_21 ? 7'h1 : _decodeList_T_606; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_608 = _decodeList_T_19 ? 7'h40 : _decodeList_T_607; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_609 = _decodeList_T_17 ? 7'hd : _decodeList_T_608; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_610 = _decodeList_T_15 ? 7'h7 : _decodeList_T_609; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_611 = _decodeList_T_13 ? 7'h6 : _decodeList_T_610; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_612 = _decodeList_T_11 ? 7'h5 : _decodeList_T_611; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_613 = _decodeList_T_9 ? 7'h4 : _decodeList_T_612; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_614 = _decodeList_T_7 ? 7'h3 : _decodeList_T_613; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_615 = _decodeList_T_5 ? 7'h2 : _decodeList_T_614; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_616 = _decodeList_T_3 ? 7'h1 : _decodeList_T_615; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] decodeList_2 = _decodeList_T_1 ? 7'h40 : _decodeList_T_616; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  hasIntr = |intrVecIDU; // @[src/main/scala/nutcore/frontend/IDU.scala 172:22]
  wire [3:0] instrType = hasIntr | io_in_bits_exceptionVec_12 | io_out_bits_cf_exceptionVec_1 ? 4'h0 : decodeList_0; // @[src/main/scala/nutcore/frontend/IDU.scala 38:75]
  wire [2:0] fuType = hasIntr | io_in_bits_exceptionVec_12 | io_out_bits_cf_exceptionVec_1 ? 3'h3 : decodeList_1; // @[src/main/scala/nutcore/frontend/IDU.scala 38:75]
  wire [6:0] fuOpType = hasIntr | io_in_bits_exceptionVec_12 | io_out_bits_cf_exceptionVec_1 ? 7'h0 : decodeList_2; // @[src/main/scala/nutcore/frontend/IDU.scala 38:75]
  wire  isRVC = io_in_bits_instr[1:0] != 2'h3; // @[src/main/scala/nutcore/frontend/IDU.scala 40:45]
  wire [4:0] _T_72 = _decodeList_T_193 ? 5'h3 : 5'h10; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _T_73 = _decodeList_T_191 ? 5'h2 : _T_72; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _T_74 = _decodeList_T_189 ? 5'h10 : _T_73; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _T_75 = _decodeList_T_187 ? 5'h10 : _T_74; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _T_76 = _decodeList_T_185 ? 5'hf : _T_75; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _T_77 = _decodeList_T_183 ? 5'h10 : _T_76; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _T_78 = _decodeList_T_181 ? 5'h10 : _T_77; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _T_79 = _decodeList_T_179 ? 5'h1 : _T_78; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _T_80 = _decodeList_T_177 ? 5'h0 : _T_79; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _T_81 = _decodeList_T_175 ? 5'ha : _T_80; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _T_82 = _decodeList_T_173 ? 5'h9 : _T_81; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _T_83 = _decodeList_T_171 ? 5'h9 : _T_82; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _T_84 = _decodeList_T_169 ? 5'h8 : _T_83; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _T_85 = _decodeList_T_167 ? 5'h10 : _T_84; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _T_86 = _decodeList_T_165 ? 5'h10 : _T_85; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _T_87 = _decodeList_T_163 ? 5'h10 : _T_86; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _T_88 = _decodeList_T_161 ? 5'h10 : _T_87; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _T_89 = _decodeList_T_159 ? 5'h10 : _T_88; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _T_90 = _decodeList_T_157 ? 5'h10 : _T_89; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _T_91 = _decodeList_T_155 ? 5'ha : _T_90; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _T_92 = _decodeList_T_153 ? 5'ha : _T_91; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _T_93 = _decodeList_T_151 ? 5'ha : _T_92; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _T_94 = _decodeList_T_149 ? 5'hb : _T_93; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _T_95 = _decodeList_T_147 ? 5'hd : _T_94; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _T_96 = _decodeList_T_145 ? 5'ha : _T_95; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _T_97 = _decodeList_T_143 ? 5'hc : _T_96; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _T_98 = _decodeList_T_141 ? 5'hc : _T_97; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _T_99 = _decodeList_T_139 ? 5'h10 : _T_98; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _T_100 = _decodeList_T_137 ? 5'h5 : _T_99; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _T_101 = _decodeList_T_135 ? 5'h4 : _T_100; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _T_102 = _decodeList_T_133 ? 5'h7 : _T_101; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _T_103 = _decodeList_T_131 ? 5'h6 : _T_102; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] rvcImmType = _decodeList_T_129 ? 5'he : _T_103; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _T_104 = _decodeList_T_193 ? 4'h9 : 4'h0; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _T_105 = _decodeList_T_191 ? 4'h9 : _T_104; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _T_106 = _decodeList_T_189 ? 4'h2 : _T_105; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _T_107 = _decodeList_T_187 ? 4'h4 : _T_106; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _T_108 = _decodeList_T_185 ? 4'h0 : _T_107; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _T_109 = _decodeList_T_183 ? 4'h5 : _T_108; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _T_110 = _decodeList_T_181 ? 4'h4 : _T_109; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _T_111 = _decodeList_T_179 ? 4'h9 : _T_110; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _T_112 = _decodeList_T_177 ? 4'h9 : _T_111; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _T_113 = _decodeList_T_175 ? 4'h2 : _T_112; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _T_114 = _decodeList_T_173 ? 4'h6 : _T_113; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _T_115 = _decodeList_T_171 ? 4'h6 : _T_114; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _T_116 = _decodeList_T_169 ? 4'h0 : _T_115; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _T_117 = _decodeList_T_167 ? 4'h6 : _T_116; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _T_118 = _decodeList_T_165 ? 4'h6 : _T_117; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _T_119 = _decodeList_T_163 ? 4'h6 : _T_118; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _T_120 = _decodeList_T_161 ? 4'h6 : _T_119; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _T_121 = _decodeList_T_159 ? 4'h6 : _T_120; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _T_122 = _decodeList_T_157 ? 4'h6 : _T_121; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _T_123 = _decodeList_T_155 ? 4'h6 : _T_122; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _T_124 = _decodeList_T_153 ? 4'h6 : _T_123; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _T_125 = _decodeList_T_151 ? 4'h6 : _T_124; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _T_126 = _decodeList_T_149 ? 4'h0 : _T_125; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _T_127 = _decodeList_T_147 ? 4'h9 : _T_126; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _T_128 = _decodeList_T_145 ? 4'h0 : _T_127; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _T_129 = _decodeList_T_143 ? 4'h2 : _T_128; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _T_130 = _decodeList_T_141 ? 4'h2 : _T_129; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _T_131 = _decodeList_T_139 ? 4'h0 : _T_130; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _T_132 = _decodeList_T_137 ? 4'h6 : _T_131; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _T_133 = _decodeList_T_135 ? 4'h6 : _T_132; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _T_134 = _decodeList_T_133 ? 4'h6 : _T_133; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _T_135 = _decodeList_T_131 ? 4'h6 : _T_134; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] rvcSrc1Type = _decodeList_T_129 ? 4'h9 : _T_135; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _T_136 = _decodeList_T_193 ? 3'h5 : 3'h0; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _T_137 = _decodeList_T_191 ? 3'h5 : _T_136; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _T_138 = _decodeList_T_189 ? 3'h5 : _T_137; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _T_139 = _decodeList_T_187 ? 3'h0 : _T_138; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _T_140 = _decodeList_T_185 ? 3'h0 : _T_139; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _T_141 = _decodeList_T_183 ? 3'h0 : _T_140; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _T_142 = _decodeList_T_181 ? 3'h0 : _T_141; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _T_143 = _decodeList_T_179 ? 3'h0 : _T_142; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _T_144 = _decodeList_T_177 ? 3'h0 : _T_143; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _T_145 = _decodeList_T_175 ? 3'h0 : _T_144; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _T_146 = _decodeList_T_173 ? 3'h0 : _T_145; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _T_147 = _decodeList_T_171 ? 3'h0 : _T_146; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _T_148 = _decodeList_T_169 ? 3'h0 : _T_147; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _T_149 = _decodeList_T_167 ? 3'h7 : _T_148; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _T_150 = _decodeList_T_165 ? 3'h7 : _T_149; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _T_151 = _decodeList_T_163 ? 3'h7 : _T_150; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _T_152 = _decodeList_T_161 ? 3'h7 : _T_151; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _T_153 = _decodeList_T_159 ? 3'h7 : _T_152; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _T_154 = _decodeList_T_157 ? 3'h7 : _T_153; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _T_155 = _decodeList_T_155 ? 3'h0 : _T_154; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _T_156 = _decodeList_T_153 ? 3'h0 : _T_155; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _T_157 = _decodeList_T_151 ? 3'h0 : _T_156; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _T_158 = _decodeList_T_149 ? 3'h0 : _T_157; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _T_159 = _decodeList_T_147 ? 3'h0 : _T_158; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _T_160 = _decodeList_T_145 ? 3'h0 : _T_159; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _T_161 = _decodeList_T_143 ? 3'h0 : _T_160; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _T_162 = _decodeList_T_141 ? 3'h0 : _T_161; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _T_163 = _decodeList_T_139 ? 3'h0 : _T_162; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _T_164 = _decodeList_T_137 ? 3'h7 : _T_163; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _T_165 = _decodeList_T_135 ? 3'h7 : _T_164; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _T_166 = _decodeList_T_133 ? 3'h0 : _T_165; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _T_167 = _decodeList_T_131 ? 3'h0 : _T_166; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] rvcSrc2Type = _decodeList_T_129 ? 3'h0 : _T_167; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [1:0] _T_170 = _decodeList_T_189 ? 2'h2 : 2'h0; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _T_171 = _decodeList_T_187 ? 4'h8 : {{2'd0}, _T_170}; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _T_172 = _decodeList_T_185 ? 4'h0 : _T_171; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _T_173 = _decodeList_T_183 ? 4'h2 : _T_172; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _T_174 = _decodeList_T_181 ? 4'h0 : _T_173; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _T_175 = _decodeList_T_179 ? 4'h2 : _T_174; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _T_176 = _decodeList_T_177 ? 4'h2 : _T_175; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _T_177 = _decodeList_T_175 ? 4'h2 : _T_176; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _T_178 = _decodeList_T_173 ? 4'h0 : _T_177; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _T_179 = _decodeList_T_171 ? 4'h0 : _T_178; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _T_180 = _decodeList_T_169 ? 4'h0 : _T_179; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _T_181 = _decodeList_T_167 ? 4'h6 : _T_180; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _T_182 = _decodeList_T_165 ? 4'h6 : _T_181; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _T_183 = _decodeList_T_163 ? 4'h6 : _T_182; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _T_184 = _decodeList_T_161 ? 4'h6 : _T_183; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _T_185 = _decodeList_T_159 ? 4'h6 : _T_184; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _T_186 = _decodeList_T_157 ? 4'h6 : _T_185; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _T_187 = _decodeList_T_155 ? 4'h6 : _T_186; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _T_188 = _decodeList_T_153 ? 4'h6 : _T_187; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _T_189 = _decodeList_T_151 ? 4'h6 : _T_188; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _T_190 = _decodeList_T_149 ? 4'h2 : _T_189; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _T_191 = _decodeList_T_147 ? 4'h9 : _T_190; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _T_192 = _decodeList_T_145 ? 4'h2 : _T_191; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _T_193 = _decodeList_T_143 ? 4'h2 : _T_192; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _T_194 = _decodeList_T_141 ? 4'h2 : _T_193; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _T_195 = _decodeList_T_139 ? 4'h0 : _T_194; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _T_196 = _decodeList_T_137 ? 4'h0 : _T_195; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _T_197 = _decodeList_T_135 ? 4'h0 : _T_196; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _T_198 = _decodeList_T_133 ? 4'h7 : _T_197; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _T_199 = _decodeList_T_131 ? 4'h7 : _T_198; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] rvcDestType = _decodeList_T_129 ? 4'h7 : _T_199; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _src1Type_T = 4'h4 == instrType; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _src1Type_T_2 = 4'h2 == instrType; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _src1Type_T_3 = 4'hf == instrType; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _src1Type_T_4 = 4'h1 == instrType; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _src1Type_T_5 = 4'h6 == instrType; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _src1Type_T_6 = 4'h7 == instrType; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _src1Type_T_7 = 4'h0 == instrType; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  src1Type = _src1Type_T_5 | _src1Type_T_6 | _src1Type_T_7; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  src2Type = _src1Type_T | _src1Type_T_5 | _src1Type_T_6 | _src1Type_T_7; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [4:0] rs = io_in_bits_instr[19:15]; // @[src/main/scala/nutcore/frontend/IDU.scala 62:28]
  wire [4:0] rt = io_in_bits_instr[24:20]; // @[src/main/scala/nutcore/frontend/IDU.scala 62:43]
  wire [4:0] rd = io_in_bits_instr[11:7]; // @[src/main/scala/nutcore/frontend/IDU.scala 62:58]
  wire [4:0] rs2 = io_in_bits_instr[6:2]; // @[src/main/scala/nutcore/frontend/IDU.scala 65:24]
  wire  _rs1p_T_1 = 3'h0 == io_in_bits_instr[9:7]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _rs1p_T_2 = 3'h1 == io_in_bits_instr[9:7]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _rs1p_T_3 = 3'h2 == io_in_bits_instr[9:7]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _rs1p_T_4 = 3'h3 == io_in_bits_instr[9:7]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _rs1p_T_5 = 3'h4 == io_in_bits_instr[9:7]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _rs1p_T_6 = 3'h5 == io_in_bits_instr[9:7]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _rs1p_T_7 = 3'h6 == io_in_bits_instr[9:7]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _rs1p_T_8 = 3'h7 == io_in_bits_instr[9:7]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [3:0] _rs1p_T_9 = _rs1p_T_1 ? 4'h8 : 4'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [3:0] _rs1p_T_10 = _rs1p_T_2 ? 4'h9 : 4'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [3:0] _rs1p_T_11 = _rs1p_T_3 ? 4'ha : 4'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [3:0] _rs1p_T_12 = _rs1p_T_4 ? 4'hb : 4'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [3:0] _rs1p_T_13 = _rs1p_T_5 ? 4'hc : 4'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [3:0] _rs1p_T_14 = _rs1p_T_6 ? 4'hd : 4'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [3:0] _rs1p_T_15 = _rs1p_T_7 ? 4'he : 4'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [3:0] _rs1p_T_16 = _rs1p_T_8 ? 4'hf : 4'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [3:0] _rs1p_T_17 = _rs1p_T_9 | _rs1p_T_10; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [3:0] _rs1p_T_18 = _rs1p_T_17 | _rs1p_T_11; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [3:0] _rs1p_T_19 = _rs1p_T_18 | _rs1p_T_12; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [3:0] _rs1p_T_20 = _rs1p_T_19 | _rs1p_T_13; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [3:0] _rs1p_T_21 = _rs1p_T_20 | _rs1p_T_14; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [3:0] _rs1p_T_22 = _rs1p_T_21 | _rs1p_T_15; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [3:0] rs1p = _rs1p_T_22 | _rs1p_T_16; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rs2p_T_1 = 3'h0 == io_in_bits_instr[4:2]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _rs2p_T_2 = 3'h1 == io_in_bits_instr[4:2]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _rs2p_T_3 = 3'h2 == io_in_bits_instr[4:2]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _rs2p_T_4 = 3'h3 == io_in_bits_instr[4:2]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _rs2p_T_5 = 3'h4 == io_in_bits_instr[4:2]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _rs2p_T_6 = 3'h5 == io_in_bits_instr[4:2]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _rs2p_T_7 = 3'h6 == io_in_bits_instr[4:2]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _rs2p_T_8 = 3'h7 == io_in_bits_instr[4:2]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [3:0] _rs2p_T_9 = _rs2p_T_1 ? 4'h8 : 4'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [3:0] _rs2p_T_10 = _rs2p_T_2 ? 4'h9 : 4'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [3:0] _rs2p_T_11 = _rs2p_T_3 ? 4'ha : 4'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [3:0] _rs2p_T_12 = _rs2p_T_4 ? 4'hb : 4'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [3:0] _rs2p_T_13 = _rs2p_T_5 ? 4'hc : 4'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [3:0] _rs2p_T_14 = _rs2p_T_6 ? 4'hd : 4'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [3:0] _rs2p_T_15 = _rs2p_T_7 ? 4'he : 4'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [3:0] _rs2p_T_16 = _rs2p_T_8 ? 4'hf : 4'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [3:0] _rs2p_T_17 = _rs2p_T_9 | _rs2p_T_10; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [3:0] _rs2p_T_18 = _rs2p_T_17 | _rs2p_T_11; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [3:0] _rs2p_T_19 = _rs2p_T_18 | _rs2p_T_12; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [3:0] _rs2p_T_20 = _rs2p_T_19 | _rs2p_T_13; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [3:0] _rs2p_T_21 = _rs2p_T_20 | _rs2p_T_14; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [3:0] _rs2p_T_22 = _rs2p_T_21 | _rs2p_T_15; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [3:0] rs2p = _rs2p_T_22 | _rs2p_T_16; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [5:0] rvc_shamt = {io_in_bits_instr[12],rs2}; // @[src/main/scala/nutcore/frontend/IDU.scala 68:22]
  wire  _rvc_src1_T_1 = 4'h3 == rvcSrc1Type; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _rvc_src1_T_2 = 4'h1 == rvcSrc1Type; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _rvc_src1_T_3 = 4'h2 == rvcSrc1Type; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _rvc_src1_T_4 = 4'h4 == rvcSrc1Type; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _rvc_src1_T_5 = 4'h5 == rvcSrc1Type; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _rvc_src1_T_6 = 4'h6 == rvcSrc1Type; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _rvc_src1_T_7 = 4'h7 == rvcSrc1Type; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _rvc_src1_T_8 = 4'h8 == rvcSrc1Type; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _rvc_src1_T_9 = 4'h9 == rvcSrc1Type; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [4:0] _rvc_src1_T_11 = _rvc_src1_T_1 ? rs : 5'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [4:0] _rvc_src1_T_12 = _rvc_src1_T_2 ? rt : 5'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [4:0] _rvc_src1_T_13 = _rvc_src1_T_3 ? rd : 5'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [4:0] _rvc_src1_T_14 = _rvc_src1_T_4 ? rd : 5'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [4:0] _rvc_src1_T_15 = _rvc_src1_T_5 ? rs2 : 5'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [3:0] _rvc_src1_T_16 = _rvc_src1_T_6 ? rs1p : 4'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [3:0] _rvc_src1_T_17 = _rvc_src1_T_7 ? rs2p : 4'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [1:0] _rvc_src1_T_19 = _rvc_src1_T_9 ? 2'h2 : 2'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [4:0] _rvc_src1_T_21 = _rvc_src1_T_11 | _rvc_src1_T_12; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [4:0] _rvc_src1_T_22 = _rvc_src1_T_21 | _rvc_src1_T_13; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [4:0] _rvc_src1_T_23 = _rvc_src1_T_22 | _rvc_src1_T_14; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [4:0] _rvc_src1_T_24 = _rvc_src1_T_23 | _rvc_src1_T_15; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [4:0] _GEN_5 = {{1'd0}, _rvc_src1_T_16}; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [4:0] _rvc_src1_T_25 = _rvc_src1_T_24 | _GEN_5; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [4:0] _GEN_6 = {{1'd0}, _rvc_src1_T_17}; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [4:0] _rvc_src1_T_26 = _rvc_src1_T_25 | _GEN_6; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [4:0] _GEN_7 = {{4'd0}, _rvc_src1_T_8}; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [4:0] _rvc_src1_T_27 = _rvc_src1_T_26 | _GEN_7; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [4:0] _GEN_8 = {{3'd0}, _rvc_src1_T_19}; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [4:0] rvc_src1 = _rvc_src1_T_27 | _GEN_8; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rvc_src2_T_1 = 3'h3 == rvcSrc2Type; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _rvc_src2_T_2 = 3'h1 == rvcSrc2Type; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _rvc_src2_T_3 = 3'h2 == rvcSrc2Type; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _rvc_src2_T_4 = 3'h4 == rvcSrc2Type; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _rvc_src2_T_5 = 3'h5 == rvcSrc2Type; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _rvc_src2_T_6 = 3'h6 == rvcSrc2Type; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _rvc_src2_T_7 = 3'h7 == rvcSrc2Type; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [3:0] _GEN_9 = {{1'd0}, rvcSrc2Type}; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _rvc_src2_T_8 = 4'h8 == _GEN_9; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _rvc_src2_T_9 = 4'h9 == _GEN_9; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [4:0] _rvc_src2_T_11 = _rvc_src2_T_1 ? rs : 5'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [4:0] _rvc_src2_T_12 = _rvc_src2_T_2 ? rt : 5'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [4:0] _rvc_src2_T_13 = _rvc_src2_T_3 ? rd : 5'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [4:0] _rvc_src2_T_14 = _rvc_src2_T_4 ? rd : 5'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [4:0] _rvc_src2_T_15 = _rvc_src2_T_5 ? rs2 : 5'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [3:0] _rvc_src2_T_16 = _rvc_src2_T_6 ? rs1p : 4'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [3:0] _rvc_src2_T_17 = _rvc_src2_T_7 ? rs2p : 4'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [1:0] _rvc_src2_T_19 = _rvc_src2_T_9 ? 2'h2 : 2'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [4:0] _rvc_src2_T_21 = _rvc_src2_T_11 | _rvc_src2_T_12; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [4:0] _rvc_src2_T_22 = _rvc_src2_T_21 | _rvc_src2_T_13; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [4:0] _rvc_src2_T_23 = _rvc_src2_T_22 | _rvc_src2_T_14; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [4:0] _rvc_src2_T_24 = _rvc_src2_T_23 | _rvc_src2_T_15; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [4:0] _GEN_11 = {{1'd0}, _rvc_src2_T_16}; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [4:0] _rvc_src2_T_25 = _rvc_src2_T_24 | _GEN_11; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [4:0] _GEN_12 = {{1'd0}, _rvc_src2_T_17}; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [4:0] _rvc_src2_T_26 = _rvc_src2_T_25 | _GEN_12; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [4:0] _GEN_13 = {{4'd0}, _rvc_src2_T_8}; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [4:0] _rvc_src2_T_27 = _rvc_src2_T_26 | _GEN_13; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [4:0] _GEN_14 = {{3'd0}, _rvc_src2_T_19}; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [4:0] rvc_src2 = _rvc_src2_T_27 | _GEN_14; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rvc_dest_T_1 = 4'h3 == rvcDestType; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _rvc_dest_T_2 = 4'h1 == rvcDestType; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _rvc_dest_T_3 = 4'h2 == rvcDestType; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _rvc_dest_T_4 = 4'h4 == rvcDestType; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _rvc_dest_T_5 = 4'h5 == rvcDestType; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _rvc_dest_T_6 = 4'h6 == rvcDestType; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _rvc_dest_T_7 = 4'h7 == rvcDestType; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _rvc_dest_T_8 = 4'h8 == rvcDestType; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _rvc_dest_T_9 = 4'h9 == rvcDestType; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [4:0] _rvc_dest_T_11 = _rvc_dest_T_1 ? rs : 5'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [4:0] _rvc_dest_T_12 = _rvc_dest_T_2 ? rt : 5'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [4:0] _rvc_dest_T_13 = _rvc_dest_T_3 ? rd : 5'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [4:0] _rvc_dest_T_14 = _rvc_dest_T_4 ? rd : 5'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [4:0] _rvc_dest_T_15 = _rvc_dest_T_5 ? rs2 : 5'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [3:0] _rvc_dest_T_16 = _rvc_dest_T_6 ? rs1p : 4'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [3:0] _rvc_dest_T_17 = _rvc_dest_T_7 ? rs2p : 4'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [1:0] _rvc_dest_T_19 = _rvc_dest_T_9 ? 2'h2 : 2'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [4:0] _rvc_dest_T_21 = _rvc_dest_T_11 | _rvc_dest_T_12; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [4:0] _rvc_dest_T_22 = _rvc_dest_T_21 | _rvc_dest_T_13; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [4:0] _rvc_dest_T_23 = _rvc_dest_T_22 | _rvc_dest_T_14; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [4:0] _rvc_dest_T_24 = _rvc_dest_T_23 | _rvc_dest_T_15; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [4:0] _GEN_15 = {{1'd0}, _rvc_dest_T_16}; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [4:0] _rvc_dest_T_25 = _rvc_dest_T_24 | _GEN_15; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [4:0] _GEN_16 = {{1'd0}, _rvc_dest_T_17}; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [4:0] _rvc_dest_T_26 = _rvc_dest_T_25 | _GEN_16; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [4:0] _GEN_17 = {{4'd0}, _rvc_dest_T_8}; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [4:0] _rvc_dest_T_27 = _rvc_dest_T_26 | _GEN_17; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [4:0] _GEN_18 = {{3'd0}, _rvc_dest_T_19}; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [4:0] rvc_dest = _rvc_dest_T_27 | _GEN_18; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [4:0] rfSrc1 = isRVC ? rvc_src1 : rs; // @[src/main/scala/nutcore/frontend/IDU.scala 89:19]
  wire [4:0] rfSrc2 = isRVC ? rvc_src2 : rt; // @[src/main/scala/nutcore/frontend/IDU.scala 90:19]
  wire [4:0] rfDest = isRVC ? rvc_dest : rd; // @[src/main/scala/nutcore/frontend/IDU.scala 91:19]
  wire  imm_signBit = io_in_bits_instr[31]; // @[src/main/scala/utils/BitUtils.scala 41:20]
  wire [51:0] _imm_T_2 = imm_signBit ? 52'hfffffffffffff : 52'h0; // @[src/main/scala/utils/BitUtils.scala 42:46]
  wire [63:0] _imm_T_3 = {_imm_T_2,io_in_bits_instr[31:20]}; // @[src/main/scala/utils/BitUtils.scala 42:41]
  wire [11:0] _imm_T_6 = {io_in_bits_instr[31:25],rd}; // @[src/main/scala/nutcore/frontend/IDU.scala 102:27]
  wire  imm_signBit_1 = _imm_T_6[11]; // @[src/main/scala/utils/BitUtils.scala 41:20]
  wire [51:0] _imm_T_8 = imm_signBit_1 ? 52'hfffffffffffff : 52'h0; // @[src/main/scala/utils/BitUtils.scala 42:46]
  wire [63:0] _imm_T_9 = {_imm_T_8,io_in_bits_instr[31:25],rd}; // @[src/main/scala/utils/BitUtils.scala 42:41]
  wire [12:0] _imm_T_20 = {io_in_bits_instr[31],io_in_bits_instr[7],io_in_bits_instr[30:25],io_in_bits_instr[11:8],1'h0}
    ; // @[src/main/scala/nutcore/frontend/IDU.scala 104:27]
  wire  imm_signBit_3 = _imm_T_20[12]; // @[src/main/scala/utils/BitUtils.scala 41:20]
  wire [50:0] _imm_T_22 = imm_signBit_3 ? 51'h7ffffffffffff : 51'h0; // @[src/main/scala/utils/BitUtils.scala 42:46]
  wire [63:0] _imm_T_23 = {_imm_T_22,io_in_bits_instr[31],io_in_bits_instr[7],io_in_bits_instr[30:25],io_in_bits_instr[
    11:8],1'h0}; // @[src/main/scala/utils/BitUtils.scala 42:41]
  wire [31:0] _imm_T_25 = {io_in_bits_instr[31:12],12'h0}; // @[src/main/scala/nutcore/frontend/IDU.scala 105:27]
  wire  imm_signBit_4 = _imm_T_25[31]; // @[src/main/scala/utils/BitUtils.scala 41:20]
  wire [31:0] _imm_T_27 = imm_signBit_4 ? 32'hffffffff : 32'h0; // @[src/main/scala/utils/BitUtils.scala 42:46]
  wire [63:0] _imm_T_28 = {_imm_T_27,io_in_bits_instr[31:12],12'h0}; // @[src/main/scala/utils/BitUtils.scala 42:41]
  wire [20:0] _imm_T_33 = {io_in_bits_instr[31],io_in_bits_instr[19:12],io_in_bits_instr[20],io_in_bits_instr[30:21],1'h0
    }; // @[src/main/scala/nutcore/frontend/IDU.scala 106:27]
  wire  imm_signBit_5 = _imm_T_33[20]; // @[src/main/scala/utils/BitUtils.scala 41:20]
  wire [42:0] _imm_T_35 = imm_signBit_5 ? 43'h7ffffffffff : 43'h0; // @[src/main/scala/utils/BitUtils.scala 42:46]
  wire [63:0] _imm_T_36 = {_imm_T_35,io_in_bits_instr[31],io_in_bits_instr[19:12],io_in_bits_instr[20],io_in_bits_instr[
    30:21],1'h0}; // @[src/main/scala/utils/BitUtils.scala 42:41]
  wire [63:0] _imm_T_43 = _src1Type_T ? _imm_T_3 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _imm_T_44 = _src1Type_T_2 ? _imm_T_9 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _imm_T_45 = _src1Type_T_3 ? _imm_T_9 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _imm_T_46 = _src1Type_T_4 ? _imm_T_23 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _imm_T_47 = _src1Type_T_5 ? _imm_T_28 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _imm_T_48 = _src1Type_T_6 ? _imm_T_36 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _imm_T_49 = _imm_T_43 | _imm_T_44; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _imm_T_50 = _imm_T_49 | _imm_T_45; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _imm_T_51 = _imm_T_50 | _imm_T_46; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _imm_T_52 = _imm_T_51 | _imm_T_47; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] imm = _imm_T_52 | _imm_T_48; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _immrvc_T_4 = {56'h0,io_in_bits_instr[3:2],io_in_bits_instr[12],io_in_bits_instr[6:4],2'h0}; // @[src/main/scala/utils/BitUtils.scala 49:41]
  wire [63:0] _immrvc_T_9 = {55'h0,io_in_bits_instr[4:2],io_in_bits_instr[12],io_in_bits_instr[6:5],3'h0}; // @[src/main/scala/utils/BitUtils.scala 49:41]
  wire [63:0] _immrvc_T_13 = {56'h0,io_in_bits_instr[8:7],io_in_bits_instr[12:9],2'h0}; // @[src/main/scala/utils/BitUtils.scala 49:41]
  wire [63:0] _immrvc_T_17 = {55'h0,io_in_bits_instr[9:7],io_in_bits_instr[12:10],3'h0}; // @[src/main/scala/utils/BitUtils.scala 49:41]
  wire [63:0] _immrvc_T_22 = {57'h0,io_in_bits_instr[5],io_in_bits_instr[12:10],io_in_bits_instr[6],2'h0}; // @[src/main/scala/utils/BitUtils.scala 49:41]
  wire [63:0] _immrvc_T_26 = {56'h0,io_in_bits_instr[6:5],io_in_bits_instr[12:10],3'h0}; // @[src/main/scala/utils/BitUtils.scala 49:41]
  wire [11:0] _immrvc_T_44 = {io_in_bits_instr[12],io_in_bits_instr[8],io_in_bits_instr[10:9],io_in_bits_instr[6],
    io_in_bits_instr[7],io_in_bits_instr[2],io_in_bits_instr[11],io_in_bits_instr[5:3],1'h0}; // @[src/main/scala/nutcore/frontend/IDU.scala 119:37]
  wire  immrvc_signBit = _immrvc_T_44[11]; // @[src/main/scala/utils/BitUtils.scala 41:20]
  wire [51:0] _immrvc_T_46 = immrvc_signBit ? 52'hfffffffffffff : 52'h0; // @[src/main/scala/utils/BitUtils.scala 42:46]
  wire [63:0] _immrvc_T_47 = {_immrvc_T_46,io_in_bits_instr[12],io_in_bits_instr[8],io_in_bits_instr[10:9],
    io_in_bits_instr[6],io_in_bits_instr[7],io_in_bits_instr[2],io_in_bits_instr[11],io_in_bits_instr[5:3],1'h0}; // @[src/main/scala/utils/BitUtils.scala 42:41]
  wire [8:0] _immrvc_T_53 = {io_in_bits_instr[12],io_in_bits_instr[6:5],io_in_bits_instr[2],io_in_bits_instr[11:10],
    io_in_bits_instr[4:3],1'h0}; // @[src/main/scala/nutcore/frontend/IDU.scala 120:37]
  wire  immrvc_signBit_1 = _immrvc_T_53[8]; // @[src/main/scala/utils/BitUtils.scala 41:20]
  wire [54:0] _immrvc_T_55 = immrvc_signBit_1 ? 55'h7fffffffffffff : 55'h0; // @[src/main/scala/utils/BitUtils.scala 42:46]
  wire [63:0] _immrvc_T_56 = {_immrvc_T_55,io_in_bits_instr[12],io_in_bits_instr[6:5],io_in_bits_instr[2],
    io_in_bits_instr[11:10],io_in_bits_instr[4:3],1'h0}; // @[src/main/scala/utils/BitUtils.scala 42:41]
  wire  immrvc_signBit_2 = rvc_shamt[5]; // @[src/main/scala/utils/BitUtils.scala 41:20]
  wire [57:0] _immrvc_T_61 = immrvc_signBit_2 ? 58'h3ffffffffffffff : 58'h0; // @[src/main/scala/utils/BitUtils.scala 42:46]
  wire [63:0] _immrvc_T_62 = {_immrvc_T_61,io_in_bits_instr[12],rs2}; // @[src/main/scala/utils/BitUtils.scala 42:41]
  wire [17:0] _immrvc_T_65 = {io_in_bits_instr[12],rs2,12'h0}; // @[src/main/scala/nutcore/frontend/IDU.scala 122:37]
  wire  immrvc_signBit_3 = _immrvc_T_65[17]; // @[src/main/scala/utils/BitUtils.scala 41:20]
  wire [45:0] _immrvc_T_67 = immrvc_signBit_3 ? 46'h3fffffffffff : 46'h0; // @[src/main/scala/utils/BitUtils.scala 42:46]
  wire [63:0] _immrvc_T_68 = {_immrvc_T_67,io_in_bits_instr[12],rs2,12'h0}; // @[src/main/scala/utils/BitUtils.scala 42:41]
  wire [9:0] _immrvc_T_80 = {io_in_bits_instr[12],io_in_bits_instr[4:3],io_in_bits_instr[5],io_in_bits_instr[2],
    io_in_bits_instr[6],4'h0}; // @[src/main/scala/nutcore/frontend/IDU.scala 124:39]
  wire  immrvc_signBit_5 = _immrvc_T_80[9]; // @[src/main/scala/utils/BitUtils.scala 41:20]
  wire [53:0] _immrvc_T_82 = immrvc_signBit_5 ? 54'h3fffffffffffff : 54'h0; // @[src/main/scala/utils/BitUtils.scala 42:46]
  wire [63:0] _immrvc_T_83 = {_immrvc_T_82,io_in_bits_instr[12],io_in_bits_instr[4:3],io_in_bits_instr[5],
    io_in_bits_instr[2],io_in_bits_instr[6],4'h0}; // @[src/main/scala/utils/BitUtils.scala 42:41]
  wire [63:0] _immrvc_T_89 = {54'h0,io_in_bits_instr[10:7],io_in_bits_instr[12:11],io_in_bits_instr[5],io_in_bits_instr[
    6],2'h0}; // @[src/main/scala/utils/BitUtils.scala 49:41]
  wire  _immrvc_T_91 = 5'h0 == rvcImmType; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _immrvc_T_92 = 5'h1 == rvcImmType; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _immrvc_T_93 = 5'h2 == rvcImmType; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _immrvc_T_94 = 5'h3 == rvcImmType; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _immrvc_T_95 = 5'h4 == rvcImmType; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _immrvc_T_96 = 5'h5 == rvcImmType; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _immrvc_T_97 = 5'h6 == rvcImmType; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _immrvc_T_98 = 5'h7 == rvcImmType; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _immrvc_T_99 = 5'h8 == rvcImmType; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _immrvc_T_100 = 5'h9 == rvcImmType; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _immrvc_T_101 = 5'ha == rvcImmType; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _immrvc_T_102 = 5'hb == rvcImmType; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _immrvc_T_103 = 5'hc == rvcImmType; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _immrvc_T_104 = 5'hd == rvcImmType; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _immrvc_T_105 = 5'he == rvcImmType; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _immrvc_T_106 = 5'hf == rvcImmType; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _immrvc_T_108 = _immrvc_T_91 ? _immrvc_T_4 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _immrvc_T_109 = _immrvc_T_92 ? _immrvc_T_9 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _immrvc_T_110 = _immrvc_T_93 ? _immrvc_T_13 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _immrvc_T_111 = _immrvc_T_94 ? _immrvc_T_17 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _immrvc_T_112 = _immrvc_T_95 ? _immrvc_T_22 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _immrvc_T_113 = _immrvc_T_96 ? _immrvc_T_26 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _immrvc_T_114 = _immrvc_T_97 ? _immrvc_T_22 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _immrvc_T_115 = _immrvc_T_98 ? _immrvc_T_26 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _immrvc_T_116 = _immrvc_T_99 ? _immrvc_T_47 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _immrvc_T_117 = _immrvc_T_100 ? _immrvc_T_56 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _immrvc_T_118 = _immrvc_T_101 ? _immrvc_T_62 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _immrvc_T_119 = _immrvc_T_102 ? _immrvc_T_68 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _immrvc_T_120 = _immrvc_T_103 ? _immrvc_T_62 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _immrvc_T_121 = _immrvc_T_104 ? _immrvc_T_83 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _immrvc_T_122 = _immrvc_T_105 ? _immrvc_T_89 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _immrvc_T_123 = _immrvc_T_106 ? 64'h1 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _immrvc_T_125 = _immrvc_T_108 | _immrvc_T_109; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _immrvc_T_126 = _immrvc_T_125 | _immrvc_T_110; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _immrvc_T_127 = _immrvc_T_126 | _immrvc_T_111; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _immrvc_T_128 = _immrvc_T_127 | _immrvc_T_112; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _immrvc_T_129 = _immrvc_T_128 | _immrvc_T_113; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _immrvc_T_130 = _immrvc_T_129 | _immrvc_T_114; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _immrvc_T_131 = _immrvc_T_130 | _immrvc_T_115; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _immrvc_T_132 = _immrvc_T_131 | _immrvc_T_116; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _immrvc_T_133 = _immrvc_T_132 | _immrvc_T_117; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _immrvc_T_134 = _immrvc_T_133 | _immrvc_T_118; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _immrvc_T_135 = _immrvc_T_134 | _immrvc_T_119; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _immrvc_T_136 = _immrvc_T_135 | _immrvc_T_120; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _immrvc_T_137 = _immrvc_T_136 | _immrvc_T_121; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _immrvc_T_138 = _immrvc_T_137 | _immrvc_T_122; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] immrvc = _immrvc_T_138 | _immrvc_T_123; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _T_203 = rfDest == 5'h1 | rfDest == 5'h5; // @[src/main/scala/nutcore/frontend/IDU.scala 133:42]
  wire [6:0] _GEN_0 = _T_203 & fuOpType == 7'h58 ? 7'h5c : fuOpType; // @[src/main/scala/nutcore/frontend/IDU.scala 134:{57,85} 47:29]
  wire  _T_209 = rfSrc1 == 5'h1 | rfSrc1 == 5'h5; // @[src/main/scala/nutcore/frontend/IDU.scala 133:42]
  wire [6:0] _GEN_1 = _T_209 ? 7'h5e : _GEN_0; // @[src/main/scala/nutcore/frontend/IDU.scala 136:{29,57}]
  wire [6:0] _GEN_2 = _T_203 ? 7'h5c : _GEN_1; // @[src/main/scala/nutcore/frontend/IDU.scala 137:{29,57}]
  wire [6:0] _GEN_3 = fuOpType == 7'h5a ? _GEN_2 : _GEN_0; // @[src/main/scala/nutcore/frontend/IDU.scala 135:40]
  wire  _io_in_ready_T_1 = io_out_ready & io_out_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  wire  _io_in_ready_T_2 = ~hasIntr; // @[src/main/scala/nutcore/frontend/IDU.scala 162:49]
  reg [63:0] c; // @[src/main/scala/utils/GTimer.scala 24:20]
  wire [63:0] _c_T_1 = c + 64'h1; // @[src/main/scala/utils/GTimer.scala 25:12]
  wire  _T_214 = _io_in_ready_T_1 & DISPLAY_ENABLE; // @[src/main/scala/utils/Debug.scala 55:16]
  wire  _T_216 = ~reset; // @[src/main/scala/utils/Debug.scala 56:24]
  assign io_in_ready = ~io_in_valid | _io_in_ready_T_1 & ~hasIntr; // @[src/main/scala/nutcore/frontend/IDU.scala 162:31]
  assign io_out_valid = io_in_valid; // @[src/main/scala/nutcore/frontend/IDU.scala 161:16]
  assign io_out_bits_cf_instr = io_in_bits_instr; // @[src/main/scala/nutcore/frontend/IDU.scala 163:18]
  assign io_out_bits_cf_pc = io_in_bits_pc; // @[src/main/scala/nutcore/frontend/IDU.scala 163:18]
  assign io_out_bits_cf_pnpc = io_in_bits_pnpc; // @[src/main/scala/nutcore/frontend/IDU.scala 163:18]
  assign io_out_bits_cf_exceptionVec_1 = |io_in_bits_pc[38:32] & ~DTLBENABLE; // @[src/main/scala/nutcore/frontend/IDU.scala 181:98]
  assign io_out_bits_cf_exceptionVec_2 = instrType == 4'h0 & _io_in_ready_T_2 & io_in_valid; // @[src/main/scala/nutcore/frontend/IDU.scala 178:83]
  assign io_out_bits_cf_exceptionVec_12 = io_in_bits_exceptionVec_12; // @[src/main/scala/nutcore/frontend/IDU.scala 179:47]
  assign io_out_bits_cf_intrVec_0 = intrVecIDU[0]; // @[src/main/scala/nutcore/frontend/IDU.scala 171:38]
  assign io_out_bits_cf_intrVec_1 = intrVecIDU[1]; // @[src/main/scala/nutcore/frontend/IDU.scala 171:38]
  assign io_out_bits_cf_intrVec_2 = intrVecIDU[2]; // @[src/main/scala/nutcore/frontend/IDU.scala 171:38]
  assign io_out_bits_cf_intrVec_3 = intrVecIDU[3]; // @[src/main/scala/nutcore/frontend/IDU.scala 171:38]
  assign io_out_bits_cf_intrVec_4 = intrVecIDU[4]; // @[src/main/scala/nutcore/frontend/IDU.scala 171:38]
  assign io_out_bits_cf_intrVec_5 = intrVecIDU[5]; // @[src/main/scala/nutcore/frontend/IDU.scala 171:38]
  assign io_out_bits_cf_intrVec_6 = intrVecIDU[6]; // @[src/main/scala/nutcore/frontend/IDU.scala 171:38]
  assign io_out_bits_cf_intrVec_7 = intrVecIDU[7]; // @[src/main/scala/nutcore/frontend/IDU.scala 171:38]
  assign io_out_bits_cf_intrVec_8 = intrVecIDU[8]; // @[src/main/scala/nutcore/frontend/IDU.scala 171:38]
  assign io_out_bits_cf_intrVec_9 = intrVecIDU[9]; // @[src/main/scala/nutcore/frontend/IDU.scala 171:38]
  assign io_out_bits_cf_intrVec_10 = intrVecIDU[10]; // @[src/main/scala/nutcore/frontend/IDU.scala 171:38]
  assign io_out_bits_cf_intrVec_11 = intrVecIDU[11]; // @[src/main/scala/nutcore/frontend/IDU.scala 171:38]
  assign io_out_bits_cf_brIdx = io_in_bits_brIdx; // @[src/main/scala/nutcore/frontend/IDU.scala 163:18]
  assign io_out_bits_cf_crossPageIPFFix = io_in_bits_crossPageIPFFix; // @[src/main/scala/nutcore/frontend/IDU.scala 163:18]
  assign io_out_bits_ctrl_src1Type = io_in_bits_instr[6:0] == 7'h37 ? 1'h0 : src1Type; // @[src/main/scala/nutcore/frontend/IDU.scala 141:35]
  assign io_out_bits_ctrl_src2Type = _src1Type_T | _src1Type_T_5 | _src1Type_T_6 | _src1Type_T_7; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign io_out_bits_ctrl_fuType = hasIntr | io_in_bits_exceptionVec_12 | io_out_bits_cf_exceptionVec_1 ? 3'h3 :
    decodeList_1; // @[src/main/scala/nutcore/frontend/IDU.scala 38:75]
  assign io_out_bits_ctrl_fuOpType = fuType == 3'h0 ? _GEN_3 : fuOpType; // @[src/main/scala/nutcore/frontend/IDU.scala 132:32 47:29]
  assign io_out_bits_ctrl_rfSrc1 = src1Type ? 5'h0 : rfSrc1; // @[src/main/scala/nutcore/frontend/IDU.scala 94:33]
  assign io_out_bits_ctrl_rfSrc2 = ~src2Type ? rfSrc2 : 5'h0; // @[src/main/scala/nutcore/frontend/IDU.scala 95:33]
  assign io_out_bits_ctrl_rfWen = instrType[2]; // @[src/main/scala/nutcore/Decode.scala 33:50]
  assign io_out_bits_ctrl_rfDest = instrType[2] ? rfDest : 5'h0; // @[src/main/scala/nutcore/frontend/IDU.scala 97:33]
  assign io_out_bits_ctrl_isNutCoreTrap = _decodeList_T_99 & io_in_valid; // @[src/main/scala/nutcore/frontend/IDU.scala 186:66]
  assign io_out_bits_data_imm = isRVC ? immrvc : imm; // @[src/main/scala/nutcore/frontend/IDU.scala 130:31]
  assign io_isWFI = _decodeList_T_203 & io_in_valid; // @[src/main/scala/nutcore/frontend/IDU.scala 187:43]
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/utils/GTimer.scala 24:20]
      c <= 64'h0; // @[src/main/scala/utils/GTimer.scala 24:20]
    end else begin
      c <= _c_T_1; // @[src/main/scala/utils/GTimer.scala 25:7]
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_214 & ~reset) begin
          $fwrite(32'h80000002,"[%d] Decoder: ",c); // @[src/main/scala/utils/Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_214 & _T_216) begin
          $fwrite(32'h80000002,"issue: pc %x npc %x instr %x\n",io_out_bits_cf_pc,io_out_bits_cf_pnpc,
            io_out_bits_cf_instr); // @[src/main/scala/utils/Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  c = _RAND_0[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Decoder_1(
  input         clock,
  input         reset,
  output        io_out_valid, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  output [63:0] io_out_bits_cf_instr, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  output [38:0] io_out_bits_cf_pc, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  output [38:0] io_out_bits_cf_pnpc, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  output        io_out_bits_cf_intrVec_0, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  output        io_out_bits_cf_intrVec_1, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  output        io_out_bits_cf_intrVec_2, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  output        io_out_bits_cf_intrVec_3, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  output        io_out_bits_cf_intrVec_4, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  output        io_out_bits_cf_intrVec_5, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  output        io_out_bits_cf_intrVec_6, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  output        io_out_bits_cf_intrVec_7, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  output        io_out_bits_cf_intrVec_8, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  output        io_out_bits_cf_intrVec_9, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  output        io_out_bits_cf_intrVec_10, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  output        io_out_bits_cf_intrVec_11, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  input         DISPLAY_ENABLE,
  input  [11:0] intrVecIDU
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  reg [63:0] c; // @[src/main/scala/utils/GTimer.scala 24:20]
  wire [63:0] _c_T_1 = c + 64'h1; // @[src/main/scala/utils/GTimer.scala 25:12]
  wire  _T_214 = io_out_valid & DISPLAY_ENABLE; // @[src/main/scala/utils/Debug.scala 55:16]
  wire  _T_216 = ~reset; // @[src/main/scala/utils/Debug.scala 56:24]
  assign io_out_valid = 1'h0; // @[src/main/scala/nutcore/frontend/IDU.scala 161:16]
  assign io_out_bits_cf_instr = 64'h0; // @[src/main/scala/nutcore/frontend/IDU.scala 163:18]
  assign io_out_bits_cf_pc = 39'h0; // @[src/main/scala/nutcore/frontend/IDU.scala 163:18]
  assign io_out_bits_cf_pnpc = 39'h0; // @[src/main/scala/nutcore/frontend/IDU.scala 163:18]
  assign io_out_bits_cf_intrVec_0 = intrVecIDU[0]; // @[src/main/scala/nutcore/frontend/IDU.scala 171:38]
  assign io_out_bits_cf_intrVec_1 = intrVecIDU[1]; // @[src/main/scala/nutcore/frontend/IDU.scala 171:38]
  assign io_out_bits_cf_intrVec_2 = intrVecIDU[2]; // @[src/main/scala/nutcore/frontend/IDU.scala 171:38]
  assign io_out_bits_cf_intrVec_3 = intrVecIDU[3]; // @[src/main/scala/nutcore/frontend/IDU.scala 171:38]
  assign io_out_bits_cf_intrVec_4 = intrVecIDU[4]; // @[src/main/scala/nutcore/frontend/IDU.scala 171:38]
  assign io_out_bits_cf_intrVec_5 = intrVecIDU[5]; // @[src/main/scala/nutcore/frontend/IDU.scala 171:38]
  assign io_out_bits_cf_intrVec_6 = intrVecIDU[6]; // @[src/main/scala/nutcore/frontend/IDU.scala 171:38]
  assign io_out_bits_cf_intrVec_7 = intrVecIDU[7]; // @[src/main/scala/nutcore/frontend/IDU.scala 171:38]
  assign io_out_bits_cf_intrVec_8 = intrVecIDU[8]; // @[src/main/scala/nutcore/frontend/IDU.scala 171:38]
  assign io_out_bits_cf_intrVec_9 = intrVecIDU[9]; // @[src/main/scala/nutcore/frontend/IDU.scala 171:38]
  assign io_out_bits_cf_intrVec_10 = intrVecIDU[10]; // @[src/main/scala/nutcore/frontend/IDU.scala 171:38]
  assign io_out_bits_cf_intrVec_11 = intrVecIDU[11]; // @[src/main/scala/nutcore/frontend/IDU.scala 171:38]
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/utils/GTimer.scala 24:20]
      c <= 64'h0; // @[src/main/scala/utils/GTimer.scala 24:20]
    end else begin
      c <= _c_T_1; // @[src/main/scala/utils/GTimer.scala 25:7]
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_214 & ~reset) begin
          $fwrite(32'h80000002,"[%d] Decoder_1: ",c); // @[src/main/scala/utils/Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_214 & _T_216) begin
          $fwrite(32'h80000002,"issue: pc %x npc %x instr %x\n",io_out_bits_cf_pc,io_out_bits_cf_pnpc,
            io_out_bits_cf_instr); // @[src/main/scala/utils/Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  c = _RAND_0[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module IDU(
  input         clock,
  input         reset,
  output        io_in_0_ready, // @[src/main/scala/nutcore/frontend/IDU.scala 194:14]
  input         io_in_0_valid, // @[src/main/scala/nutcore/frontend/IDU.scala 194:14]
  input  [63:0] io_in_0_bits_instr, // @[src/main/scala/nutcore/frontend/IDU.scala 194:14]
  input  [38:0] io_in_0_bits_pc, // @[src/main/scala/nutcore/frontend/IDU.scala 194:14]
  input  [38:0] io_in_0_bits_pnpc, // @[src/main/scala/nutcore/frontend/IDU.scala 194:14]
  input         io_in_0_bits_exceptionVec_12, // @[src/main/scala/nutcore/frontend/IDU.scala 194:14]
  input  [3:0]  io_in_0_bits_brIdx, // @[src/main/scala/nutcore/frontend/IDU.scala 194:14]
  input         io_in_0_bits_crossPageIPFFix, // @[src/main/scala/nutcore/frontend/IDU.scala 194:14]
  input         io_out_0_ready, // @[src/main/scala/nutcore/frontend/IDU.scala 194:14]
  output        io_out_0_valid, // @[src/main/scala/nutcore/frontend/IDU.scala 194:14]
  output [63:0] io_out_0_bits_cf_instr, // @[src/main/scala/nutcore/frontend/IDU.scala 194:14]
  output [38:0] io_out_0_bits_cf_pc, // @[src/main/scala/nutcore/frontend/IDU.scala 194:14]
  output [38:0] io_out_0_bits_cf_pnpc, // @[src/main/scala/nutcore/frontend/IDU.scala 194:14]
  output        io_out_0_bits_cf_exceptionVec_1, // @[src/main/scala/nutcore/frontend/IDU.scala 194:14]
  output        io_out_0_bits_cf_exceptionVec_2, // @[src/main/scala/nutcore/frontend/IDU.scala 194:14]
  output        io_out_0_bits_cf_exceptionVec_12, // @[src/main/scala/nutcore/frontend/IDU.scala 194:14]
  output        io_out_0_bits_cf_intrVec_0, // @[src/main/scala/nutcore/frontend/IDU.scala 194:14]
  output        io_out_0_bits_cf_intrVec_1, // @[src/main/scala/nutcore/frontend/IDU.scala 194:14]
  output        io_out_0_bits_cf_intrVec_2, // @[src/main/scala/nutcore/frontend/IDU.scala 194:14]
  output        io_out_0_bits_cf_intrVec_3, // @[src/main/scala/nutcore/frontend/IDU.scala 194:14]
  output        io_out_0_bits_cf_intrVec_4, // @[src/main/scala/nutcore/frontend/IDU.scala 194:14]
  output        io_out_0_bits_cf_intrVec_5, // @[src/main/scala/nutcore/frontend/IDU.scala 194:14]
  output        io_out_0_bits_cf_intrVec_6, // @[src/main/scala/nutcore/frontend/IDU.scala 194:14]
  output        io_out_0_bits_cf_intrVec_7, // @[src/main/scala/nutcore/frontend/IDU.scala 194:14]
  output        io_out_0_bits_cf_intrVec_8, // @[src/main/scala/nutcore/frontend/IDU.scala 194:14]
  output        io_out_0_bits_cf_intrVec_9, // @[src/main/scala/nutcore/frontend/IDU.scala 194:14]
  output        io_out_0_bits_cf_intrVec_10, // @[src/main/scala/nutcore/frontend/IDU.scala 194:14]
  output        io_out_0_bits_cf_intrVec_11, // @[src/main/scala/nutcore/frontend/IDU.scala 194:14]
  output [3:0]  io_out_0_bits_cf_brIdx, // @[src/main/scala/nutcore/frontend/IDU.scala 194:14]
  output        io_out_0_bits_cf_crossPageIPFFix, // @[src/main/scala/nutcore/frontend/IDU.scala 194:14]
  output        io_out_0_bits_ctrl_src1Type, // @[src/main/scala/nutcore/frontend/IDU.scala 194:14]
  output        io_out_0_bits_ctrl_src2Type, // @[src/main/scala/nutcore/frontend/IDU.scala 194:14]
  output [2:0]  io_out_0_bits_ctrl_fuType, // @[src/main/scala/nutcore/frontend/IDU.scala 194:14]
  output [6:0]  io_out_0_bits_ctrl_fuOpType, // @[src/main/scala/nutcore/frontend/IDU.scala 194:14]
  output [4:0]  io_out_0_bits_ctrl_rfSrc1, // @[src/main/scala/nutcore/frontend/IDU.scala 194:14]
  output [4:0]  io_out_0_bits_ctrl_rfSrc2, // @[src/main/scala/nutcore/frontend/IDU.scala 194:14]
  output        io_out_0_bits_ctrl_rfWen, // @[src/main/scala/nutcore/frontend/IDU.scala 194:14]
  output [4:0]  io_out_0_bits_ctrl_rfDest, // @[src/main/scala/nutcore/frontend/IDU.scala 194:14]
  output        io_out_0_bits_ctrl_isNutCoreTrap, // @[src/main/scala/nutcore/frontend/IDU.scala 194:14]
  output [63:0] io_out_0_bits_data_imm, // @[src/main/scala/nutcore/frontend/IDU.scala 194:14]
  output        io_out_1_bits_cf_intrVec_0, // @[src/main/scala/nutcore/frontend/IDU.scala 194:14]
  output        io_out_1_bits_cf_intrVec_1, // @[src/main/scala/nutcore/frontend/IDU.scala 194:14]
  output        io_out_1_bits_cf_intrVec_2, // @[src/main/scala/nutcore/frontend/IDU.scala 194:14]
  output        io_out_1_bits_cf_intrVec_3, // @[src/main/scala/nutcore/frontend/IDU.scala 194:14]
  output        io_out_1_bits_cf_intrVec_4, // @[src/main/scala/nutcore/frontend/IDU.scala 194:14]
  output        io_out_1_bits_cf_intrVec_5, // @[src/main/scala/nutcore/frontend/IDU.scala 194:14]
  output        io_out_1_bits_cf_intrVec_6, // @[src/main/scala/nutcore/frontend/IDU.scala 194:14]
  output        io_out_1_bits_cf_intrVec_7, // @[src/main/scala/nutcore/frontend/IDU.scala 194:14]
  output        io_out_1_bits_cf_intrVec_8, // @[src/main/scala/nutcore/frontend/IDU.scala 194:14]
  output        io_out_1_bits_cf_intrVec_9, // @[src/main/scala/nutcore/frontend/IDU.scala 194:14]
  output        io_out_1_bits_cf_intrVec_10, // @[src/main/scala/nutcore/frontend/IDU.scala 194:14]
  output        io_out_1_bits_cf_intrVec_11, // @[src/main/scala/nutcore/frontend/IDU.scala 194:14]
  output        _WIRE_1,
  input         _WIRE_5,
  input  [11:0] _WIRE_14,
  input         _WIRE_2_2
);
  wire  decoder1_clock; // @[src/main/scala/nutcore/frontend/IDU.scala 198:25]
  wire  decoder1_reset; // @[src/main/scala/nutcore/frontend/IDU.scala 198:25]
  wire  decoder1_io_in_ready; // @[src/main/scala/nutcore/frontend/IDU.scala 198:25]
  wire  decoder1_io_in_valid; // @[src/main/scala/nutcore/frontend/IDU.scala 198:25]
  wire [63:0] decoder1_io_in_bits_instr; // @[src/main/scala/nutcore/frontend/IDU.scala 198:25]
  wire [38:0] decoder1_io_in_bits_pc; // @[src/main/scala/nutcore/frontend/IDU.scala 198:25]
  wire [38:0] decoder1_io_in_bits_pnpc; // @[src/main/scala/nutcore/frontend/IDU.scala 198:25]
  wire  decoder1_io_in_bits_exceptionVec_12; // @[src/main/scala/nutcore/frontend/IDU.scala 198:25]
  wire [3:0] decoder1_io_in_bits_brIdx; // @[src/main/scala/nutcore/frontend/IDU.scala 198:25]
  wire  decoder1_io_in_bits_crossPageIPFFix; // @[src/main/scala/nutcore/frontend/IDU.scala 198:25]
  wire  decoder1_io_out_ready; // @[src/main/scala/nutcore/frontend/IDU.scala 198:25]
  wire  decoder1_io_out_valid; // @[src/main/scala/nutcore/frontend/IDU.scala 198:25]
  wire [63:0] decoder1_io_out_bits_cf_instr; // @[src/main/scala/nutcore/frontend/IDU.scala 198:25]
  wire [38:0] decoder1_io_out_bits_cf_pc; // @[src/main/scala/nutcore/frontend/IDU.scala 198:25]
  wire [38:0] decoder1_io_out_bits_cf_pnpc; // @[src/main/scala/nutcore/frontend/IDU.scala 198:25]
  wire  decoder1_io_out_bits_cf_exceptionVec_1; // @[src/main/scala/nutcore/frontend/IDU.scala 198:25]
  wire  decoder1_io_out_bits_cf_exceptionVec_2; // @[src/main/scala/nutcore/frontend/IDU.scala 198:25]
  wire  decoder1_io_out_bits_cf_exceptionVec_12; // @[src/main/scala/nutcore/frontend/IDU.scala 198:25]
  wire  decoder1_io_out_bits_cf_intrVec_0; // @[src/main/scala/nutcore/frontend/IDU.scala 198:25]
  wire  decoder1_io_out_bits_cf_intrVec_1; // @[src/main/scala/nutcore/frontend/IDU.scala 198:25]
  wire  decoder1_io_out_bits_cf_intrVec_2; // @[src/main/scala/nutcore/frontend/IDU.scala 198:25]
  wire  decoder1_io_out_bits_cf_intrVec_3; // @[src/main/scala/nutcore/frontend/IDU.scala 198:25]
  wire  decoder1_io_out_bits_cf_intrVec_4; // @[src/main/scala/nutcore/frontend/IDU.scala 198:25]
  wire  decoder1_io_out_bits_cf_intrVec_5; // @[src/main/scala/nutcore/frontend/IDU.scala 198:25]
  wire  decoder1_io_out_bits_cf_intrVec_6; // @[src/main/scala/nutcore/frontend/IDU.scala 198:25]
  wire  decoder1_io_out_bits_cf_intrVec_7; // @[src/main/scala/nutcore/frontend/IDU.scala 198:25]
  wire  decoder1_io_out_bits_cf_intrVec_8; // @[src/main/scala/nutcore/frontend/IDU.scala 198:25]
  wire  decoder1_io_out_bits_cf_intrVec_9; // @[src/main/scala/nutcore/frontend/IDU.scala 198:25]
  wire  decoder1_io_out_bits_cf_intrVec_10; // @[src/main/scala/nutcore/frontend/IDU.scala 198:25]
  wire  decoder1_io_out_bits_cf_intrVec_11; // @[src/main/scala/nutcore/frontend/IDU.scala 198:25]
  wire [3:0] decoder1_io_out_bits_cf_brIdx; // @[src/main/scala/nutcore/frontend/IDU.scala 198:25]
  wire  decoder1_io_out_bits_cf_crossPageIPFFix; // @[src/main/scala/nutcore/frontend/IDU.scala 198:25]
  wire  decoder1_io_out_bits_ctrl_src1Type; // @[src/main/scala/nutcore/frontend/IDU.scala 198:25]
  wire  decoder1_io_out_bits_ctrl_src2Type; // @[src/main/scala/nutcore/frontend/IDU.scala 198:25]
  wire [2:0] decoder1_io_out_bits_ctrl_fuType; // @[src/main/scala/nutcore/frontend/IDU.scala 198:25]
  wire [6:0] decoder1_io_out_bits_ctrl_fuOpType; // @[src/main/scala/nutcore/frontend/IDU.scala 198:25]
  wire [4:0] decoder1_io_out_bits_ctrl_rfSrc1; // @[src/main/scala/nutcore/frontend/IDU.scala 198:25]
  wire [4:0] decoder1_io_out_bits_ctrl_rfSrc2; // @[src/main/scala/nutcore/frontend/IDU.scala 198:25]
  wire  decoder1_io_out_bits_ctrl_rfWen; // @[src/main/scala/nutcore/frontend/IDU.scala 198:25]
  wire [4:0] decoder1_io_out_bits_ctrl_rfDest; // @[src/main/scala/nutcore/frontend/IDU.scala 198:25]
  wire  decoder1_io_out_bits_ctrl_isNutCoreTrap; // @[src/main/scala/nutcore/frontend/IDU.scala 198:25]
  wire [63:0] decoder1_io_out_bits_data_imm; // @[src/main/scala/nutcore/frontend/IDU.scala 198:25]
  wire  decoder1_io_isWFI; // @[src/main/scala/nutcore/frontend/IDU.scala 198:25]
  wire  decoder1_DISPLAY_ENABLE; // @[src/main/scala/nutcore/frontend/IDU.scala 198:25]
  wire [11:0] decoder1_intrVecIDU; // @[src/main/scala/nutcore/frontend/IDU.scala 198:25]
  wire  decoder1_DTLBENABLE; // @[src/main/scala/nutcore/frontend/IDU.scala 198:25]
  wire  decoder2_clock; // @[src/main/scala/nutcore/frontend/IDU.scala 199:25]
  wire  decoder2_reset; // @[src/main/scala/nutcore/frontend/IDU.scala 199:25]
  wire  decoder2_io_out_valid; // @[src/main/scala/nutcore/frontend/IDU.scala 199:25]
  wire [63:0] decoder2_io_out_bits_cf_instr; // @[src/main/scala/nutcore/frontend/IDU.scala 199:25]
  wire [38:0] decoder2_io_out_bits_cf_pc; // @[src/main/scala/nutcore/frontend/IDU.scala 199:25]
  wire [38:0] decoder2_io_out_bits_cf_pnpc; // @[src/main/scala/nutcore/frontend/IDU.scala 199:25]
  wire  decoder2_io_out_bits_cf_intrVec_0; // @[src/main/scala/nutcore/frontend/IDU.scala 199:25]
  wire  decoder2_io_out_bits_cf_intrVec_1; // @[src/main/scala/nutcore/frontend/IDU.scala 199:25]
  wire  decoder2_io_out_bits_cf_intrVec_2; // @[src/main/scala/nutcore/frontend/IDU.scala 199:25]
  wire  decoder2_io_out_bits_cf_intrVec_3; // @[src/main/scala/nutcore/frontend/IDU.scala 199:25]
  wire  decoder2_io_out_bits_cf_intrVec_4; // @[src/main/scala/nutcore/frontend/IDU.scala 199:25]
  wire  decoder2_io_out_bits_cf_intrVec_5; // @[src/main/scala/nutcore/frontend/IDU.scala 199:25]
  wire  decoder2_io_out_bits_cf_intrVec_6; // @[src/main/scala/nutcore/frontend/IDU.scala 199:25]
  wire  decoder2_io_out_bits_cf_intrVec_7; // @[src/main/scala/nutcore/frontend/IDU.scala 199:25]
  wire  decoder2_io_out_bits_cf_intrVec_8; // @[src/main/scala/nutcore/frontend/IDU.scala 199:25]
  wire  decoder2_io_out_bits_cf_intrVec_9; // @[src/main/scala/nutcore/frontend/IDU.scala 199:25]
  wire  decoder2_io_out_bits_cf_intrVec_10; // @[src/main/scala/nutcore/frontend/IDU.scala 199:25]
  wire  decoder2_io_out_bits_cf_intrVec_11; // @[src/main/scala/nutcore/frontend/IDU.scala 199:25]
  wire  decoder2_DISPLAY_ENABLE; // @[src/main/scala/nutcore/frontend/IDU.scala 199:25]
  wire [11:0] decoder2_intrVecIDU; // @[src/main/scala/nutcore/frontend/IDU.scala 199:25]
  wire  _WIRE = decoder1_io_isWFI; // @[src/main/scala/nutcore/frontend/IDU.scala 219:54]
  Decoder decoder1 ( // @[src/main/scala/nutcore/frontend/IDU.scala 198:25]
    .clock(decoder1_clock),
    .reset(decoder1_reset),
    .io_in_ready(decoder1_io_in_ready),
    .io_in_valid(decoder1_io_in_valid),
    .io_in_bits_instr(decoder1_io_in_bits_instr),
    .io_in_bits_pc(decoder1_io_in_bits_pc),
    .io_in_bits_pnpc(decoder1_io_in_bits_pnpc),
    .io_in_bits_exceptionVec_12(decoder1_io_in_bits_exceptionVec_12),
    .io_in_bits_brIdx(decoder1_io_in_bits_brIdx),
    .io_in_bits_crossPageIPFFix(decoder1_io_in_bits_crossPageIPFFix),
    .io_out_ready(decoder1_io_out_ready),
    .io_out_valid(decoder1_io_out_valid),
    .io_out_bits_cf_instr(decoder1_io_out_bits_cf_instr),
    .io_out_bits_cf_pc(decoder1_io_out_bits_cf_pc),
    .io_out_bits_cf_pnpc(decoder1_io_out_bits_cf_pnpc),
    .io_out_bits_cf_exceptionVec_1(decoder1_io_out_bits_cf_exceptionVec_1),
    .io_out_bits_cf_exceptionVec_2(decoder1_io_out_bits_cf_exceptionVec_2),
    .io_out_bits_cf_exceptionVec_12(decoder1_io_out_bits_cf_exceptionVec_12),
    .io_out_bits_cf_intrVec_0(decoder1_io_out_bits_cf_intrVec_0),
    .io_out_bits_cf_intrVec_1(decoder1_io_out_bits_cf_intrVec_1),
    .io_out_bits_cf_intrVec_2(decoder1_io_out_bits_cf_intrVec_2),
    .io_out_bits_cf_intrVec_3(decoder1_io_out_bits_cf_intrVec_3),
    .io_out_bits_cf_intrVec_4(decoder1_io_out_bits_cf_intrVec_4),
    .io_out_bits_cf_intrVec_5(decoder1_io_out_bits_cf_intrVec_5),
    .io_out_bits_cf_intrVec_6(decoder1_io_out_bits_cf_intrVec_6),
    .io_out_bits_cf_intrVec_7(decoder1_io_out_bits_cf_intrVec_7),
    .io_out_bits_cf_intrVec_8(decoder1_io_out_bits_cf_intrVec_8),
    .io_out_bits_cf_intrVec_9(decoder1_io_out_bits_cf_intrVec_9),
    .io_out_bits_cf_intrVec_10(decoder1_io_out_bits_cf_intrVec_10),
    .io_out_bits_cf_intrVec_11(decoder1_io_out_bits_cf_intrVec_11),
    .io_out_bits_cf_brIdx(decoder1_io_out_bits_cf_brIdx),
    .io_out_bits_cf_crossPageIPFFix(decoder1_io_out_bits_cf_crossPageIPFFix),
    .io_out_bits_ctrl_src1Type(decoder1_io_out_bits_ctrl_src1Type),
    .io_out_bits_ctrl_src2Type(decoder1_io_out_bits_ctrl_src2Type),
    .io_out_bits_ctrl_fuType(decoder1_io_out_bits_ctrl_fuType),
    .io_out_bits_ctrl_fuOpType(decoder1_io_out_bits_ctrl_fuOpType),
    .io_out_bits_ctrl_rfSrc1(decoder1_io_out_bits_ctrl_rfSrc1),
    .io_out_bits_ctrl_rfSrc2(decoder1_io_out_bits_ctrl_rfSrc2),
    .io_out_bits_ctrl_rfWen(decoder1_io_out_bits_ctrl_rfWen),
    .io_out_bits_ctrl_rfDest(decoder1_io_out_bits_ctrl_rfDest),
    .io_out_bits_ctrl_isNutCoreTrap(decoder1_io_out_bits_ctrl_isNutCoreTrap),
    .io_out_bits_data_imm(decoder1_io_out_bits_data_imm),
    .io_isWFI(decoder1_io_isWFI),
    .DISPLAY_ENABLE(decoder1_DISPLAY_ENABLE),
    .intrVecIDU(decoder1_intrVecIDU),
    .DTLBENABLE(decoder1_DTLBENABLE)
  );
  Decoder_1 decoder2 ( // @[src/main/scala/nutcore/frontend/IDU.scala 199:25]
    .clock(decoder2_clock),
    .reset(decoder2_reset),
    .io_out_valid(decoder2_io_out_valid),
    .io_out_bits_cf_instr(decoder2_io_out_bits_cf_instr),
    .io_out_bits_cf_pc(decoder2_io_out_bits_cf_pc),
    .io_out_bits_cf_pnpc(decoder2_io_out_bits_cf_pnpc),
    .io_out_bits_cf_intrVec_0(decoder2_io_out_bits_cf_intrVec_0),
    .io_out_bits_cf_intrVec_1(decoder2_io_out_bits_cf_intrVec_1),
    .io_out_bits_cf_intrVec_2(decoder2_io_out_bits_cf_intrVec_2),
    .io_out_bits_cf_intrVec_3(decoder2_io_out_bits_cf_intrVec_3),
    .io_out_bits_cf_intrVec_4(decoder2_io_out_bits_cf_intrVec_4),
    .io_out_bits_cf_intrVec_5(decoder2_io_out_bits_cf_intrVec_5),
    .io_out_bits_cf_intrVec_6(decoder2_io_out_bits_cf_intrVec_6),
    .io_out_bits_cf_intrVec_7(decoder2_io_out_bits_cf_intrVec_7),
    .io_out_bits_cf_intrVec_8(decoder2_io_out_bits_cf_intrVec_8),
    .io_out_bits_cf_intrVec_9(decoder2_io_out_bits_cf_intrVec_9),
    .io_out_bits_cf_intrVec_10(decoder2_io_out_bits_cf_intrVec_10),
    .io_out_bits_cf_intrVec_11(decoder2_io_out_bits_cf_intrVec_11),
    .DISPLAY_ENABLE(decoder2_DISPLAY_ENABLE),
    .intrVecIDU(decoder2_intrVecIDU)
  );
  assign io_in_0_ready = decoder1_io_in_ready; // @[src/main/scala/nutcore/frontend/IDU.scala 200:12]
  assign io_out_0_valid = decoder1_io_out_valid; // @[src/main/scala/nutcore/frontend/IDU.scala 202:13]
  assign io_out_0_bits_cf_instr = decoder1_io_out_bits_cf_instr; // @[src/main/scala/nutcore/frontend/IDU.scala 202:13]
  assign io_out_0_bits_cf_pc = decoder1_io_out_bits_cf_pc; // @[src/main/scala/nutcore/frontend/IDU.scala 202:13]
  assign io_out_0_bits_cf_pnpc = decoder1_io_out_bits_cf_pnpc; // @[src/main/scala/nutcore/frontend/IDU.scala 202:13]
  assign io_out_0_bits_cf_exceptionVec_1 = decoder1_io_out_bits_cf_exceptionVec_1; // @[src/main/scala/nutcore/frontend/IDU.scala 202:13]
  assign io_out_0_bits_cf_exceptionVec_2 = decoder1_io_out_bits_cf_exceptionVec_2; // @[src/main/scala/nutcore/frontend/IDU.scala 202:13]
  assign io_out_0_bits_cf_exceptionVec_12 = decoder1_io_out_bits_cf_exceptionVec_12; // @[src/main/scala/nutcore/frontend/IDU.scala 202:13]
  assign io_out_0_bits_cf_intrVec_0 = decoder1_io_out_bits_cf_intrVec_0; // @[src/main/scala/nutcore/frontend/IDU.scala 202:13]
  assign io_out_0_bits_cf_intrVec_1 = decoder1_io_out_bits_cf_intrVec_1; // @[src/main/scala/nutcore/frontend/IDU.scala 202:13]
  assign io_out_0_bits_cf_intrVec_2 = decoder1_io_out_bits_cf_intrVec_2; // @[src/main/scala/nutcore/frontend/IDU.scala 202:13]
  assign io_out_0_bits_cf_intrVec_3 = decoder1_io_out_bits_cf_intrVec_3; // @[src/main/scala/nutcore/frontend/IDU.scala 202:13]
  assign io_out_0_bits_cf_intrVec_4 = decoder1_io_out_bits_cf_intrVec_4; // @[src/main/scala/nutcore/frontend/IDU.scala 202:13]
  assign io_out_0_bits_cf_intrVec_5 = decoder1_io_out_bits_cf_intrVec_5; // @[src/main/scala/nutcore/frontend/IDU.scala 202:13]
  assign io_out_0_bits_cf_intrVec_6 = decoder1_io_out_bits_cf_intrVec_6; // @[src/main/scala/nutcore/frontend/IDU.scala 202:13]
  assign io_out_0_bits_cf_intrVec_7 = decoder1_io_out_bits_cf_intrVec_7; // @[src/main/scala/nutcore/frontend/IDU.scala 202:13]
  assign io_out_0_bits_cf_intrVec_8 = decoder1_io_out_bits_cf_intrVec_8; // @[src/main/scala/nutcore/frontend/IDU.scala 202:13]
  assign io_out_0_bits_cf_intrVec_9 = decoder1_io_out_bits_cf_intrVec_9; // @[src/main/scala/nutcore/frontend/IDU.scala 202:13]
  assign io_out_0_bits_cf_intrVec_10 = decoder1_io_out_bits_cf_intrVec_10; // @[src/main/scala/nutcore/frontend/IDU.scala 202:13]
  assign io_out_0_bits_cf_intrVec_11 = decoder1_io_out_bits_cf_intrVec_11; // @[src/main/scala/nutcore/frontend/IDU.scala 202:13]
  assign io_out_0_bits_cf_brIdx = decoder1_io_out_bits_cf_brIdx; // @[src/main/scala/nutcore/frontend/IDU.scala 202:13]
  assign io_out_0_bits_cf_crossPageIPFFix = decoder1_io_out_bits_cf_crossPageIPFFix; // @[src/main/scala/nutcore/frontend/IDU.scala 202:13]
  assign io_out_0_bits_ctrl_src1Type = decoder1_io_out_bits_ctrl_src1Type; // @[src/main/scala/nutcore/frontend/IDU.scala 202:13]
  assign io_out_0_bits_ctrl_src2Type = decoder1_io_out_bits_ctrl_src2Type; // @[src/main/scala/nutcore/frontend/IDU.scala 202:13]
  assign io_out_0_bits_ctrl_fuType = decoder1_io_out_bits_ctrl_fuType; // @[src/main/scala/nutcore/frontend/IDU.scala 202:13]
  assign io_out_0_bits_ctrl_fuOpType = decoder1_io_out_bits_ctrl_fuOpType; // @[src/main/scala/nutcore/frontend/IDU.scala 202:13]
  assign io_out_0_bits_ctrl_rfSrc1 = decoder1_io_out_bits_ctrl_rfSrc1; // @[src/main/scala/nutcore/frontend/IDU.scala 202:13]
  assign io_out_0_bits_ctrl_rfSrc2 = decoder1_io_out_bits_ctrl_rfSrc2; // @[src/main/scala/nutcore/frontend/IDU.scala 202:13]
  assign io_out_0_bits_ctrl_rfWen = decoder1_io_out_bits_ctrl_rfWen; // @[src/main/scala/nutcore/frontend/IDU.scala 202:13]
  assign io_out_0_bits_ctrl_rfDest = decoder1_io_out_bits_ctrl_rfDest; // @[src/main/scala/nutcore/frontend/IDU.scala 202:13]
  assign io_out_0_bits_ctrl_isNutCoreTrap = decoder1_io_out_bits_ctrl_isNutCoreTrap; // @[src/main/scala/nutcore/frontend/IDU.scala 202:13]
  assign io_out_0_bits_data_imm = decoder1_io_out_bits_data_imm; // @[src/main/scala/nutcore/frontend/IDU.scala 202:13]
  assign io_out_1_bits_cf_intrVec_0 = decoder2_io_out_bits_cf_intrVec_0; // @[src/main/scala/nutcore/frontend/IDU.scala 203:13]
  assign io_out_1_bits_cf_intrVec_1 = decoder2_io_out_bits_cf_intrVec_1; // @[src/main/scala/nutcore/frontend/IDU.scala 203:13]
  assign io_out_1_bits_cf_intrVec_2 = decoder2_io_out_bits_cf_intrVec_2; // @[src/main/scala/nutcore/frontend/IDU.scala 203:13]
  assign io_out_1_bits_cf_intrVec_3 = decoder2_io_out_bits_cf_intrVec_3; // @[src/main/scala/nutcore/frontend/IDU.scala 203:13]
  assign io_out_1_bits_cf_intrVec_4 = decoder2_io_out_bits_cf_intrVec_4; // @[src/main/scala/nutcore/frontend/IDU.scala 203:13]
  assign io_out_1_bits_cf_intrVec_5 = decoder2_io_out_bits_cf_intrVec_5; // @[src/main/scala/nutcore/frontend/IDU.scala 203:13]
  assign io_out_1_bits_cf_intrVec_6 = decoder2_io_out_bits_cf_intrVec_6; // @[src/main/scala/nutcore/frontend/IDU.scala 203:13]
  assign io_out_1_bits_cf_intrVec_7 = decoder2_io_out_bits_cf_intrVec_7; // @[src/main/scala/nutcore/frontend/IDU.scala 203:13]
  assign io_out_1_bits_cf_intrVec_8 = decoder2_io_out_bits_cf_intrVec_8; // @[src/main/scala/nutcore/frontend/IDU.scala 203:13]
  assign io_out_1_bits_cf_intrVec_9 = decoder2_io_out_bits_cf_intrVec_9; // @[src/main/scala/nutcore/frontend/IDU.scala 203:13]
  assign io_out_1_bits_cf_intrVec_10 = decoder2_io_out_bits_cf_intrVec_10; // @[src/main/scala/nutcore/frontend/IDU.scala 203:13]
  assign io_out_1_bits_cf_intrVec_11 = decoder2_io_out_bits_cf_intrVec_11; // @[src/main/scala/nutcore/frontend/IDU.scala 203:13]
  assign _WIRE_1 = _WIRE;
  assign decoder1_clock = clock;
  assign decoder1_reset = reset;
  assign decoder1_io_in_valid = io_in_0_valid; // @[src/main/scala/nutcore/frontend/IDU.scala 200:12]
  assign decoder1_io_in_bits_instr = io_in_0_bits_instr; // @[src/main/scala/nutcore/frontend/IDU.scala 200:12]
  assign decoder1_io_in_bits_pc = io_in_0_bits_pc; // @[src/main/scala/nutcore/frontend/IDU.scala 200:12]
  assign decoder1_io_in_bits_pnpc = io_in_0_bits_pnpc; // @[src/main/scala/nutcore/frontend/IDU.scala 200:12]
  assign decoder1_io_in_bits_exceptionVec_12 = io_in_0_bits_exceptionVec_12; // @[src/main/scala/nutcore/frontend/IDU.scala 200:12]
  assign decoder1_io_in_bits_brIdx = io_in_0_bits_brIdx; // @[src/main/scala/nutcore/frontend/IDU.scala 200:12]
  assign decoder1_io_in_bits_crossPageIPFFix = io_in_0_bits_crossPageIPFFix; // @[src/main/scala/nutcore/frontend/IDU.scala 200:12]
  assign decoder1_io_out_ready = io_out_0_ready; // @[src/main/scala/nutcore/frontend/IDU.scala 202:13]
  assign decoder1_DISPLAY_ENABLE = _WIRE_5;
  assign decoder1_intrVecIDU = _WIRE_14;
  assign decoder1_DTLBENABLE = _WIRE_2_2;
  assign decoder2_clock = clock;
  assign decoder2_reset = reset;
  assign decoder2_DISPLAY_ENABLE = _WIRE_5;
  assign decoder2_intrVecIDU = _WIRE_14;
endmodule
module FlushableQueue(
  input         clock,
  input         reset,
  output        io_enq_ready, // @[src/main/scala/utils/FlushableQueue.scala 21:14]
  input         io_enq_valid, // @[src/main/scala/utils/FlushableQueue.scala 21:14]
  input  [63:0] io_enq_bits_instr, // @[src/main/scala/utils/FlushableQueue.scala 21:14]
  input  [38:0] io_enq_bits_pc, // @[src/main/scala/utils/FlushableQueue.scala 21:14]
  input  [38:0] io_enq_bits_pnpc, // @[src/main/scala/utils/FlushableQueue.scala 21:14]
  input         io_enq_bits_exceptionVec_12, // @[src/main/scala/utils/FlushableQueue.scala 21:14]
  input  [3:0]  io_enq_bits_brIdx, // @[src/main/scala/utils/FlushableQueue.scala 21:14]
  input         io_deq_ready, // @[src/main/scala/utils/FlushableQueue.scala 21:14]
  output        io_deq_valid, // @[src/main/scala/utils/FlushableQueue.scala 21:14]
  output [63:0] io_deq_bits_instr, // @[src/main/scala/utils/FlushableQueue.scala 21:14]
  output [38:0] io_deq_bits_pc, // @[src/main/scala/utils/FlushableQueue.scala 21:14]
  output [38:0] io_deq_bits_pnpc, // @[src/main/scala/utils/FlushableQueue.scala 21:14]
  output        io_deq_bits_exceptionVec_12, // @[src/main/scala/utils/FlushableQueue.scala 21:14]
  output [3:0]  io_deq_bits_brIdx, // @[src/main/scala/utils/FlushableQueue.scala 21:14]
  input         io_flush // @[src/main/scala/utils/FlushableQueue.scala 21:14]
);
`ifdef RANDOMIZE_MEM_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
`endif // RANDOMIZE_REG_INIT
  reg [63:0] ram_instr [0:3]; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_instr_io_deq_bits_MPORT_en; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire [1:0] ram_instr_io_deq_bits_MPORT_addr; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire [63:0] ram_instr_io_deq_bits_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire [63:0] ram_instr_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire [1:0] ram_instr_MPORT_addr; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_instr_MPORT_mask; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_instr_MPORT_en; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  reg [38:0] ram_pc [0:3]; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_pc_io_deq_bits_MPORT_en; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire [1:0] ram_pc_io_deq_bits_MPORT_addr; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire [38:0] ram_pc_io_deq_bits_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire [38:0] ram_pc_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire [1:0] ram_pc_MPORT_addr; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_pc_MPORT_mask; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_pc_MPORT_en; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  reg [38:0] ram_pnpc [0:3]; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_pnpc_io_deq_bits_MPORT_en; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire [1:0] ram_pnpc_io_deq_bits_MPORT_addr; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire [38:0] ram_pnpc_io_deq_bits_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire [38:0] ram_pnpc_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire [1:0] ram_pnpc_MPORT_addr; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_pnpc_MPORT_mask; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_pnpc_MPORT_en; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  reg  ram_exceptionVec_12 [0:3]; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_12_io_deq_bits_MPORT_en; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire [1:0] ram_exceptionVec_12_io_deq_bits_MPORT_addr; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_12_io_deq_bits_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_12_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire [1:0] ram_exceptionVec_12_MPORT_addr; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_12_MPORT_mask; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_12_MPORT_en; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  reg [3:0] ram_brIdx [0:3]; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_brIdx_io_deq_bits_MPORT_en; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire [1:0] ram_brIdx_io_deq_bits_MPORT_addr; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire [3:0] ram_brIdx_io_deq_bits_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire [3:0] ram_brIdx_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire [1:0] ram_brIdx_MPORT_addr; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_brIdx_MPORT_mask; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_brIdx_MPORT_en; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  reg [1:0] enq_ptr_value; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
  reg [1:0] deq_ptr_value; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
  reg  maybe_full; // @[src/main/scala/utils/FlushableQueue.scala 26:35]
  wire  ptr_match = enq_ptr_value == deq_ptr_value; // @[src/main/scala/utils/FlushableQueue.scala 28:41]
  wire  empty = ptr_match & ~maybe_full; // @[src/main/scala/utils/FlushableQueue.scala 29:33]
  wire  full = ptr_match & maybe_full; // @[src/main/scala/utils/FlushableQueue.scala 30:32]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  wire [1:0] _value_T_1 = enq_ptr_value + 2'h1; // @[src/main/scala/chisel3/util/Counter.scala 77:24]
  wire [1:0] _value_T_3 = deq_ptr_value + 2'h1; // @[src/main/scala/chisel3/util/Counter.scala 77:24]
  assign ram_instr_io_deq_bits_MPORT_en = 1'h1;
  assign ram_instr_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_instr_io_deq_bits_MPORT_data = ram_instr[ram_instr_io_deq_bits_MPORT_addr]; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  assign ram_instr_MPORT_data = io_enq_bits_instr;
  assign ram_instr_MPORT_addr = enq_ptr_value;
  assign ram_instr_MPORT_mask = 1'h1;
  assign ram_instr_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_pc_io_deq_bits_MPORT_en = 1'h1;
  assign ram_pc_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_pc_io_deq_bits_MPORT_data = ram_pc[ram_pc_io_deq_bits_MPORT_addr]; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  assign ram_pc_MPORT_data = io_enq_bits_pc;
  assign ram_pc_MPORT_addr = enq_ptr_value;
  assign ram_pc_MPORT_mask = 1'h1;
  assign ram_pc_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_pnpc_io_deq_bits_MPORT_en = 1'h1;
  assign ram_pnpc_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_pnpc_io_deq_bits_MPORT_data = ram_pnpc[ram_pnpc_io_deq_bits_MPORT_addr]; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  assign ram_pnpc_MPORT_data = io_enq_bits_pnpc;
  assign ram_pnpc_MPORT_addr = enq_ptr_value;
  assign ram_pnpc_MPORT_mask = 1'h1;
  assign ram_pnpc_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_exceptionVec_12_io_deq_bits_MPORT_en = 1'h1;
  assign ram_exceptionVec_12_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_exceptionVec_12_io_deq_bits_MPORT_data = ram_exceptionVec_12[ram_exceptionVec_12_io_deq_bits_MPORT_addr]; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  assign ram_exceptionVec_12_MPORT_data = io_enq_bits_exceptionVec_12;
  assign ram_exceptionVec_12_MPORT_addr = enq_ptr_value;
  assign ram_exceptionVec_12_MPORT_mask = 1'h1;
  assign ram_exceptionVec_12_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_brIdx_io_deq_bits_MPORT_en = 1'h1;
  assign ram_brIdx_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_brIdx_io_deq_bits_MPORT_data = ram_brIdx[ram_brIdx_io_deq_bits_MPORT_addr]; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  assign ram_brIdx_MPORT_data = io_enq_bits_brIdx;
  assign ram_brIdx_MPORT_addr = enq_ptr_value;
  assign ram_brIdx_MPORT_mask = 1'h1;
  assign ram_brIdx_MPORT_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = ~full; // @[src/main/scala/utils/FlushableQueue.scala 46:19]
  assign io_deq_valid = ~empty; // @[src/main/scala/utils/FlushableQueue.scala 45:19]
  assign io_deq_bits_instr = ram_instr_io_deq_bits_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 47:15]
  assign io_deq_bits_pc = ram_pc_io_deq_bits_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 47:15]
  assign io_deq_bits_pnpc = ram_pnpc_io_deq_bits_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 47:15]
  assign io_deq_bits_exceptionVec_12 = ram_exceptionVec_12_io_deq_bits_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 47:15]
  assign io_deq_bits_brIdx = ram_brIdx_io_deq_bits_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 47:15]
  always @(posedge clock) begin
    if (ram_instr_MPORT_en & ram_instr_MPORT_mask) begin
      ram_instr[ram_instr_MPORT_addr] <= ram_instr_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
    end
    if (ram_pc_MPORT_en & ram_pc_MPORT_mask) begin
      ram_pc[ram_pc_MPORT_addr] <= ram_pc_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
    end
    if (ram_pnpc_MPORT_en & ram_pnpc_MPORT_mask) begin
      ram_pnpc[ram_pnpc_MPORT_addr] <= ram_pnpc_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
    end
    if (ram_exceptionVec_12_MPORT_en & ram_exceptionVec_12_MPORT_mask) begin
      ram_exceptionVec_12[ram_exceptionVec_12_MPORT_addr] <= ram_exceptionVec_12_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
    end
    if (ram_brIdx_MPORT_en & ram_brIdx_MPORT_mask) begin
      ram_brIdx[ram_brIdx_MPORT_addr] <= ram_brIdx_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
    end
    if (reset) begin // @[src/main/scala/chisel3/util/Counter.scala 61:40]
      enq_ptr_value <= 2'h0; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end else if (io_flush) begin // @[src/main/scala/utils/FlushableQueue.scala 62:19]
      enq_ptr_value <= 2'h0; // @[src/main/scala/utils/FlushableQueue.scala 64:21]
    end else if (do_enq) begin // @[src/main/scala/utils/FlushableQueue.scala 34:17]
      enq_ptr_value <= _value_T_1; // @[src/main/scala/chisel3/util/Counter.scala 77:15]
    end
    if (reset) begin // @[src/main/scala/chisel3/util/Counter.scala 61:40]
      deq_ptr_value <= 2'h0; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end else if (io_flush) begin // @[src/main/scala/utils/FlushableQueue.scala 62:19]
      deq_ptr_value <= 2'h0; // @[src/main/scala/utils/FlushableQueue.scala 65:21]
    end else if (do_deq) begin // @[src/main/scala/utils/FlushableQueue.scala 38:17]
      deq_ptr_value <= _value_T_3; // @[src/main/scala/chisel3/util/Counter.scala 77:15]
    end
    if (reset) begin // @[src/main/scala/utils/FlushableQueue.scala 26:35]
      maybe_full <= 1'h0; // @[src/main/scala/utils/FlushableQueue.scala 26:35]
    end else if (io_flush) begin // @[src/main/scala/utils/FlushableQueue.scala 62:19]
      maybe_full <= 1'h0; // @[src/main/scala/utils/FlushableQueue.scala 67:16]
    end else if (do_enq != do_deq) begin // @[src/main/scala/utils/FlushableQueue.scala 41:28]
      maybe_full <= do_enq; // @[src/main/scala/utils/FlushableQueue.scala 42:16]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {2{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    ram_instr[initvar] = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    ram_pc[initvar] = _RAND_1[38:0];
  _RAND_2 = {2{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    ram_pnpc[initvar] = _RAND_2[38:0];
  _RAND_3 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    ram_exceptionVec_12[initvar] = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    ram_brIdx[initvar] = _RAND_4[3:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  enq_ptr_value = _RAND_5[1:0];
  _RAND_6 = {1{`RANDOM}};
  deq_ptr_value = _RAND_6[1:0];
  _RAND_7 = {1{`RANDOM}};
  maybe_full = _RAND_7[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Frontend_inorder(
  input         clock,
  input         reset,
  input         io_imem_req_ready, // @[src/main/scala/nutcore/frontend/Frontend.scala 36:14]
  output        io_imem_req_valid, // @[src/main/scala/nutcore/frontend/Frontend.scala 36:14]
  output [38:0] io_imem_req_bits_addr, // @[src/main/scala/nutcore/frontend/Frontend.scala 36:14]
  output [86:0] io_imem_req_bits_user, // @[src/main/scala/nutcore/frontend/Frontend.scala 36:14]
  output        io_imem_resp_ready, // @[src/main/scala/nutcore/frontend/Frontend.scala 36:14]
  input         io_imem_resp_valid, // @[src/main/scala/nutcore/frontend/Frontend.scala 36:14]
  input  [63:0] io_imem_resp_bits_rdata, // @[src/main/scala/nutcore/frontend/Frontend.scala 36:14]
  input  [86:0] io_imem_resp_bits_user, // @[src/main/scala/nutcore/frontend/Frontend.scala 36:14]
  input         io_out_0_ready, // @[src/main/scala/nutcore/frontend/Frontend.scala 36:14]
  output        io_out_0_valid, // @[src/main/scala/nutcore/frontend/Frontend.scala 36:14]
  output [63:0] io_out_0_bits_cf_instr, // @[src/main/scala/nutcore/frontend/Frontend.scala 36:14]
  output [38:0] io_out_0_bits_cf_pc, // @[src/main/scala/nutcore/frontend/Frontend.scala 36:14]
  output [38:0] io_out_0_bits_cf_pnpc, // @[src/main/scala/nutcore/frontend/Frontend.scala 36:14]
  output        io_out_0_bits_cf_exceptionVec_1, // @[src/main/scala/nutcore/frontend/Frontend.scala 36:14]
  output        io_out_0_bits_cf_exceptionVec_2, // @[src/main/scala/nutcore/frontend/Frontend.scala 36:14]
  output        io_out_0_bits_cf_exceptionVec_12, // @[src/main/scala/nutcore/frontend/Frontend.scala 36:14]
  output        io_out_0_bits_cf_intrVec_0, // @[src/main/scala/nutcore/frontend/Frontend.scala 36:14]
  output        io_out_0_bits_cf_intrVec_1, // @[src/main/scala/nutcore/frontend/Frontend.scala 36:14]
  output        io_out_0_bits_cf_intrVec_2, // @[src/main/scala/nutcore/frontend/Frontend.scala 36:14]
  output        io_out_0_bits_cf_intrVec_3, // @[src/main/scala/nutcore/frontend/Frontend.scala 36:14]
  output        io_out_0_bits_cf_intrVec_4, // @[src/main/scala/nutcore/frontend/Frontend.scala 36:14]
  output        io_out_0_bits_cf_intrVec_5, // @[src/main/scala/nutcore/frontend/Frontend.scala 36:14]
  output        io_out_0_bits_cf_intrVec_6, // @[src/main/scala/nutcore/frontend/Frontend.scala 36:14]
  output        io_out_0_bits_cf_intrVec_7, // @[src/main/scala/nutcore/frontend/Frontend.scala 36:14]
  output        io_out_0_bits_cf_intrVec_8, // @[src/main/scala/nutcore/frontend/Frontend.scala 36:14]
  output        io_out_0_bits_cf_intrVec_9, // @[src/main/scala/nutcore/frontend/Frontend.scala 36:14]
  output        io_out_0_bits_cf_intrVec_10, // @[src/main/scala/nutcore/frontend/Frontend.scala 36:14]
  output        io_out_0_bits_cf_intrVec_11, // @[src/main/scala/nutcore/frontend/Frontend.scala 36:14]
  output [3:0]  io_out_0_bits_cf_brIdx, // @[src/main/scala/nutcore/frontend/Frontend.scala 36:14]
  output        io_out_0_bits_cf_crossPageIPFFix, // @[src/main/scala/nutcore/frontend/Frontend.scala 36:14]
  output        io_out_0_bits_ctrl_src1Type, // @[src/main/scala/nutcore/frontend/Frontend.scala 36:14]
  output        io_out_0_bits_ctrl_src2Type, // @[src/main/scala/nutcore/frontend/Frontend.scala 36:14]
  output [2:0]  io_out_0_bits_ctrl_fuType, // @[src/main/scala/nutcore/frontend/Frontend.scala 36:14]
  output [6:0]  io_out_0_bits_ctrl_fuOpType, // @[src/main/scala/nutcore/frontend/Frontend.scala 36:14]
  output [4:0]  io_out_0_bits_ctrl_rfSrc1, // @[src/main/scala/nutcore/frontend/Frontend.scala 36:14]
  output [4:0]  io_out_0_bits_ctrl_rfSrc2, // @[src/main/scala/nutcore/frontend/Frontend.scala 36:14]
  output        io_out_0_bits_ctrl_rfWen, // @[src/main/scala/nutcore/frontend/Frontend.scala 36:14]
  output [4:0]  io_out_0_bits_ctrl_rfDest, // @[src/main/scala/nutcore/frontend/Frontend.scala 36:14]
  output        io_out_0_bits_ctrl_isNutCoreTrap, // @[src/main/scala/nutcore/frontend/Frontend.scala 36:14]
  output [63:0] io_out_0_bits_data_imm, // @[src/main/scala/nutcore/frontend/Frontend.scala 36:14]
  output        io_out_1_bits_cf_intrVec_0, // @[src/main/scala/nutcore/frontend/Frontend.scala 36:14]
  output        io_out_1_bits_cf_intrVec_1, // @[src/main/scala/nutcore/frontend/Frontend.scala 36:14]
  output        io_out_1_bits_cf_intrVec_2, // @[src/main/scala/nutcore/frontend/Frontend.scala 36:14]
  output        io_out_1_bits_cf_intrVec_3, // @[src/main/scala/nutcore/frontend/Frontend.scala 36:14]
  output        io_out_1_bits_cf_intrVec_4, // @[src/main/scala/nutcore/frontend/Frontend.scala 36:14]
  output        io_out_1_bits_cf_intrVec_5, // @[src/main/scala/nutcore/frontend/Frontend.scala 36:14]
  output        io_out_1_bits_cf_intrVec_6, // @[src/main/scala/nutcore/frontend/Frontend.scala 36:14]
  output        io_out_1_bits_cf_intrVec_7, // @[src/main/scala/nutcore/frontend/Frontend.scala 36:14]
  output        io_out_1_bits_cf_intrVec_8, // @[src/main/scala/nutcore/frontend/Frontend.scala 36:14]
  output        io_out_1_bits_cf_intrVec_9, // @[src/main/scala/nutcore/frontend/Frontend.scala 36:14]
  output        io_out_1_bits_cf_intrVec_10, // @[src/main/scala/nutcore/frontend/Frontend.scala 36:14]
  output        io_out_1_bits_cf_intrVec_11, // @[src/main/scala/nutcore/frontend/Frontend.scala 36:14]
  output [3:0]  io_flushVec, // @[src/main/scala/nutcore/frontend/Frontend.scala 36:14]
  input  [38:0] io_redirect_target, // @[src/main/scala/nutcore/frontend/Frontend.scala 36:14]
  input         io_redirect_valid, // @[src/main/scala/nutcore/frontend/Frontend.scala 36:14]
  input         io_ipf, // @[src/main/scala/nutcore/frontend/Frontend.scala 36:14]
  input         REG_valid,
  input  [38:0] REG_pc,
  input         REG_isMissPredict,
  input  [38:0] REG_actualTarget,
  input         REG_actualTaken,
  input  [6:0]  REG_fuOpType,
  input  [1:0]  REG_btbType,
  input         REG_isRVC,
  output        _WIRE_0,
  input         DISPLAY_ENABLE,
  output        _WIRE_7,
  input         _WIRE_11,
  input         _WIRE_1_4,
  input  [11:0] _WIRE_14,
  input         _WIRE_2_2,
  output        r_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [63:0] _RAND_10;
`endif // RANDOMIZE_REG_INIT
  wire  ifu_clock; // @[src/main/scala/nutcore/frontend/Frontend.scala 94:20]
  wire  ifu_reset; // @[src/main/scala/nutcore/frontend/Frontend.scala 94:20]
  wire  ifu_io_imem_req_ready; // @[src/main/scala/nutcore/frontend/Frontend.scala 94:20]
  wire  ifu_io_imem_req_valid; // @[src/main/scala/nutcore/frontend/Frontend.scala 94:20]
  wire [38:0] ifu_io_imem_req_bits_addr; // @[src/main/scala/nutcore/frontend/Frontend.scala 94:20]
  wire [81:0] ifu_io_imem_req_bits_user; // @[src/main/scala/nutcore/frontend/Frontend.scala 94:20]
  wire  ifu_io_imem_resp_ready; // @[src/main/scala/nutcore/frontend/Frontend.scala 94:20]
  wire  ifu_io_imem_resp_valid; // @[src/main/scala/nutcore/frontend/Frontend.scala 94:20]
  wire [63:0] ifu_io_imem_resp_bits_rdata; // @[src/main/scala/nutcore/frontend/Frontend.scala 94:20]
  wire [81:0] ifu_io_imem_resp_bits_user; // @[src/main/scala/nutcore/frontend/Frontend.scala 94:20]
  wire  ifu_io_out_ready; // @[src/main/scala/nutcore/frontend/Frontend.scala 94:20]
  wire  ifu_io_out_valid; // @[src/main/scala/nutcore/frontend/Frontend.scala 94:20]
  wire [63:0] ifu_io_out_bits_instr; // @[src/main/scala/nutcore/frontend/Frontend.scala 94:20]
  wire [38:0] ifu_io_out_bits_pc; // @[src/main/scala/nutcore/frontend/Frontend.scala 94:20]
  wire [38:0] ifu_io_out_bits_pnpc; // @[src/main/scala/nutcore/frontend/Frontend.scala 94:20]
  wire  ifu_io_out_bits_exceptionVec_12; // @[src/main/scala/nutcore/frontend/Frontend.scala 94:20]
  wire [3:0] ifu_io_out_bits_brIdx; // @[src/main/scala/nutcore/frontend/Frontend.scala 94:20]
  wire [38:0] ifu_io_redirect_target; // @[src/main/scala/nutcore/frontend/Frontend.scala 94:20]
  wire  ifu_io_redirect_valid; // @[src/main/scala/nutcore/frontend/Frontend.scala 94:20]
  wire [3:0] ifu_io_flushVec; // @[src/main/scala/nutcore/frontend/Frontend.scala 94:20]
  wire  ifu_io_ipf; // @[src/main/scala/nutcore/frontend/Frontend.scala 94:20]
  wire  ifu_REG_valid; // @[src/main/scala/nutcore/frontend/Frontend.scala 94:20]
  wire [38:0] ifu_REG_pc; // @[src/main/scala/nutcore/frontend/Frontend.scala 94:20]
  wire  ifu_REG_isMissPredict; // @[src/main/scala/nutcore/frontend/Frontend.scala 94:20]
  wire [38:0] ifu_REG_actualTarget; // @[src/main/scala/nutcore/frontend/Frontend.scala 94:20]
  wire  ifu_REG_actualTaken; // @[src/main/scala/nutcore/frontend/Frontend.scala 94:20]
  wire [6:0] ifu_REG_fuOpType; // @[src/main/scala/nutcore/frontend/Frontend.scala 94:20]
  wire [1:0] ifu_REG_btbType; // @[src/main/scala/nutcore/frontend/Frontend.scala 94:20]
  wire  ifu_REG_isRVC; // @[src/main/scala/nutcore/frontend/Frontend.scala 94:20]
  wire  ifu_DISPLAY_ENABLE; // @[src/main/scala/nutcore/frontend/Frontend.scala 94:20]
  wire  ifu__WIRE_7; // @[src/main/scala/nutcore/frontend/Frontend.scala 94:20]
  wire  ifu__WIRE_11; // @[src/main/scala/nutcore/frontend/Frontend.scala 94:20]
  wire  ifu__WIRE_1_4; // @[src/main/scala/nutcore/frontend/Frontend.scala 94:20]
  wire  ifu_r_2; // @[src/main/scala/nutcore/frontend/Frontend.scala 94:20]
  wire  ibf_clock; // @[src/main/scala/nutcore/frontend/Frontend.scala 95:19]
  wire  ibf_reset; // @[src/main/scala/nutcore/frontend/Frontend.scala 95:19]
  wire  ibf_io_in_ready; // @[src/main/scala/nutcore/frontend/Frontend.scala 95:19]
  wire  ibf_io_in_valid; // @[src/main/scala/nutcore/frontend/Frontend.scala 95:19]
  wire [63:0] ibf_io_in_bits_instr; // @[src/main/scala/nutcore/frontend/Frontend.scala 95:19]
  wire [38:0] ibf_io_in_bits_pc; // @[src/main/scala/nutcore/frontend/Frontend.scala 95:19]
  wire [38:0] ibf_io_in_bits_pnpc; // @[src/main/scala/nutcore/frontend/Frontend.scala 95:19]
  wire  ibf_io_in_bits_exceptionVec_12; // @[src/main/scala/nutcore/frontend/Frontend.scala 95:19]
  wire [3:0] ibf_io_in_bits_brIdx; // @[src/main/scala/nutcore/frontend/Frontend.scala 95:19]
  wire  ibf_io_out_ready; // @[src/main/scala/nutcore/frontend/Frontend.scala 95:19]
  wire  ibf_io_out_valid; // @[src/main/scala/nutcore/frontend/Frontend.scala 95:19]
  wire [63:0] ibf_io_out_bits_instr; // @[src/main/scala/nutcore/frontend/Frontend.scala 95:19]
  wire [38:0] ibf_io_out_bits_pc; // @[src/main/scala/nutcore/frontend/Frontend.scala 95:19]
  wire [38:0] ibf_io_out_bits_pnpc; // @[src/main/scala/nutcore/frontend/Frontend.scala 95:19]
  wire  ibf_io_out_bits_exceptionVec_12; // @[src/main/scala/nutcore/frontend/Frontend.scala 95:19]
  wire [3:0] ibf_io_out_bits_brIdx; // @[src/main/scala/nutcore/frontend/Frontend.scala 95:19]
  wire  ibf_io_out_bits_crossPageIPFFix; // @[src/main/scala/nutcore/frontend/Frontend.scala 95:19]
  wire  ibf_io_flush; // @[src/main/scala/nutcore/frontend/Frontend.scala 95:19]
  wire  ibf_DISPLAY_ENABLE; // @[src/main/scala/nutcore/frontend/Frontend.scala 95:19]
  wire  idu_clock; // @[src/main/scala/nutcore/frontend/Frontend.scala 96:20]
  wire  idu_reset; // @[src/main/scala/nutcore/frontend/Frontend.scala 96:20]
  wire  idu_io_in_0_ready; // @[src/main/scala/nutcore/frontend/Frontend.scala 96:20]
  wire  idu_io_in_0_valid; // @[src/main/scala/nutcore/frontend/Frontend.scala 96:20]
  wire [63:0] idu_io_in_0_bits_instr; // @[src/main/scala/nutcore/frontend/Frontend.scala 96:20]
  wire [38:0] idu_io_in_0_bits_pc; // @[src/main/scala/nutcore/frontend/Frontend.scala 96:20]
  wire [38:0] idu_io_in_0_bits_pnpc; // @[src/main/scala/nutcore/frontend/Frontend.scala 96:20]
  wire  idu_io_in_0_bits_exceptionVec_12; // @[src/main/scala/nutcore/frontend/Frontend.scala 96:20]
  wire [3:0] idu_io_in_0_bits_brIdx; // @[src/main/scala/nutcore/frontend/Frontend.scala 96:20]
  wire  idu_io_in_0_bits_crossPageIPFFix; // @[src/main/scala/nutcore/frontend/Frontend.scala 96:20]
  wire  idu_io_out_0_ready; // @[src/main/scala/nutcore/frontend/Frontend.scala 96:20]
  wire  idu_io_out_0_valid; // @[src/main/scala/nutcore/frontend/Frontend.scala 96:20]
  wire [63:0] idu_io_out_0_bits_cf_instr; // @[src/main/scala/nutcore/frontend/Frontend.scala 96:20]
  wire [38:0] idu_io_out_0_bits_cf_pc; // @[src/main/scala/nutcore/frontend/Frontend.scala 96:20]
  wire [38:0] idu_io_out_0_bits_cf_pnpc; // @[src/main/scala/nutcore/frontend/Frontend.scala 96:20]
  wire  idu_io_out_0_bits_cf_exceptionVec_1; // @[src/main/scala/nutcore/frontend/Frontend.scala 96:20]
  wire  idu_io_out_0_bits_cf_exceptionVec_2; // @[src/main/scala/nutcore/frontend/Frontend.scala 96:20]
  wire  idu_io_out_0_bits_cf_exceptionVec_12; // @[src/main/scala/nutcore/frontend/Frontend.scala 96:20]
  wire  idu_io_out_0_bits_cf_intrVec_0; // @[src/main/scala/nutcore/frontend/Frontend.scala 96:20]
  wire  idu_io_out_0_bits_cf_intrVec_1; // @[src/main/scala/nutcore/frontend/Frontend.scala 96:20]
  wire  idu_io_out_0_bits_cf_intrVec_2; // @[src/main/scala/nutcore/frontend/Frontend.scala 96:20]
  wire  idu_io_out_0_bits_cf_intrVec_3; // @[src/main/scala/nutcore/frontend/Frontend.scala 96:20]
  wire  idu_io_out_0_bits_cf_intrVec_4; // @[src/main/scala/nutcore/frontend/Frontend.scala 96:20]
  wire  idu_io_out_0_bits_cf_intrVec_5; // @[src/main/scala/nutcore/frontend/Frontend.scala 96:20]
  wire  idu_io_out_0_bits_cf_intrVec_6; // @[src/main/scala/nutcore/frontend/Frontend.scala 96:20]
  wire  idu_io_out_0_bits_cf_intrVec_7; // @[src/main/scala/nutcore/frontend/Frontend.scala 96:20]
  wire  idu_io_out_0_bits_cf_intrVec_8; // @[src/main/scala/nutcore/frontend/Frontend.scala 96:20]
  wire  idu_io_out_0_bits_cf_intrVec_9; // @[src/main/scala/nutcore/frontend/Frontend.scala 96:20]
  wire  idu_io_out_0_bits_cf_intrVec_10; // @[src/main/scala/nutcore/frontend/Frontend.scala 96:20]
  wire  idu_io_out_0_bits_cf_intrVec_11; // @[src/main/scala/nutcore/frontend/Frontend.scala 96:20]
  wire [3:0] idu_io_out_0_bits_cf_brIdx; // @[src/main/scala/nutcore/frontend/Frontend.scala 96:20]
  wire  idu_io_out_0_bits_cf_crossPageIPFFix; // @[src/main/scala/nutcore/frontend/Frontend.scala 96:20]
  wire  idu_io_out_0_bits_ctrl_src1Type; // @[src/main/scala/nutcore/frontend/Frontend.scala 96:20]
  wire  idu_io_out_0_bits_ctrl_src2Type; // @[src/main/scala/nutcore/frontend/Frontend.scala 96:20]
  wire [2:0] idu_io_out_0_bits_ctrl_fuType; // @[src/main/scala/nutcore/frontend/Frontend.scala 96:20]
  wire [6:0] idu_io_out_0_bits_ctrl_fuOpType; // @[src/main/scala/nutcore/frontend/Frontend.scala 96:20]
  wire [4:0] idu_io_out_0_bits_ctrl_rfSrc1; // @[src/main/scala/nutcore/frontend/Frontend.scala 96:20]
  wire [4:0] idu_io_out_0_bits_ctrl_rfSrc2; // @[src/main/scala/nutcore/frontend/Frontend.scala 96:20]
  wire  idu_io_out_0_bits_ctrl_rfWen; // @[src/main/scala/nutcore/frontend/Frontend.scala 96:20]
  wire [4:0] idu_io_out_0_bits_ctrl_rfDest; // @[src/main/scala/nutcore/frontend/Frontend.scala 96:20]
  wire  idu_io_out_0_bits_ctrl_isNutCoreTrap; // @[src/main/scala/nutcore/frontend/Frontend.scala 96:20]
  wire [63:0] idu_io_out_0_bits_data_imm; // @[src/main/scala/nutcore/frontend/Frontend.scala 96:20]
  wire  idu_io_out_1_bits_cf_intrVec_0; // @[src/main/scala/nutcore/frontend/Frontend.scala 96:20]
  wire  idu_io_out_1_bits_cf_intrVec_1; // @[src/main/scala/nutcore/frontend/Frontend.scala 96:20]
  wire  idu_io_out_1_bits_cf_intrVec_2; // @[src/main/scala/nutcore/frontend/Frontend.scala 96:20]
  wire  idu_io_out_1_bits_cf_intrVec_3; // @[src/main/scala/nutcore/frontend/Frontend.scala 96:20]
  wire  idu_io_out_1_bits_cf_intrVec_4; // @[src/main/scala/nutcore/frontend/Frontend.scala 96:20]
  wire  idu_io_out_1_bits_cf_intrVec_5; // @[src/main/scala/nutcore/frontend/Frontend.scala 96:20]
  wire  idu_io_out_1_bits_cf_intrVec_6; // @[src/main/scala/nutcore/frontend/Frontend.scala 96:20]
  wire  idu_io_out_1_bits_cf_intrVec_7; // @[src/main/scala/nutcore/frontend/Frontend.scala 96:20]
  wire  idu_io_out_1_bits_cf_intrVec_8; // @[src/main/scala/nutcore/frontend/Frontend.scala 96:20]
  wire  idu_io_out_1_bits_cf_intrVec_9; // @[src/main/scala/nutcore/frontend/Frontend.scala 96:20]
  wire  idu_io_out_1_bits_cf_intrVec_10; // @[src/main/scala/nutcore/frontend/Frontend.scala 96:20]
  wire  idu_io_out_1_bits_cf_intrVec_11; // @[src/main/scala/nutcore/frontend/Frontend.scala 96:20]
  wire  idu__WIRE_1; // @[src/main/scala/nutcore/frontend/Frontend.scala 96:20]
  wire  idu__WIRE_5; // @[src/main/scala/nutcore/frontend/Frontend.scala 96:20]
  wire [11:0] idu__WIRE_14; // @[src/main/scala/nutcore/frontend/Frontend.scala 96:20]
  wire  idu__WIRE_2_2; // @[src/main/scala/nutcore/frontend/Frontend.scala 96:20]
  wire  ibf_io_in_q_clock; // @[src/main/scala/utils/FlushableQueue.scala 94:21]
  wire  ibf_io_in_q_reset; // @[src/main/scala/utils/FlushableQueue.scala 94:21]
  wire  ibf_io_in_q_io_enq_ready; // @[src/main/scala/utils/FlushableQueue.scala 94:21]
  wire  ibf_io_in_q_io_enq_valid; // @[src/main/scala/utils/FlushableQueue.scala 94:21]
  wire [63:0] ibf_io_in_q_io_enq_bits_instr; // @[src/main/scala/utils/FlushableQueue.scala 94:21]
  wire [38:0] ibf_io_in_q_io_enq_bits_pc; // @[src/main/scala/utils/FlushableQueue.scala 94:21]
  wire [38:0] ibf_io_in_q_io_enq_bits_pnpc; // @[src/main/scala/utils/FlushableQueue.scala 94:21]
  wire  ibf_io_in_q_io_enq_bits_exceptionVec_12; // @[src/main/scala/utils/FlushableQueue.scala 94:21]
  wire [3:0] ibf_io_in_q_io_enq_bits_brIdx; // @[src/main/scala/utils/FlushableQueue.scala 94:21]
  wire  ibf_io_in_q_io_deq_ready; // @[src/main/scala/utils/FlushableQueue.scala 94:21]
  wire  ibf_io_in_q_io_deq_valid; // @[src/main/scala/utils/FlushableQueue.scala 94:21]
  wire [63:0] ibf_io_in_q_io_deq_bits_instr; // @[src/main/scala/utils/FlushableQueue.scala 94:21]
  wire [38:0] ibf_io_in_q_io_deq_bits_pc; // @[src/main/scala/utils/FlushableQueue.scala 94:21]
  wire [38:0] ibf_io_in_q_io_deq_bits_pnpc; // @[src/main/scala/utils/FlushableQueue.scala 94:21]
  wire  ibf_io_in_q_io_deq_bits_exceptionVec_12; // @[src/main/scala/utils/FlushableQueue.scala 94:21]
  wire [3:0] ibf_io_in_q_io_deq_bits_brIdx; // @[src/main/scala/utils/FlushableQueue.scala 94:21]
  wire  ibf_io_in_q_io_flush; // @[src/main/scala/utils/FlushableQueue.scala 94:21]
  wire  _T_1 = idu_io_out_0_ready & idu_io_out_0_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  reg  valid; // @[src/main/scala/utils/Pipeline.scala 24:24]
  wire  _GEN_0 = _T_1 ? 1'h0 : valid; // @[src/main/scala/utils/Pipeline.scala 24:24 25:{25,33}]
  wire  _T_3 = ibf_io_out_valid & idu_io_in_0_ready; // @[src/main/scala/utils/Pipeline.scala 26:22]
  wire  _GEN_1 = ibf_io_out_valid & idu_io_in_0_ready | _GEN_0; // @[src/main/scala/utils/Pipeline.scala 26:{38,46}]
  reg [63:0] idu_io_in_0_bits_r_instr; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg [38:0] idu_io_in_0_bits_r_pc; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg [38:0] idu_io_in_0_bits_r_pnpc; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg  idu_io_in_0_bits_r_exceptionVec_12; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg [3:0] idu_io_in_0_bits_r_brIdx; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg  idu_io_in_0_bits_r_crossPageIPFFix; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg [63:0] c; // @[src/main/scala/utils/GTimer.scala 24:20]
  wire [63:0] _c_T_1 = c + 64'h1; // @[src/main/scala/utils/GTimer.scala 25:12]
  wire  _T_6 = ~reset; // @[src/main/scala/utils/Debug.scala 56:24]
  reg [63:0] c_1; // @[src/main/scala/utils/GTimer.scala 24:20]
  wire [63:0] _c_T_3 = c_1 + 64'h1; // @[src/main/scala/utils/GTimer.scala 25:12]
  reg [63:0] c_2; // @[src/main/scala/utils/GTimer.scala 24:20]
  wire [63:0] _c_T_5 = c_2 + 64'h1; // @[src/main/scala/utils/GTimer.scala 25:12]
  wire  _T_14 = ifu_io_out_valid & DISPLAY_ENABLE; // @[src/main/scala/utils/Debug.scala 55:16]
  reg [63:0] c_3; // @[src/main/scala/utils/GTimer.scala 24:20]
  wire [63:0] _c_T_7 = c_3 + 64'h1; // @[src/main/scala/utils/GTimer.scala 25:12]
  wire  _T_19 = idu_io_in_0_valid & DISPLAY_ENABLE; // @[src/main/scala/utils/Debug.scala 55:16]
  IFU_inorder ifu ( // @[src/main/scala/nutcore/frontend/Frontend.scala 94:20]
    .clock(ifu_clock),
    .reset(ifu_reset),
    .io_imem_req_ready(ifu_io_imem_req_ready),
    .io_imem_req_valid(ifu_io_imem_req_valid),
    .io_imem_req_bits_addr(ifu_io_imem_req_bits_addr),
    .io_imem_req_bits_user(ifu_io_imem_req_bits_user),
    .io_imem_resp_ready(ifu_io_imem_resp_ready),
    .io_imem_resp_valid(ifu_io_imem_resp_valid),
    .io_imem_resp_bits_rdata(ifu_io_imem_resp_bits_rdata),
    .io_imem_resp_bits_user(ifu_io_imem_resp_bits_user),
    .io_out_ready(ifu_io_out_ready),
    .io_out_valid(ifu_io_out_valid),
    .io_out_bits_instr(ifu_io_out_bits_instr),
    .io_out_bits_pc(ifu_io_out_bits_pc),
    .io_out_bits_pnpc(ifu_io_out_bits_pnpc),
    .io_out_bits_exceptionVec_12(ifu_io_out_bits_exceptionVec_12),
    .io_out_bits_brIdx(ifu_io_out_bits_brIdx),
    .io_redirect_target(ifu_io_redirect_target),
    .io_redirect_valid(ifu_io_redirect_valid),
    .io_flushVec(ifu_io_flushVec),
    .io_ipf(ifu_io_ipf),
    .REG_valid(ifu_REG_valid),
    .REG_pc(ifu_REG_pc),
    .REG_isMissPredict(ifu_REG_isMissPredict),
    .REG_actualTarget(ifu_REG_actualTarget),
    .REG_actualTaken(ifu_REG_actualTaken),
    .REG_fuOpType(ifu_REG_fuOpType),
    .REG_btbType(ifu_REG_btbType),
    .REG_isRVC(ifu_REG_isRVC),
    .DISPLAY_ENABLE(ifu_DISPLAY_ENABLE),
    ._WIRE_7(ifu__WIRE_7),
    ._WIRE_11(ifu__WIRE_11),
    ._WIRE_1_4(ifu__WIRE_1_4),
    .r_2(ifu_r_2)
  );
  NaiveRVCAlignBuffer ibf ( // @[src/main/scala/nutcore/frontend/Frontend.scala 95:19]
    .clock(ibf_clock),
    .reset(ibf_reset),
    .io_in_ready(ibf_io_in_ready),
    .io_in_valid(ibf_io_in_valid),
    .io_in_bits_instr(ibf_io_in_bits_instr),
    .io_in_bits_pc(ibf_io_in_bits_pc),
    .io_in_bits_pnpc(ibf_io_in_bits_pnpc),
    .io_in_bits_exceptionVec_12(ibf_io_in_bits_exceptionVec_12),
    .io_in_bits_brIdx(ibf_io_in_bits_brIdx),
    .io_out_ready(ibf_io_out_ready),
    .io_out_valid(ibf_io_out_valid),
    .io_out_bits_instr(ibf_io_out_bits_instr),
    .io_out_bits_pc(ibf_io_out_bits_pc),
    .io_out_bits_pnpc(ibf_io_out_bits_pnpc),
    .io_out_bits_exceptionVec_12(ibf_io_out_bits_exceptionVec_12),
    .io_out_bits_brIdx(ibf_io_out_bits_brIdx),
    .io_out_bits_crossPageIPFFix(ibf_io_out_bits_crossPageIPFFix),
    .io_flush(ibf_io_flush),
    .DISPLAY_ENABLE(ibf_DISPLAY_ENABLE)
  );
  IDU idu ( // @[src/main/scala/nutcore/frontend/Frontend.scala 96:20]
    .clock(idu_clock),
    .reset(idu_reset),
    .io_in_0_ready(idu_io_in_0_ready),
    .io_in_0_valid(idu_io_in_0_valid),
    .io_in_0_bits_instr(idu_io_in_0_bits_instr),
    .io_in_0_bits_pc(idu_io_in_0_bits_pc),
    .io_in_0_bits_pnpc(idu_io_in_0_bits_pnpc),
    .io_in_0_bits_exceptionVec_12(idu_io_in_0_bits_exceptionVec_12),
    .io_in_0_bits_brIdx(idu_io_in_0_bits_brIdx),
    .io_in_0_bits_crossPageIPFFix(idu_io_in_0_bits_crossPageIPFFix),
    .io_out_0_ready(idu_io_out_0_ready),
    .io_out_0_valid(idu_io_out_0_valid),
    .io_out_0_bits_cf_instr(idu_io_out_0_bits_cf_instr),
    .io_out_0_bits_cf_pc(idu_io_out_0_bits_cf_pc),
    .io_out_0_bits_cf_pnpc(idu_io_out_0_bits_cf_pnpc),
    .io_out_0_bits_cf_exceptionVec_1(idu_io_out_0_bits_cf_exceptionVec_1),
    .io_out_0_bits_cf_exceptionVec_2(idu_io_out_0_bits_cf_exceptionVec_2),
    .io_out_0_bits_cf_exceptionVec_12(idu_io_out_0_bits_cf_exceptionVec_12),
    .io_out_0_bits_cf_intrVec_0(idu_io_out_0_bits_cf_intrVec_0),
    .io_out_0_bits_cf_intrVec_1(idu_io_out_0_bits_cf_intrVec_1),
    .io_out_0_bits_cf_intrVec_2(idu_io_out_0_bits_cf_intrVec_2),
    .io_out_0_bits_cf_intrVec_3(idu_io_out_0_bits_cf_intrVec_3),
    .io_out_0_bits_cf_intrVec_4(idu_io_out_0_bits_cf_intrVec_4),
    .io_out_0_bits_cf_intrVec_5(idu_io_out_0_bits_cf_intrVec_5),
    .io_out_0_bits_cf_intrVec_6(idu_io_out_0_bits_cf_intrVec_6),
    .io_out_0_bits_cf_intrVec_7(idu_io_out_0_bits_cf_intrVec_7),
    .io_out_0_bits_cf_intrVec_8(idu_io_out_0_bits_cf_intrVec_8),
    .io_out_0_bits_cf_intrVec_9(idu_io_out_0_bits_cf_intrVec_9),
    .io_out_0_bits_cf_intrVec_10(idu_io_out_0_bits_cf_intrVec_10),
    .io_out_0_bits_cf_intrVec_11(idu_io_out_0_bits_cf_intrVec_11),
    .io_out_0_bits_cf_brIdx(idu_io_out_0_bits_cf_brIdx),
    .io_out_0_bits_cf_crossPageIPFFix(idu_io_out_0_bits_cf_crossPageIPFFix),
    .io_out_0_bits_ctrl_src1Type(idu_io_out_0_bits_ctrl_src1Type),
    .io_out_0_bits_ctrl_src2Type(idu_io_out_0_bits_ctrl_src2Type),
    .io_out_0_bits_ctrl_fuType(idu_io_out_0_bits_ctrl_fuType),
    .io_out_0_bits_ctrl_fuOpType(idu_io_out_0_bits_ctrl_fuOpType),
    .io_out_0_bits_ctrl_rfSrc1(idu_io_out_0_bits_ctrl_rfSrc1),
    .io_out_0_bits_ctrl_rfSrc2(idu_io_out_0_bits_ctrl_rfSrc2),
    .io_out_0_bits_ctrl_rfWen(idu_io_out_0_bits_ctrl_rfWen),
    .io_out_0_bits_ctrl_rfDest(idu_io_out_0_bits_ctrl_rfDest),
    .io_out_0_bits_ctrl_isNutCoreTrap(idu_io_out_0_bits_ctrl_isNutCoreTrap),
    .io_out_0_bits_data_imm(idu_io_out_0_bits_data_imm),
    .io_out_1_bits_cf_intrVec_0(idu_io_out_1_bits_cf_intrVec_0),
    .io_out_1_bits_cf_intrVec_1(idu_io_out_1_bits_cf_intrVec_1),
    .io_out_1_bits_cf_intrVec_2(idu_io_out_1_bits_cf_intrVec_2),
    .io_out_1_bits_cf_intrVec_3(idu_io_out_1_bits_cf_intrVec_3),
    .io_out_1_bits_cf_intrVec_4(idu_io_out_1_bits_cf_intrVec_4),
    .io_out_1_bits_cf_intrVec_5(idu_io_out_1_bits_cf_intrVec_5),
    .io_out_1_bits_cf_intrVec_6(idu_io_out_1_bits_cf_intrVec_6),
    .io_out_1_bits_cf_intrVec_7(idu_io_out_1_bits_cf_intrVec_7),
    .io_out_1_bits_cf_intrVec_8(idu_io_out_1_bits_cf_intrVec_8),
    .io_out_1_bits_cf_intrVec_9(idu_io_out_1_bits_cf_intrVec_9),
    .io_out_1_bits_cf_intrVec_10(idu_io_out_1_bits_cf_intrVec_10),
    .io_out_1_bits_cf_intrVec_11(idu_io_out_1_bits_cf_intrVec_11),
    ._WIRE_1(idu__WIRE_1),
    ._WIRE_5(idu__WIRE_5),
    ._WIRE_14(idu__WIRE_14),
    ._WIRE_2_2(idu__WIRE_2_2)
  );
  FlushableQueue ibf_io_in_q ( // @[src/main/scala/utils/FlushableQueue.scala 94:21]
    .clock(ibf_io_in_q_clock),
    .reset(ibf_io_in_q_reset),
    .io_enq_ready(ibf_io_in_q_io_enq_ready),
    .io_enq_valid(ibf_io_in_q_io_enq_valid),
    .io_enq_bits_instr(ibf_io_in_q_io_enq_bits_instr),
    .io_enq_bits_pc(ibf_io_in_q_io_enq_bits_pc),
    .io_enq_bits_pnpc(ibf_io_in_q_io_enq_bits_pnpc),
    .io_enq_bits_exceptionVec_12(ibf_io_in_q_io_enq_bits_exceptionVec_12),
    .io_enq_bits_brIdx(ibf_io_in_q_io_enq_bits_brIdx),
    .io_deq_ready(ibf_io_in_q_io_deq_ready),
    .io_deq_valid(ibf_io_in_q_io_deq_valid),
    .io_deq_bits_instr(ibf_io_in_q_io_deq_bits_instr),
    .io_deq_bits_pc(ibf_io_in_q_io_deq_bits_pc),
    .io_deq_bits_pnpc(ibf_io_in_q_io_deq_bits_pnpc),
    .io_deq_bits_exceptionVec_12(ibf_io_in_q_io_deq_bits_exceptionVec_12),
    .io_deq_bits_brIdx(ibf_io_in_q_io_deq_bits_brIdx),
    .io_flush(ibf_io_in_q_io_flush)
  );
  assign io_imem_req_valid = ifu_io_imem_req_valid; // @[src/main/scala/nutcore/frontend/Frontend.scala 115:11]
  assign io_imem_req_bits_addr = ifu_io_imem_req_bits_addr; // @[src/main/scala/nutcore/frontend/Frontend.scala 115:11]
  assign io_imem_req_bits_user = {{5'd0}, ifu_io_imem_req_bits_user}; // @[src/main/scala/nutcore/frontend/Frontend.scala 115:11]
  assign io_imem_resp_ready = ifu_io_imem_resp_ready; // @[src/main/scala/nutcore/frontend/Frontend.scala 115:11]
  assign io_out_0_valid = idu_io_out_0_valid; // @[src/main/scala/nutcore/frontend/Frontend.scala 110:10]
  assign io_out_0_bits_cf_instr = idu_io_out_0_bits_cf_instr; // @[src/main/scala/nutcore/frontend/Frontend.scala 110:10]
  assign io_out_0_bits_cf_pc = idu_io_out_0_bits_cf_pc; // @[src/main/scala/nutcore/frontend/Frontend.scala 110:10]
  assign io_out_0_bits_cf_pnpc = idu_io_out_0_bits_cf_pnpc; // @[src/main/scala/nutcore/frontend/Frontend.scala 110:10]
  assign io_out_0_bits_cf_exceptionVec_1 = idu_io_out_0_bits_cf_exceptionVec_1; // @[src/main/scala/nutcore/frontend/Frontend.scala 110:10]
  assign io_out_0_bits_cf_exceptionVec_2 = idu_io_out_0_bits_cf_exceptionVec_2; // @[src/main/scala/nutcore/frontend/Frontend.scala 110:10]
  assign io_out_0_bits_cf_exceptionVec_12 = idu_io_out_0_bits_cf_exceptionVec_12; // @[src/main/scala/nutcore/frontend/Frontend.scala 110:10]
  assign io_out_0_bits_cf_intrVec_0 = idu_io_out_0_bits_cf_intrVec_0; // @[src/main/scala/nutcore/frontend/Frontend.scala 110:10]
  assign io_out_0_bits_cf_intrVec_1 = idu_io_out_0_bits_cf_intrVec_1; // @[src/main/scala/nutcore/frontend/Frontend.scala 110:10]
  assign io_out_0_bits_cf_intrVec_2 = idu_io_out_0_bits_cf_intrVec_2; // @[src/main/scala/nutcore/frontend/Frontend.scala 110:10]
  assign io_out_0_bits_cf_intrVec_3 = idu_io_out_0_bits_cf_intrVec_3; // @[src/main/scala/nutcore/frontend/Frontend.scala 110:10]
  assign io_out_0_bits_cf_intrVec_4 = idu_io_out_0_bits_cf_intrVec_4; // @[src/main/scala/nutcore/frontend/Frontend.scala 110:10]
  assign io_out_0_bits_cf_intrVec_5 = idu_io_out_0_bits_cf_intrVec_5; // @[src/main/scala/nutcore/frontend/Frontend.scala 110:10]
  assign io_out_0_bits_cf_intrVec_6 = idu_io_out_0_bits_cf_intrVec_6; // @[src/main/scala/nutcore/frontend/Frontend.scala 110:10]
  assign io_out_0_bits_cf_intrVec_7 = idu_io_out_0_bits_cf_intrVec_7; // @[src/main/scala/nutcore/frontend/Frontend.scala 110:10]
  assign io_out_0_bits_cf_intrVec_8 = idu_io_out_0_bits_cf_intrVec_8; // @[src/main/scala/nutcore/frontend/Frontend.scala 110:10]
  assign io_out_0_bits_cf_intrVec_9 = idu_io_out_0_bits_cf_intrVec_9; // @[src/main/scala/nutcore/frontend/Frontend.scala 110:10]
  assign io_out_0_bits_cf_intrVec_10 = idu_io_out_0_bits_cf_intrVec_10; // @[src/main/scala/nutcore/frontend/Frontend.scala 110:10]
  assign io_out_0_bits_cf_intrVec_11 = idu_io_out_0_bits_cf_intrVec_11; // @[src/main/scala/nutcore/frontend/Frontend.scala 110:10]
  assign io_out_0_bits_cf_brIdx = idu_io_out_0_bits_cf_brIdx; // @[src/main/scala/nutcore/frontend/Frontend.scala 110:10]
  assign io_out_0_bits_cf_crossPageIPFFix = idu_io_out_0_bits_cf_crossPageIPFFix; // @[src/main/scala/nutcore/frontend/Frontend.scala 110:10]
  assign io_out_0_bits_ctrl_src1Type = idu_io_out_0_bits_ctrl_src1Type; // @[src/main/scala/nutcore/frontend/Frontend.scala 110:10]
  assign io_out_0_bits_ctrl_src2Type = idu_io_out_0_bits_ctrl_src2Type; // @[src/main/scala/nutcore/frontend/Frontend.scala 110:10]
  assign io_out_0_bits_ctrl_fuType = idu_io_out_0_bits_ctrl_fuType; // @[src/main/scala/nutcore/frontend/Frontend.scala 110:10]
  assign io_out_0_bits_ctrl_fuOpType = idu_io_out_0_bits_ctrl_fuOpType; // @[src/main/scala/nutcore/frontend/Frontend.scala 110:10]
  assign io_out_0_bits_ctrl_rfSrc1 = idu_io_out_0_bits_ctrl_rfSrc1; // @[src/main/scala/nutcore/frontend/Frontend.scala 110:10]
  assign io_out_0_bits_ctrl_rfSrc2 = idu_io_out_0_bits_ctrl_rfSrc2; // @[src/main/scala/nutcore/frontend/Frontend.scala 110:10]
  assign io_out_0_bits_ctrl_rfWen = idu_io_out_0_bits_ctrl_rfWen; // @[src/main/scala/nutcore/frontend/Frontend.scala 110:10]
  assign io_out_0_bits_ctrl_rfDest = idu_io_out_0_bits_ctrl_rfDest; // @[src/main/scala/nutcore/frontend/Frontend.scala 110:10]
  assign io_out_0_bits_ctrl_isNutCoreTrap = idu_io_out_0_bits_ctrl_isNutCoreTrap; // @[src/main/scala/nutcore/frontend/Frontend.scala 110:10]
  assign io_out_0_bits_data_imm = idu_io_out_0_bits_data_imm; // @[src/main/scala/nutcore/frontend/Frontend.scala 110:10]
  assign io_out_1_bits_cf_intrVec_0 = idu_io_out_1_bits_cf_intrVec_0; // @[src/main/scala/nutcore/frontend/Frontend.scala 110:10]
  assign io_out_1_bits_cf_intrVec_1 = idu_io_out_1_bits_cf_intrVec_1; // @[src/main/scala/nutcore/frontend/Frontend.scala 110:10]
  assign io_out_1_bits_cf_intrVec_2 = idu_io_out_1_bits_cf_intrVec_2; // @[src/main/scala/nutcore/frontend/Frontend.scala 110:10]
  assign io_out_1_bits_cf_intrVec_3 = idu_io_out_1_bits_cf_intrVec_3; // @[src/main/scala/nutcore/frontend/Frontend.scala 110:10]
  assign io_out_1_bits_cf_intrVec_4 = idu_io_out_1_bits_cf_intrVec_4; // @[src/main/scala/nutcore/frontend/Frontend.scala 110:10]
  assign io_out_1_bits_cf_intrVec_5 = idu_io_out_1_bits_cf_intrVec_5; // @[src/main/scala/nutcore/frontend/Frontend.scala 110:10]
  assign io_out_1_bits_cf_intrVec_6 = idu_io_out_1_bits_cf_intrVec_6; // @[src/main/scala/nutcore/frontend/Frontend.scala 110:10]
  assign io_out_1_bits_cf_intrVec_7 = idu_io_out_1_bits_cf_intrVec_7; // @[src/main/scala/nutcore/frontend/Frontend.scala 110:10]
  assign io_out_1_bits_cf_intrVec_8 = idu_io_out_1_bits_cf_intrVec_8; // @[src/main/scala/nutcore/frontend/Frontend.scala 110:10]
  assign io_out_1_bits_cf_intrVec_9 = idu_io_out_1_bits_cf_intrVec_9; // @[src/main/scala/nutcore/frontend/Frontend.scala 110:10]
  assign io_out_1_bits_cf_intrVec_10 = idu_io_out_1_bits_cf_intrVec_10; // @[src/main/scala/nutcore/frontend/Frontend.scala 110:10]
  assign io_out_1_bits_cf_intrVec_11 = idu_io_out_1_bits_cf_intrVec_11; // @[src/main/scala/nutcore/frontend/Frontend.scala 110:10]
  assign io_flushVec = ifu_io_flushVec; // @[src/main/scala/nutcore/frontend/Frontend.scala 112:15]
  assign _WIRE_0 = idu__WIRE_1;
  assign _WIRE_7 = ifu__WIRE_7;
  assign r_0 = ifu_r_2;
  assign ifu_clock = clock;
  assign ifu_reset = reset;
  assign ifu_io_imem_req_ready = io_imem_req_ready; // @[src/main/scala/nutcore/frontend/Frontend.scala 115:11]
  assign ifu_io_imem_resp_valid = io_imem_resp_valid; // @[src/main/scala/nutcore/frontend/Frontend.scala 115:11]
  assign ifu_io_imem_resp_bits_rdata = io_imem_resp_bits_rdata; // @[src/main/scala/nutcore/frontend/Frontend.scala 115:11]
  assign ifu_io_imem_resp_bits_user = io_imem_resp_bits_user[81:0]; // @[src/main/scala/nutcore/frontend/Frontend.scala 115:11]
  assign ifu_io_out_ready = ibf_io_in_q_io_enq_ready; // @[src/main/scala/utils/FlushableQueue.scala 98:17]
  assign ifu_io_redirect_target = io_redirect_target; // @[src/main/scala/nutcore/frontend/Frontend.scala 111:15]
  assign ifu_io_redirect_valid = io_redirect_valid; // @[src/main/scala/nutcore/frontend/Frontend.scala 111:15]
  assign ifu_io_ipf = io_ipf; // @[src/main/scala/nutcore/frontend/Frontend.scala 114:10]
  assign ifu_REG_valid = REG_valid;
  assign ifu_REG_pc = REG_pc;
  assign ifu_REG_isMissPredict = REG_isMissPredict;
  assign ifu_REG_actualTarget = REG_actualTarget;
  assign ifu_REG_actualTaken = REG_actualTaken;
  assign ifu_REG_fuOpType = REG_fuOpType;
  assign ifu_REG_btbType = REG_btbType;
  assign ifu_REG_isRVC = REG_isRVC;
  assign ifu_DISPLAY_ENABLE = DISPLAY_ENABLE;
  assign ifu__WIRE_11 = _WIRE_11;
  assign ifu__WIRE_1_4 = _WIRE_1_4;
  assign ibf_clock = clock;
  assign ibf_reset = reset;
  assign ibf_io_in_valid = ibf_io_in_q_io_deq_valid; // @[src/main/scala/nutcore/frontend/Frontend.scala 102:11]
  assign ibf_io_in_bits_instr = ibf_io_in_q_io_deq_bits_instr; // @[src/main/scala/nutcore/frontend/Frontend.scala 102:11]
  assign ibf_io_in_bits_pc = ibf_io_in_q_io_deq_bits_pc; // @[src/main/scala/nutcore/frontend/Frontend.scala 102:11]
  assign ibf_io_in_bits_pnpc = ibf_io_in_q_io_deq_bits_pnpc; // @[src/main/scala/nutcore/frontend/Frontend.scala 102:11]
  assign ibf_io_in_bits_exceptionVec_12 = ibf_io_in_q_io_deq_bits_exceptionVec_12; // @[src/main/scala/nutcore/frontend/Frontend.scala 102:11]
  assign ibf_io_in_bits_brIdx = ibf_io_in_q_io_deq_bits_brIdx; // @[src/main/scala/nutcore/frontend/Frontend.scala 102:11]
  assign ibf_io_out_ready = idu_io_in_0_ready; // @[src/main/scala/utils/Pipeline.scala 29:16]
  assign ibf_io_flush = ifu_io_flushVec[1]; // @[src/main/scala/nutcore/frontend/Frontend.scala 109:34]
  assign ibf_DISPLAY_ENABLE = DISPLAY_ENABLE;
  assign idu_clock = clock;
  assign idu_reset = reset;
  assign idu_io_in_0_valid = valid; // @[src/main/scala/utils/Pipeline.scala 31:17]
  assign idu_io_in_0_bits_instr = idu_io_in_0_bits_r_instr; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign idu_io_in_0_bits_pc = idu_io_in_0_bits_r_pc; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign idu_io_in_0_bits_pnpc = idu_io_in_0_bits_r_pnpc; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign idu_io_in_0_bits_exceptionVec_12 = idu_io_in_0_bits_r_exceptionVec_12; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign idu_io_in_0_bits_brIdx = idu_io_in_0_bits_r_brIdx; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign idu_io_in_0_bits_crossPageIPFFix = idu_io_in_0_bits_r_crossPageIPFFix; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign idu_io_out_0_ready = io_out_0_ready; // @[src/main/scala/nutcore/frontend/Frontend.scala 110:10]
  assign idu__WIRE_5 = DISPLAY_ENABLE;
  assign idu__WIRE_14 = _WIRE_14;
  assign idu__WIRE_2_2 = _WIRE_2_2;
  assign ibf_io_in_q_clock = clock;
  assign ibf_io_in_q_reset = reset;
  assign ibf_io_in_q_io_enq_valid = ifu_io_out_valid; // @[src/main/scala/utils/FlushableQueue.scala 95:22]
  assign ibf_io_in_q_io_enq_bits_instr = ifu_io_out_bits_instr; // @[src/main/scala/utils/FlushableQueue.scala 96:21]
  assign ibf_io_in_q_io_enq_bits_pc = ifu_io_out_bits_pc; // @[src/main/scala/utils/FlushableQueue.scala 96:21]
  assign ibf_io_in_q_io_enq_bits_pnpc = ifu_io_out_bits_pnpc; // @[src/main/scala/utils/FlushableQueue.scala 96:21]
  assign ibf_io_in_q_io_enq_bits_exceptionVec_12 = ifu_io_out_bits_exceptionVec_12; // @[src/main/scala/utils/FlushableQueue.scala 96:21]
  assign ibf_io_in_q_io_enq_bits_brIdx = ifu_io_out_bits_brIdx; // @[src/main/scala/utils/FlushableQueue.scala 96:21]
  assign ibf_io_in_q_io_deq_ready = ibf_io_in_ready; // @[src/main/scala/nutcore/frontend/Frontend.scala 102:11]
  assign ibf_io_in_q_io_flush = ifu_io_flushVec[0]; // @[src/main/scala/nutcore/frontend/Frontend.scala 105:58]
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/utils/Pipeline.scala 24:24]
      valid <= 1'h0; // @[src/main/scala/utils/Pipeline.scala 24:24]
    end else if (ifu_io_flushVec[1]) begin // @[src/main/scala/utils/Pipeline.scala 27:20]
      valid <= 1'h0; // @[src/main/scala/utils/Pipeline.scala 27:28]
    end else begin
      valid <= _GEN_1;
    end
    if (_T_3) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      idu_io_in_0_bits_r_instr <= ibf_io_out_bits_instr; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_3) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      idu_io_in_0_bits_r_pc <= ibf_io_out_bits_pc; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_3) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      idu_io_in_0_bits_r_pnpc <= ibf_io_out_bits_pnpc; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_3) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      idu_io_in_0_bits_r_exceptionVec_12 <= ibf_io_out_bits_exceptionVec_12; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_3) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      idu_io_in_0_bits_r_brIdx <= ibf_io_out_bits_brIdx; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_3) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      idu_io_in_0_bits_r_crossPageIPFFix <= ibf_io_out_bits_crossPageIPFFix; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (reset) begin // @[src/main/scala/utils/GTimer.scala 24:20]
      c <= 64'h0; // @[src/main/scala/utils/GTimer.scala 24:20]
    end else begin
      c <= _c_T_1; // @[src/main/scala/utils/GTimer.scala 25:7]
    end
    if (reset) begin // @[src/main/scala/utils/GTimer.scala 24:20]
      c_1 <= 64'h0; // @[src/main/scala/utils/GTimer.scala 24:20]
    end else begin
      c_1 <= _c_T_3; // @[src/main/scala/utils/GTimer.scala 25:7]
    end
    if (reset) begin // @[src/main/scala/utils/GTimer.scala 24:20]
      c_2 <= 64'h0; // @[src/main/scala/utils/GTimer.scala 24:20]
    end else begin
      c_2 <= _c_T_5; // @[src/main/scala/utils/GTimer.scala 25:7]
    end
    if (reset) begin // @[src/main/scala/utils/GTimer.scala 24:20]
      c_3 <= 64'h0; // @[src/main/scala/utils/GTimer.scala 24:20]
    end else begin
      c_3 <= _c_T_7; // @[src/main/scala/utils/GTimer.scala 25:7]
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & ~reset) begin
          $fwrite(32'h80000002,"[%d] Frontend_inorder: ",c); // @[src/main/scala/utils/Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_6) begin
          $fwrite(32'h80000002,"------------------------ FRONTEND:------------------------\n"); // @[src/main/scala/utils/Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & ~reset) begin
          $fwrite(32'h80000002,"[%d] Frontend_inorder: ",c_1); // @[src/main/scala/utils/Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_6) begin
          $fwrite(32'h80000002,"flush = %b, ifu:(%d,%d), idu:(%d,%d)\n",ifu_io_flushVec,ifu_io_out_valid,
            ifu_io_out_ready,idu_io_in_0_valid,idu_io_in_0_ready); // @[src/main/scala/utils/Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_14 & ~reset) begin
          $fwrite(32'h80000002,"[%d] Frontend_inorder: ",c_2); // @[src/main/scala/utils/Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_14 & _T_6) begin
          $fwrite(32'h80000002,"IFU: pc = 0x%x, instr = 0x%x\n",ifu_io_out_bits_pc,ifu_io_out_bits_instr); // @[src/main/scala/utils/Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_19 & ~reset) begin
          $fwrite(32'h80000002,"[%d] Frontend_inorder: ",c_3); // @[src/main/scala/utils/Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_19 & _T_6) begin
          $fwrite(32'h80000002,"IDU1: pc = 0x%x, instr = 0x%x, pnpc = 0x%x\n",idu_io_in_0_bits_pc,idu_io_in_0_bits_instr
            ,idu_io_in_0_bits_pnpc); // @[src/main/scala/utils/Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  valid = _RAND_0[0:0];
  _RAND_1 = {2{`RANDOM}};
  idu_io_in_0_bits_r_instr = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  idu_io_in_0_bits_r_pc = _RAND_2[38:0];
  _RAND_3 = {2{`RANDOM}};
  idu_io_in_0_bits_r_pnpc = _RAND_3[38:0];
  _RAND_4 = {1{`RANDOM}};
  idu_io_in_0_bits_r_exceptionVec_12 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  idu_io_in_0_bits_r_brIdx = _RAND_5[3:0];
  _RAND_6 = {1{`RANDOM}};
  idu_io_in_0_bits_r_crossPageIPFFix = _RAND_6[0:0];
  _RAND_7 = {2{`RANDOM}};
  c = _RAND_7[63:0];
  _RAND_8 = {2{`RANDOM}};
  c_1 = _RAND_8[63:0];
  _RAND_9 = {2{`RANDOM}};
  c_2 = _RAND_9[63:0];
  _RAND_10 = {2{`RANDOM}};
  c_3 = _RAND_10[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ISU(
  input         clock,
  input         reset,
  output        io_in_0_ready, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  input         io_in_0_valid, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  input  [63:0] io_in_0_bits_cf_instr, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  input  [38:0] io_in_0_bits_cf_pc, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  input  [38:0] io_in_0_bits_cf_pnpc, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  input         io_in_0_bits_cf_exceptionVec_1, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  input         io_in_0_bits_cf_exceptionVec_2, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  input         io_in_0_bits_cf_exceptionVec_12, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  input         io_in_0_bits_cf_intrVec_0, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  input         io_in_0_bits_cf_intrVec_1, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  input         io_in_0_bits_cf_intrVec_2, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  input         io_in_0_bits_cf_intrVec_3, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  input         io_in_0_bits_cf_intrVec_4, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  input         io_in_0_bits_cf_intrVec_5, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  input         io_in_0_bits_cf_intrVec_6, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  input         io_in_0_bits_cf_intrVec_7, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  input         io_in_0_bits_cf_intrVec_8, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  input         io_in_0_bits_cf_intrVec_9, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  input         io_in_0_bits_cf_intrVec_10, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  input         io_in_0_bits_cf_intrVec_11, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  input  [3:0]  io_in_0_bits_cf_brIdx, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  input         io_in_0_bits_cf_crossPageIPFFix, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  input         io_in_0_bits_ctrl_src1Type, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  input         io_in_0_bits_ctrl_src2Type, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  input  [2:0]  io_in_0_bits_ctrl_fuType, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  input  [6:0]  io_in_0_bits_ctrl_fuOpType, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  input  [4:0]  io_in_0_bits_ctrl_rfSrc1, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  input  [4:0]  io_in_0_bits_ctrl_rfSrc2, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  input         io_in_0_bits_ctrl_rfWen, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  input  [4:0]  io_in_0_bits_ctrl_rfDest, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  input         io_in_0_bits_ctrl_isNutCoreTrap, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  input  [63:0] io_in_0_bits_data_imm, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  input         io_out_ready, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  output        io_out_valid, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  output [63:0] io_out_bits_cf_instr, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  output [38:0] io_out_bits_cf_pc, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  output [38:0] io_out_bits_cf_pnpc, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  output        io_out_bits_cf_exceptionVec_1, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  output        io_out_bits_cf_exceptionVec_2, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  output        io_out_bits_cf_exceptionVec_12, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  output        io_out_bits_cf_intrVec_0, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  output        io_out_bits_cf_intrVec_1, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  output        io_out_bits_cf_intrVec_2, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  output        io_out_bits_cf_intrVec_3, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  output        io_out_bits_cf_intrVec_4, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  output        io_out_bits_cf_intrVec_5, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  output        io_out_bits_cf_intrVec_6, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  output        io_out_bits_cf_intrVec_7, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  output        io_out_bits_cf_intrVec_8, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  output        io_out_bits_cf_intrVec_9, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  output        io_out_bits_cf_intrVec_10, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  output        io_out_bits_cf_intrVec_11, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  output [3:0]  io_out_bits_cf_brIdx, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  output        io_out_bits_cf_crossPageIPFFix, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  output [2:0]  io_out_bits_ctrl_fuType, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  output [6:0]  io_out_bits_ctrl_fuOpType, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  output        io_out_bits_ctrl_rfWen, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  output [4:0]  io_out_bits_ctrl_rfDest, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  output        io_out_bits_ctrl_isNutCoreTrap, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  output [63:0] io_out_bits_data_src1, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  output [63:0] io_out_bits_data_src2, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  output [63:0] io_out_bits_data_imm, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  input         io_wb_rfWen, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  input  [4:0]  io_wb_rfDest, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  input  [63:0] io_wb_rfData, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  input         io_forward_valid, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  input         io_forward_wb_rfWen, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  input  [4:0]  io_forward_wb_rfDest, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  input  [63:0] io_forward_wb_rfData, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  input  [2:0]  io_forward_fuType, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  input         io_flush, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  output        _WIRE_1_0,
  input         DISPLAY_ENABLE,
  output        _WIRE_8,
  output        _WIRE_2_2
);
`ifdef RANDOMIZE_MEM_INIT
  reg [63:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [63:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg [63:0] rf [0:31]; // @[src/main/scala/nutcore/RF.scala 30:15]
  wire  rf_io_out_bits_data_src1_MPORT_en; // @[src/main/scala/nutcore/RF.scala 30:15]
  wire [4:0] rf_io_out_bits_data_src1_MPORT_addr; // @[src/main/scala/nutcore/RF.scala 30:15]
  wire [63:0] rf_io_out_bits_data_src1_MPORT_data; // @[src/main/scala/nutcore/RF.scala 30:15]
  wire  rf_io_out_bits_data_src2_MPORT_en; // @[src/main/scala/nutcore/RF.scala 30:15]
  wire [4:0] rf_io_out_bits_data_src2_MPORT_addr; // @[src/main/scala/nutcore/RF.scala 30:15]
  wire [63:0] rf_io_out_bits_data_src2_MPORT_data; // @[src/main/scala/nutcore/RF.scala 30:15]
  wire  rf_MPORT_1_en; // @[src/main/scala/nutcore/RF.scala 30:15]
  wire [4:0] rf_MPORT_1_addr; // @[src/main/scala/nutcore/RF.scala 30:15]
  wire [63:0] rf_MPORT_1_data; // @[src/main/scala/nutcore/RF.scala 30:15]
  wire  rf_MPORT_2_en; // @[src/main/scala/nutcore/RF.scala 30:15]
  wire [4:0] rf_MPORT_2_addr; // @[src/main/scala/nutcore/RF.scala 30:15]
  wire [63:0] rf_MPORT_2_data; // @[src/main/scala/nutcore/RF.scala 30:15]
  wire  rf_MPORT_3_en; // @[src/main/scala/nutcore/RF.scala 30:15]
  wire [4:0] rf_MPORT_3_addr; // @[src/main/scala/nutcore/RF.scala 30:15]
  wire [63:0] rf_MPORT_3_data; // @[src/main/scala/nutcore/RF.scala 30:15]
  wire  rf_MPORT_4_en; // @[src/main/scala/nutcore/RF.scala 30:15]
  wire [4:0] rf_MPORT_4_addr; // @[src/main/scala/nutcore/RF.scala 30:15]
  wire [63:0] rf_MPORT_4_data; // @[src/main/scala/nutcore/RF.scala 30:15]
  wire  rf_MPORT_5_en; // @[src/main/scala/nutcore/RF.scala 30:15]
  wire [4:0] rf_MPORT_5_addr; // @[src/main/scala/nutcore/RF.scala 30:15]
  wire [63:0] rf_MPORT_5_data; // @[src/main/scala/nutcore/RF.scala 30:15]
  wire  rf_MPORT_6_en; // @[src/main/scala/nutcore/RF.scala 30:15]
  wire [4:0] rf_MPORT_6_addr; // @[src/main/scala/nutcore/RF.scala 30:15]
  wire [63:0] rf_MPORT_6_data; // @[src/main/scala/nutcore/RF.scala 30:15]
  wire  rf_MPORT_7_en; // @[src/main/scala/nutcore/RF.scala 30:15]
  wire [4:0] rf_MPORT_7_addr; // @[src/main/scala/nutcore/RF.scala 30:15]
  wire [63:0] rf_MPORT_7_data; // @[src/main/scala/nutcore/RF.scala 30:15]
  wire  rf_MPORT_8_en; // @[src/main/scala/nutcore/RF.scala 30:15]
  wire [4:0] rf_MPORT_8_addr; // @[src/main/scala/nutcore/RF.scala 30:15]
  wire [63:0] rf_MPORT_8_data; // @[src/main/scala/nutcore/RF.scala 30:15]
  wire  rf_MPORT_9_en; // @[src/main/scala/nutcore/RF.scala 30:15]
  wire [4:0] rf_MPORT_9_addr; // @[src/main/scala/nutcore/RF.scala 30:15]
  wire [63:0] rf_MPORT_9_data; // @[src/main/scala/nutcore/RF.scala 30:15]
  wire  rf_MPORT_10_en; // @[src/main/scala/nutcore/RF.scala 30:15]
  wire [4:0] rf_MPORT_10_addr; // @[src/main/scala/nutcore/RF.scala 30:15]
  wire [63:0] rf_MPORT_10_data; // @[src/main/scala/nutcore/RF.scala 30:15]
  wire  rf_MPORT_11_en; // @[src/main/scala/nutcore/RF.scala 30:15]
  wire [4:0] rf_MPORT_11_addr; // @[src/main/scala/nutcore/RF.scala 30:15]
  wire [63:0] rf_MPORT_11_data; // @[src/main/scala/nutcore/RF.scala 30:15]
  wire  rf_MPORT_12_en; // @[src/main/scala/nutcore/RF.scala 30:15]
  wire [4:0] rf_MPORT_12_addr; // @[src/main/scala/nutcore/RF.scala 30:15]
  wire [63:0] rf_MPORT_12_data; // @[src/main/scala/nutcore/RF.scala 30:15]
  wire  rf_MPORT_13_en; // @[src/main/scala/nutcore/RF.scala 30:15]
  wire [4:0] rf_MPORT_13_addr; // @[src/main/scala/nutcore/RF.scala 30:15]
  wire [63:0] rf_MPORT_13_data; // @[src/main/scala/nutcore/RF.scala 30:15]
  wire  rf_MPORT_14_en; // @[src/main/scala/nutcore/RF.scala 30:15]
  wire [4:0] rf_MPORT_14_addr; // @[src/main/scala/nutcore/RF.scala 30:15]
  wire [63:0] rf_MPORT_14_data; // @[src/main/scala/nutcore/RF.scala 30:15]
  wire  rf_MPORT_15_en; // @[src/main/scala/nutcore/RF.scala 30:15]
  wire [4:0] rf_MPORT_15_addr; // @[src/main/scala/nutcore/RF.scala 30:15]
  wire [63:0] rf_MPORT_15_data; // @[src/main/scala/nutcore/RF.scala 30:15]
  wire  rf_MPORT_16_en; // @[src/main/scala/nutcore/RF.scala 30:15]
  wire [4:0] rf_MPORT_16_addr; // @[src/main/scala/nutcore/RF.scala 30:15]
  wire [63:0] rf_MPORT_16_data; // @[src/main/scala/nutcore/RF.scala 30:15]
  wire  rf_MPORT_17_en; // @[src/main/scala/nutcore/RF.scala 30:15]
  wire [4:0] rf_MPORT_17_addr; // @[src/main/scala/nutcore/RF.scala 30:15]
  wire [63:0] rf_MPORT_17_data; // @[src/main/scala/nutcore/RF.scala 30:15]
  wire  rf_MPORT_18_en; // @[src/main/scala/nutcore/RF.scala 30:15]
  wire [4:0] rf_MPORT_18_addr; // @[src/main/scala/nutcore/RF.scala 30:15]
  wire [63:0] rf_MPORT_18_data; // @[src/main/scala/nutcore/RF.scala 30:15]
  wire  rf_MPORT_19_en; // @[src/main/scala/nutcore/RF.scala 30:15]
  wire [4:0] rf_MPORT_19_addr; // @[src/main/scala/nutcore/RF.scala 30:15]
  wire [63:0] rf_MPORT_19_data; // @[src/main/scala/nutcore/RF.scala 30:15]
  wire  rf_MPORT_20_en; // @[src/main/scala/nutcore/RF.scala 30:15]
  wire [4:0] rf_MPORT_20_addr; // @[src/main/scala/nutcore/RF.scala 30:15]
  wire [63:0] rf_MPORT_20_data; // @[src/main/scala/nutcore/RF.scala 30:15]
  wire  rf_MPORT_21_en; // @[src/main/scala/nutcore/RF.scala 30:15]
  wire [4:0] rf_MPORT_21_addr; // @[src/main/scala/nutcore/RF.scala 30:15]
  wire [63:0] rf_MPORT_21_data; // @[src/main/scala/nutcore/RF.scala 30:15]
  wire  rf_MPORT_22_en; // @[src/main/scala/nutcore/RF.scala 30:15]
  wire [4:0] rf_MPORT_22_addr; // @[src/main/scala/nutcore/RF.scala 30:15]
  wire [63:0] rf_MPORT_22_data; // @[src/main/scala/nutcore/RF.scala 30:15]
  wire  rf_MPORT_23_en; // @[src/main/scala/nutcore/RF.scala 30:15]
  wire [4:0] rf_MPORT_23_addr; // @[src/main/scala/nutcore/RF.scala 30:15]
  wire [63:0] rf_MPORT_23_data; // @[src/main/scala/nutcore/RF.scala 30:15]
  wire  rf_MPORT_24_en; // @[src/main/scala/nutcore/RF.scala 30:15]
  wire [4:0] rf_MPORT_24_addr; // @[src/main/scala/nutcore/RF.scala 30:15]
  wire [63:0] rf_MPORT_24_data; // @[src/main/scala/nutcore/RF.scala 30:15]
  wire  rf_MPORT_25_en; // @[src/main/scala/nutcore/RF.scala 30:15]
  wire [4:0] rf_MPORT_25_addr; // @[src/main/scala/nutcore/RF.scala 30:15]
  wire [63:0] rf_MPORT_25_data; // @[src/main/scala/nutcore/RF.scala 30:15]
  wire  rf_MPORT_26_en; // @[src/main/scala/nutcore/RF.scala 30:15]
  wire [4:0] rf_MPORT_26_addr; // @[src/main/scala/nutcore/RF.scala 30:15]
  wire [63:0] rf_MPORT_26_data; // @[src/main/scala/nutcore/RF.scala 30:15]
  wire  rf_MPORT_27_en; // @[src/main/scala/nutcore/RF.scala 30:15]
  wire [4:0] rf_MPORT_27_addr; // @[src/main/scala/nutcore/RF.scala 30:15]
  wire [63:0] rf_MPORT_27_data; // @[src/main/scala/nutcore/RF.scala 30:15]
  wire  rf_MPORT_28_en; // @[src/main/scala/nutcore/RF.scala 30:15]
  wire [4:0] rf_MPORT_28_addr; // @[src/main/scala/nutcore/RF.scala 30:15]
  wire [63:0] rf_MPORT_28_data; // @[src/main/scala/nutcore/RF.scala 30:15]
  wire  rf_MPORT_29_en; // @[src/main/scala/nutcore/RF.scala 30:15]
  wire [4:0] rf_MPORT_29_addr; // @[src/main/scala/nutcore/RF.scala 30:15]
  wire [63:0] rf_MPORT_29_data; // @[src/main/scala/nutcore/RF.scala 30:15]
  wire  rf_MPORT_30_en; // @[src/main/scala/nutcore/RF.scala 30:15]
  wire [4:0] rf_MPORT_30_addr; // @[src/main/scala/nutcore/RF.scala 30:15]
  wire [63:0] rf_MPORT_30_data; // @[src/main/scala/nutcore/RF.scala 30:15]
  wire  rf_MPORT_31_en; // @[src/main/scala/nutcore/RF.scala 30:15]
  wire [4:0] rf_MPORT_31_addr; // @[src/main/scala/nutcore/RF.scala 30:15]
  wire [63:0] rf_MPORT_31_data; // @[src/main/scala/nutcore/RF.scala 30:15]
  wire  rf_MPORT_32_en; // @[src/main/scala/nutcore/RF.scala 30:15]
  wire [4:0] rf_MPORT_32_addr; // @[src/main/scala/nutcore/RF.scala 30:15]
  wire [63:0] rf_MPORT_32_data; // @[src/main/scala/nutcore/RF.scala 30:15]
  wire [63:0] rf_MPORT_data; // @[src/main/scala/nutcore/RF.scala 30:15]
  wire [4:0] rf_MPORT_addr; // @[src/main/scala/nutcore/RF.scala 30:15]
  wire  rf_MPORT_mask; // @[src/main/scala/nutcore/RF.scala 30:15]
  wire  rf_MPORT_en; // @[src/main/scala/nutcore/RF.scala 30:15]
  wire  forwardRfWen = io_forward_wb_rfWen & io_forward_valid; // @[src/main/scala/nutcore/backend/seq/ISU.scala 43:42]
  wire  dontForward1 = io_forward_fuType != 3'h0 & io_forward_fuType != 3'h1; // @[src/main/scala/nutcore/backend/seq/ISU.scala 44:57]
  wire  src1DependEX = io_in_0_bits_ctrl_rfSrc1 != 5'h0 & io_in_0_bits_ctrl_rfSrc1 == io_forward_wb_rfDest &
    forwardRfWen; // @[src/main/scala/nutcore/backend/seq/ISU.scala 41:100]
  wire  src2DependEX = io_in_0_bits_ctrl_rfSrc2 != 5'h0 & io_in_0_bits_ctrl_rfSrc2 == io_forward_wb_rfDest &
    forwardRfWen; // @[src/main/scala/nutcore/backend/seq/ISU.scala 41:100]
  wire  src1DependWB = io_in_0_bits_ctrl_rfSrc1 != 5'h0 & io_in_0_bits_ctrl_rfSrc1 == io_wb_rfDest & io_wb_rfWen; // @[src/main/scala/nutcore/backend/seq/ISU.scala 41:100]
  wire  src2DependWB = io_in_0_bits_ctrl_rfSrc2 != 5'h0 & io_in_0_bits_ctrl_rfSrc2 == io_wb_rfDest & io_wb_rfWen; // @[src/main/scala/nutcore/backend/seq/ISU.scala 41:100]
  wire  _src1ForwardNextCycle_T = ~dontForward1; // @[src/main/scala/nutcore/backend/seq/ISU.scala 50:46]
  wire  src1ForwardNextCycle = src1DependEX & ~dontForward1; // @[src/main/scala/nutcore/backend/seq/ISU.scala 50:43]
  wire  src2ForwardNextCycle = src2DependEX & _src1ForwardNextCycle_T; // @[src/main/scala/nutcore/backend/seq/ISU.scala 51:43]
  wire  _src1Forward_T_1 = dontForward1 ? ~src1DependEX : 1'h1; // @[src/main/scala/nutcore/backend/seq/ISU.scala 52:40]
  wire  src1Forward = src1DependWB & _src1Forward_T_1; // @[src/main/scala/nutcore/backend/seq/ISU.scala 52:34]
  wire  _src2Forward_T_1 = dontForward1 ? ~src2DependEX : 1'h1; // @[src/main/scala/nutcore/backend/seq/ISU.scala 53:40]
  wire  src2Forward = src2DependWB & _src2Forward_T_1; // @[src/main/scala/nutcore/backend/seq/ISU.scala 53:34]
  reg [31:0] busy; // @[src/main/scala/nutcore/RF.scala 36:21]
  wire [31:0] _src1Ready_T = busy >> io_in_0_bits_ctrl_rfSrc1; // @[src/main/scala/nutcore/RF.scala 37:37]
  wire  src1Ready = ~_src1Ready_T[0] | src1ForwardNextCycle | src1Forward; // @[src/main/scala/nutcore/backend/seq/ISU.scala 56:62]
  wire [31:0] _src2Ready_T = busy >> io_in_0_bits_ctrl_rfSrc2; // @[src/main/scala/nutcore/RF.scala 37:37]
  wire  src2Ready = ~_src2Ready_T[0] | src2ForwardNextCycle | src2Forward; // @[src/main/scala/nutcore/backend/seq/ISU.scala 57:62]
  wire  io_out_bits_data_src1_signBit = io_in_0_bits_cf_pc[38]; // @[src/main/scala/utils/BitUtils.scala 41:20]
  wire [24:0] _io_out_bits_data_src1_T_2 = io_out_bits_data_src1_signBit ? 25'h1ffffff : 25'h0; // @[src/main/scala/utils/BitUtils.scala 42:46]
  wire [63:0] _io_out_bits_data_src1_T_3 = {_io_out_bits_data_src1_T_2,io_in_0_bits_cf_pc}; // @[src/main/scala/utils/BitUtils.scala 42:41]
  wire  _io_out_bits_data_src1_T_4 = ~src1ForwardNextCycle; // @[src/main/scala/nutcore/backend/seq/ISU.scala 66:21]
  wire  _io_out_bits_data_src1_T_5 = src1Forward & ~src1ForwardNextCycle; // @[src/main/scala/nutcore/backend/seq/ISU.scala 66:18]
  wire  _io_out_bits_data_src1_T_10 = ~io_in_0_bits_ctrl_src1Type & _io_out_bits_data_src1_T_4 & ~src1Forward; // @[src/main/scala/nutcore/backend/seq/ISU.scala 67:76]
  wire [63:0] _io_out_bits_data_src1_T_12 = io_in_0_bits_ctrl_rfSrc1 == 5'h0 ? 64'h0 :
    rf_io_out_bits_data_src1_MPORT_data; // @[src/main/scala/nutcore/RF.scala 31:36]
  wire [63:0] _io_out_bits_data_src1_T_13 = io_in_0_bits_ctrl_src1Type ? _io_out_bits_data_src1_T_3 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_out_bits_data_src1_T_14 = src1ForwardNextCycle ? io_forward_wb_rfData : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_out_bits_data_src1_T_15 = _io_out_bits_data_src1_T_5 ? io_wb_rfData : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_out_bits_data_src1_T_16 = _io_out_bits_data_src1_T_10 ? _io_out_bits_data_src1_T_12 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_out_bits_data_src1_T_17 = _io_out_bits_data_src1_T_13 | _io_out_bits_data_src1_T_14; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_out_bits_data_src1_T_18 = _io_out_bits_data_src1_T_17 | _io_out_bits_data_src1_T_15; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _io_out_bits_data_src2_T_1 = ~src2ForwardNextCycle; // @[src/main/scala/nutcore/backend/seq/ISU.scala 72:21]
  wire  _io_out_bits_data_src2_T_2 = src2Forward & ~src2ForwardNextCycle; // @[src/main/scala/nutcore/backend/seq/ISU.scala 72:18]
  wire  _io_out_bits_data_src2_T_7 = ~io_in_0_bits_ctrl_src2Type & _io_out_bits_data_src2_T_1 & ~src2Forward; // @[src/main/scala/nutcore/backend/seq/ISU.scala 73:77]
  wire [63:0] _io_out_bits_data_src2_T_9 = io_in_0_bits_ctrl_rfSrc2 == 5'h0 ? 64'h0 :
    rf_io_out_bits_data_src2_MPORT_data; // @[src/main/scala/nutcore/RF.scala 31:36]
  wire [63:0] _io_out_bits_data_src2_T_10 = io_in_0_bits_ctrl_src2Type ? io_in_0_bits_data_imm : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_out_bits_data_src2_T_11 = src2ForwardNextCycle ? io_forward_wb_rfData : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_out_bits_data_src2_T_12 = _io_out_bits_data_src2_T_2 ? io_wb_rfData : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_out_bits_data_src2_T_13 = _io_out_bits_data_src2_T_7 ? _io_out_bits_data_src2_T_9 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_out_bits_data_src2_T_14 = _io_out_bits_data_src2_T_10 | _io_out_bits_data_src2_T_11; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_out_bits_data_src2_T_15 = _io_out_bits_data_src2_T_14 | _io_out_bits_data_src2_T_12; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _wbClearMask_T_3 = io_wb_rfDest != 5'h0 & io_wb_rfDest == io_forward_wb_rfDest & forwardRfWen; // @[src/main/scala/nutcore/backend/seq/ISU.scala 41:100]
  wire [62:0] _wbClearMask_T_6 = 63'h1 << io_wb_rfDest; // @[src/main/scala/nutcore/RF.scala 38:39]
  wire [31:0] wbClearMask = io_wb_rfWen & ~_wbClearMask_T_3 ? _wbClearMask_T_6[31:0] : 32'h0; // @[src/main/scala/nutcore/backend/seq/ISU.scala 85:24]
  wire  _isuFireSetMask_T = io_out_ready & io_out_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  wire [62:0] _isuFireSetMask_T_1 = 63'h1 << io_in_0_bits_ctrl_rfDest; // @[src/main/scala/nutcore/RF.scala 38:39]
  wire [31:0] isuFireSetMask = _isuFireSetMask_T ? _isuFireSetMask_T_1[31:0] : 32'h0; // @[src/main/scala/nutcore/backend/seq/ISU.scala 87:27]
  wire [31:0] _busy_T_5 = ~wbClearMask; // @[src/main/scala/nutcore/RF.scala 44:26]
  wire [31:0] _busy_T_6 = busy & _busy_T_5; // @[src/main/scala/nutcore/RF.scala 44:24]
  wire [31:0] _busy_T_7 = _busy_T_6 | isuFireSetMask; // @[src/main/scala/nutcore/RF.scala 44:38]
  wire [31:0] _busy_T_9 = {_busy_T_7[31:1],1'h0}; // @[src/main/scala/nutcore/RF.scala 44:16]
  reg [63:0] c; // @[src/main/scala/utils/GTimer.scala 24:20]
  wire [63:0] _c_T_1 = c + 64'h1; // @[src/main/scala/utils/GTimer.scala 25:12]
  wire  _T_3 = _isuFireSetMask_T & DISPLAY_ENABLE; // @[src/main/scala/utils/Debug.scala 55:16]
  wire  _T_5 = ~reset; // @[src/main/scala/utils/Debug.scala 56:24]
  wire  _WIRE = io_in_0_valid & ~io_out_valid; // @[src/main/scala/nutcore/backend/seq/ISU.scala 97:49]
  wire  _WIRE_1 = io_out_valid & ~_isuFireSetMask_T; // @[src/main/scala/nutcore/backend/seq/ISU.scala 98:47]
  wire  _WIRE_2 = io_out_ready & io_out_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  assign rf_io_out_bits_data_src1_MPORT_en = 1'h1;
  assign rf_io_out_bits_data_src1_MPORT_addr = io_in_0_bits_ctrl_rfSrc1;
  assign rf_io_out_bits_data_src1_MPORT_data = rf[rf_io_out_bits_data_src1_MPORT_addr]; // @[src/main/scala/nutcore/RF.scala 30:15]
  assign rf_io_out_bits_data_src2_MPORT_en = 1'h1;
  assign rf_io_out_bits_data_src2_MPORT_addr = io_in_0_bits_ctrl_rfSrc2;
  assign rf_io_out_bits_data_src2_MPORT_data = rf[rf_io_out_bits_data_src2_MPORT_addr]; // @[src/main/scala/nutcore/RF.scala 30:15]
  assign rf_MPORT_1_en = 1'h1;
  assign rf_MPORT_1_addr = 5'h0;
  assign rf_MPORT_1_data = rf[rf_MPORT_1_addr]; // @[src/main/scala/nutcore/RF.scala 30:15]
  assign rf_MPORT_2_en = 1'h1;
  assign rf_MPORT_2_addr = 5'h1;
  assign rf_MPORT_2_data = rf[rf_MPORT_2_addr]; // @[src/main/scala/nutcore/RF.scala 30:15]
  assign rf_MPORT_3_en = 1'h1;
  assign rf_MPORT_3_addr = 5'h2;
  assign rf_MPORT_3_data = rf[rf_MPORT_3_addr]; // @[src/main/scala/nutcore/RF.scala 30:15]
  assign rf_MPORT_4_en = 1'h1;
  assign rf_MPORT_4_addr = 5'h3;
  assign rf_MPORT_4_data = rf[rf_MPORT_4_addr]; // @[src/main/scala/nutcore/RF.scala 30:15]
  assign rf_MPORT_5_en = 1'h1;
  assign rf_MPORT_5_addr = 5'h4;
  assign rf_MPORT_5_data = rf[rf_MPORT_5_addr]; // @[src/main/scala/nutcore/RF.scala 30:15]
  assign rf_MPORT_6_en = 1'h1;
  assign rf_MPORT_6_addr = 5'h5;
  assign rf_MPORT_6_data = rf[rf_MPORT_6_addr]; // @[src/main/scala/nutcore/RF.scala 30:15]
  assign rf_MPORT_7_en = 1'h1;
  assign rf_MPORT_7_addr = 5'h6;
  assign rf_MPORT_7_data = rf[rf_MPORT_7_addr]; // @[src/main/scala/nutcore/RF.scala 30:15]
  assign rf_MPORT_8_en = 1'h1;
  assign rf_MPORT_8_addr = 5'h7;
  assign rf_MPORT_8_data = rf[rf_MPORT_8_addr]; // @[src/main/scala/nutcore/RF.scala 30:15]
  assign rf_MPORT_9_en = 1'h1;
  assign rf_MPORT_9_addr = 5'h8;
  assign rf_MPORT_9_data = rf[rf_MPORT_9_addr]; // @[src/main/scala/nutcore/RF.scala 30:15]
  assign rf_MPORT_10_en = 1'h1;
  assign rf_MPORT_10_addr = 5'h9;
  assign rf_MPORT_10_data = rf[rf_MPORT_10_addr]; // @[src/main/scala/nutcore/RF.scala 30:15]
  assign rf_MPORT_11_en = 1'h1;
  assign rf_MPORT_11_addr = 5'ha;
  assign rf_MPORT_11_data = rf[rf_MPORT_11_addr]; // @[src/main/scala/nutcore/RF.scala 30:15]
  assign rf_MPORT_12_en = 1'h1;
  assign rf_MPORT_12_addr = 5'hb;
  assign rf_MPORT_12_data = rf[rf_MPORT_12_addr]; // @[src/main/scala/nutcore/RF.scala 30:15]
  assign rf_MPORT_13_en = 1'h1;
  assign rf_MPORT_13_addr = 5'hc;
  assign rf_MPORT_13_data = rf[rf_MPORT_13_addr]; // @[src/main/scala/nutcore/RF.scala 30:15]
  assign rf_MPORT_14_en = 1'h1;
  assign rf_MPORT_14_addr = 5'hd;
  assign rf_MPORT_14_data = rf[rf_MPORT_14_addr]; // @[src/main/scala/nutcore/RF.scala 30:15]
  assign rf_MPORT_15_en = 1'h1;
  assign rf_MPORT_15_addr = 5'he;
  assign rf_MPORT_15_data = rf[rf_MPORT_15_addr]; // @[src/main/scala/nutcore/RF.scala 30:15]
  assign rf_MPORT_16_en = 1'h1;
  assign rf_MPORT_16_addr = 5'hf;
  assign rf_MPORT_16_data = rf[rf_MPORT_16_addr]; // @[src/main/scala/nutcore/RF.scala 30:15]
  assign rf_MPORT_17_en = 1'h1;
  assign rf_MPORT_17_addr = 5'h10;
  assign rf_MPORT_17_data = rf[rf_MPORT_17_addr]; // @[src/main/scala/nutcore/RF.scala 30:15]
  assign rf_MPORT_18_en = 1'h1;
  assign rf_MPORT_18_addr = 5'h11;
  assign rf_MPORT_18_data = rf[rf_MPORT_18_addr]; // @[src/main/scala/nutcore/RF.scala 30:15]
  assign rf_MPORT_19_en = 1'h1;
  assign rf_MPORT_19_addr = 5'h12;
  assign rf_MPORT_19_data = rf[rf_MPORT_19_addr]; // @[src/main/scala/nutcore/RF.scala 30:15]
  assign rf_MPORT_20_en = 1'h1;
  assign rf_MPORT_20_addr = 5'h13;
  assign rf_MPORT_20_data = rf[rf_MPORT_20_addr]; // @[src/main/scala/nutcore/RF.scala 30:15]
  assign rf_MPORT_21_en = 1'h1;
  assign rf_MPORT_21_addr = 5'h14;
  assign rf_MPORT_21_data = rf[rf_MPORT_21_addr]; // @[src/main/scala/nutcore/RF.scala 30:15]
  assign rf_MPORT_22_en = 1'h1;
  assign rf_MPORT_22_addr = 5'h15;
  assign rf_MPORT_22_data = rf[rf_MPORT_22_addr]; // @[src/main/scala/nutcore/RF.scala 30:15]
  assign rf_MPORT_23_en = 1'h1;
  assign rf_MPORT_23_addr = 5'h16;
  assign rf_MPORT_23_data = rf[rf_MPORT_23_addr]; // @[src/main/scala/nutcore/RF.scala 30:15]
  assign rf_MPORT_24_en = 1'h1;
  assign rf_MPORT_24_addr = 5'h17;
  assign rf_MPORT_24_data = rf[rf_MPORT_24_addr]; // @[src/main/scala/nutcore/RF.scala 30:15]
  assign rf_MPORT_25_en = 1'h1;
  assign rf_MPORT_25_addr = 5'h18;
  assign rf_MPORT_25_data = rf[rf_MPORT_25_addr]; // @[src/main/scala/nutcore/RF.scala 30:15]
  assign rf_MPORT_26_en = 1'h1;
  assign rf_MPORT_26_addr = 5'h19;
  assign rf_MPORT_26_data = rf[rf_MPORT_26_addr]; // @[src/main/scala/nutcore/RF.scala 30:15]
  assign rf_MPORT_27_en = 1'h1;
  assign rf_MPORT_27_addr = 5'h1a;
  assign rf_MPORT_27_data = rf[rf_MPORT_27_addr]; // @[src/main/scala/nutcore/RF.scala 30:15]
  assign rf_MPORT_28_en = 1'h1;
  assign rf_MPORT_28_addr = 5'h1b;
  assign rf_MPORT_28_data = rf[rf_MPORT_28_addr]; // @[src/main/scala/nutcore/RF.scala 30:15]
  assign rf_MPORT_29_en = 1'h1;
  assign rf_MPORT_29_addr = 5'h1c;
  assign rf_MPORT_29_data = rf[rf_MPORT_29_addr]; // @[src/main/scala/nutcore/RF.scala 30:15]
  assign rf_MPORT_30_en = 1'h1;
  assign rf_MPORT_30_addr = 5'h1d;
  assign rf_MPORT_30_data = rf[rf_MPORT_30_addr]; // @[src/main/scala/nutcore/RF.scala 30:15]
  assign rf_MPORT_31_en = 1'h1;
  assign rf_MPORT_31_addr = 5'h1e;
  assign rf_MPORT_31_data = rf[rf_MPORT_31_addr]; // @[src/main/scala/nutcore/RF.scala 30:15]
  assign rf_MPORT_32_en = 1'h1;
  assign rf_MPORT_32_addr = 5'h1f;
  assign rf_MPORT_32_data = rf[rf_MPORT_32_addr]; // @[src/main/scala/nutcore/RF.scala 30:15]
  assign rf_MPORT_data = io_wb_rfData;
  assign rf_MPORT_addr = io_wb_rfDest;
  assign rf_MPORT_mask = 1'h1;
  assign rf_MPORT_en = io_wb_rfWen;
  assign io_in_0_ready = ~io_in_0_valid | _isuFireSetMask_T; // @[src/main/scala/nutcore/backend/seq/ISU.scala 91:37]
  assign io_out_valid = io_in_0_valid & src1Ready & src2Ready; // @[src/main/scala/nutcore/backend/seq/ISU.scala 58:47]
  assign io_out_bits_cf_instr = io_in_0_bits_cf_instr; // @[src/main/scala/nutcore/backend/seq/ISU.scala 77:18]
  assign io_out_bits_cf_pc = io_in_0_bits_cf_pc; // @[src/main/scala/nutcore/backend/seq/ISU.scala 77:18]
  assign io_out_bits_cf_pnpc = io_in_0_bits_cf_pnpc; // @[src/main/scala/nutcore/backend/seq/ISU.scala 77:18]
  assign io_out_bits_cf_exceptionVec_1 = io_in_0_bits_cf_exceptionVec_1; // @[src/main/scala/nutcore/backend/seq/ISU.scala 77:18]
  assign io_out_bits_cf_exceptionVec_2 = io_in_0_bits_cf_exceptionVec_2; // @[src/main/scala/nutcore/backend/seq/ISU.scala 77:18]
  assign io_out_bits_cf_exceptionVec_12 = io_in_0_bits_cf_exceptionVec_12; // @[src/main/scala/nutcore/backend/seq/ISU.scala 77:18]
  assign io_out_bits_cf_intrVec_0 = io_in_0_bits_cf_intrVec_0; // @[src/main/scala/nutcore/backend/seq/ISU.scala 77:18]
  assign io_out_bits_cf_intrVec_1 = io_in_0_bits_cf_intrVec_1; // @[src/main/scala/nutcore/backend/seq/ISU.scala 77:18]
  assign io_out_bits_cf_intrVec_2 = io_in_0_bits_cf_intrVec_2; // @[src/main/scala/nutcore/backend/seq/ISU.scala 77:18]
  assign io_out_bits_cf_intrVec_3 = io_in_0_bits_cf_intrVec_3; // @[src/main/scala/nutcore/backend/seq/ISU.scala 77:18]
  assign io_out_bits_cf_intrVec_4 = io_in_0_bits_cf_intrVec_4; // @[src/main/scala/nutcore/backend/seq/ISU.scala 77:18]
  assign io_out_bits_cf_intrVec_5 = io_in_0_bits_cf_intrVec_5; // @[src/main/scala/nutcore/backend/seq/ISU.scala 77:18]
  assign io_out_bits_cf_intrVec_6 = io_in_0_bits_cf_intrVec_6; // @[src/main/scala/nutcore/backend/seq/ISU.scala 77:18]
  assign io_out_bits_cf_intrVec_7 = io_in_0_bits_cf_intrVec_7; // @[src/main/scala/nutcore/backend/seq/ISU.scala 77:18]
  assign io_out_bits_cf_intrVec_8 = io_in_0_bits_cf_intrVec_8; // @[src/main/scala/nutcore/backend/seq/ISU.scala 77:18]
  assign io_out_bits_cf_intrVec_9 = io_in_0_bits_cf_intrVec_9; // @[src/main/scala/nutcore/backend/seq/ISU.scala 77:18]
  assign io_out_bits_cf_intrVec_10 = io_in_0_bits_cf_intrVec_10; // @[src/main/scala/nutcore/backend/seq/ISU.scala 77:18]
  assign io_out_bits_cf_intrVec_11 = io_in_0_bits_cf_intrVec_11; // @[src/main/scala/nutcore/backend/seq/ISU.scala 77:18]
  assign io_out_bits_cf_brIdx = io_in_0_bits_cf_brIdx; // @[src/main/scala/nutcore/backend/seq/ISU.scala 77:18]
  assign io_out_bits_cf_crossPageIPFFix = io_in_0_bits_cf_crossPageIPFFix; // @[src/main/scala/nutcore/backend/seq/ISU.scala 77:18]
  assign io_out_bits_ctrl_fuType = io_in_0_bits_ctrl_fuType; // @[src/main/scala/nutcore/backend/seq/ISU.scala 78:20]
  assign io_out_bits_ctrl_fuOpType = io_in_0_bits_ctrl_fuOpType; // @[src/main/scala/nutcore/backend/seq/ISU.scala 78:20]
  assign io_out_bits_ctrl_rfWen = io_in_0_bits_ctrl_rfWen; // @[src/main/scala/nutcore/backend/seq/ISU.scala 78:20]
  assign io_out_bits_ctrl_rfDest = io_in_0_bits_ctrl_rfDest; // @[src/main/scala/nutcore/backend/seq/ISU.scala 78:20]
  assign io_out_bits_ctrl_isNutCoreTrap = io_in_0_bits_ctrl_isNutCoreTrap; // @[src/main/scala/nutcore/backend/seq/ISU.scala 78:20]
  assign io_out_bits_data_src1 = _io_out_bits_data_src1_T_18 | _io_out_bits_data_src1_T_16; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign io_out_bits_data_src2 = _io_out_bits_data_src2_T_15 | _io_out_bits_data_src2_T_13; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign io_out_bits_data_imm = io_in_0_bits_data_imm; // @[src/main/scala/nutcore/backend/seq/ISU.scala 75:25]
  assign _WIRE_1_0 = _WIRE_1;
  assign _WIRE_8 = _WIRE;
  assign _WIRE_2_2 = _WIRE_2;
  always @(posedge clock) begin
    if (rf_MPORT_en & rf_MPORT_mask) begin
      rf[rf_MPORT_addr] <= rf_MPORT_data; // @[src/main/scala/nutcore/RF.scala 30:15]
    end
    if (reset) begin // @[src/main/scala/nutcore/RF.scala 36:21]
      busy <= 32'h0; // @[src/main/scala/nutcore/RF.scala 36:21]
    end else if (io_flush) begin // @[src/main/scala/nutcore/backend/seq/ISU.scala 88:19]
      busy <= 32'h0; // @[src/main/scala/nutcore/RF.scala 44:10]
    end else begin
      busy <= _busy_T_9; // @[src/main/scala/nutcore/RF.scala 44:10]
    end
    if (reset) begin // @[src/main/scala/utils/GTimer.scala 24:20]
      c <= 64'h0; // @[src/main/scala/utils/GTimer.scala 24:20]
    end else begin
      c <= _c_T_1; // @[src/main/scala/utils/GTimer.scala 25:7]
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3 & ~reset) begin
          $fwrite(32'h80000002,"[%d] ISU: ",c); // @[src/main/scala/utils/Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3 & _T_5) begin
          $fwrite(32'h80000002,"issue: pc %x npc %x instr %x src1 %x src2 %x imm %x\n",io_out_bits_cf_pc,
            io_out_bits_cf_pnpc,io_out_bits_cf_instr,io_out_bits_data_src1,io_out_bits_data_src2,io_out_bits_data_imm); // @[src/main/scala/utils/Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {2{`RANDOM}};
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    rf[initvar] = _RAND_0[63:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  busy = _RAND_1[31:0];
  _RAND_2 = {2{`RANDOM}};
  c = _RAND_2[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ALU(
  input         clock,
  input         reset,
  input         io_in_valid, // @[src/main/scala/nutcore/backend/fu/ALU.scala 76:14]
  input  [63:0] io_in_bits_src1, // @[src/main/scala/nutcore/backend/fu/ALU.scala 76:14]
  input  [63:0] io_in_bits_src2, // @[src/main/scala/nutcore/backend/fu/ALU.scala 76:14]
  input  [6:0]  io_in_bits_func, // @[src/main/scala/nutcore/backend/fu/ALU.scala 76:14]
  input         io_out_ready, // @[src/main/scala/nutcore/backend/fu/ALU.scala 76:14]
  output        io_out_valid, // @[src/main/scala/nutcore/backend/fu/ALU.scala 76:14]
  output [63:0] io_out_bits, // @[src/main/scala/nutcore/backend/fu/ALU.scala 76:14]
  input  [63:0] io_cfIn_instr, // @[src/main/scala/nutcore/backend/fu/ALU.scala 76:14]
  input  [38:0] io_cfIn_pc, // @[src/main/scala/nutcore/backend/fu/ALU.scala 76:14]
  input  [38:0] io_cfIn_pnpc, // @[src/main/scala/nutcore/backend/fu/ALU.scala 76:14]
  input  [3:0]  io_cfIn_brIdx, // @[src/main/scala/nutcore/backend/fu/ALU.scala 76:14]
  output [38:0] io_redirect_target, // @[src/main/scala/nutcore/backend/fu/ALU.scala 76:14]
  output        io_redirect_valid, // @[src/main/scala/nutcore/backend/fu/ALU.scala 76:14]
  input  [63:0] io_offset, // @[src/main/scala/nutcore/backend/fu/ALU.scala 76:14]
  output        _WIRE_2_0,
  output        REG_0_valid,
  output [38:0] REG_0_pc,
  output        REG_0_isMissPredict,
  output [38:0] REG_0_actualTarget,
  output        REG_0_actualTaken,
  output [6:0]  REG_0_fuOpType,
  output [1:0]  REG_0_btbType,
  output        REG_0_isRVC,
  output        _WIRE_15_0,
  input         DISPLAY_ENABLE,
  output        _WIRE_13_0,
  output        _WIRE_6_0,
  output        _WIRE_5_0,
  output        _WIRE_4_1,
  output        _WIRE_3_0,
  output        _WIRE_10_0,
  output        _WIRE_9_0,
  output        _WIRE_8_0,
  output        _WIRE_7_0,
  output        _WIRE_1_2,
  output        _WIRE_12_0,
  output        _WIRE_14_0,
  output        _WIRE_11_0,
  output        _WIRE_16_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
`endif // RANDOMIZE_REG_INIT
  wire  isAdderSub = ~io_in_bits_func[6]; // @[src/main/scala/nutcore/backend/fu/ALU.scala 87:20]
  wire [63:0] _adderRes_T_1 = isAdderSub ? 64'hffffffffffffffff : 64'h0; // @[src/main/scala/nutcore/backend/fu/ALU.scala 88:39]
  wire [63:0] _adderRes_T_2 = io_in_bits_src2 ^ _adderRes_T_1; // @[src/main/scala/nutcore/backend/fu/ALU.scala 88:33]
  wire [64:0] _adderRes_T_3 = io_in_bits_src1 + _adderRes_T_2; // @[src/main/scala/nutcore/backend/fu/ALU.scala 88:24]
  wire [64:0] _GEN_0 = {{64'd0}, isAdderSub}; // @[src/main/scala/nutcore/backend/fu/ALU.scala 88:60]
  wire [64:0] adderRes = _adderRes_T_3 + _GEN_0; // @[src/main/scala/nutcore/backend/fu/ALU.scala 88:60]
  wire [63:0] xorRes = io_in_bits_src1 ^ io_in_bits_src2; // @[src/main/scala/nutcore/backend/fu/ALU.scala 89:21]
  wire  sltu = ~adderRes[64]; // @[src/main/scala/nutcore/backend/fu/ALU.scala 90:14]
  wire  slt = xorRes[63] ^ sltu; // @[src/main/scala/nutcore/backend/fu/ALU.scala 91:28]
  wire [63:0] _shsrc1_T_2 = {32'h0,io_in_bits_src1[31:0]}; // @[src/main/scala/utils/BitUtils.scala 49:41]
  wire  shsrc1_signBit = io_in_bits_src1[31]; // @[src/main/scala/utils/BitUtils.scala 41:20]
  wire [31:0] _shsrc1_T_5 = shsrc1_signBit ? 32'hffffffff : 32'h0; // @[src/main/scala/utils/BitUtils.scala 42:46]
  wire [63:0] _shsrc1_T_6 = {_shsrc1_T_5,io_in_bits_src1[31:0]}; // @[src/main/scala/utils/BitUtils.scala 42:41]
  wire [63:0] _shsrc1_T_8 = 7'h25 == io_in_bits_func ? _shsrc1_T_2 : io_in_bits_src1; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [63:0] shsrc1 = 7'h2d == io_in_bits_func ? _shsrc1_T_6 : _shsrc1_T_8; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [5:0] shamt = io_in_bits_func[5] ? {{1'd0}, io_in_bits_src2[4:0]} : io_in_bits_src2[5:0]; // @[src/main/scala/nutcore/backend/fu/ALU.scala 97:18]
  wire [126:0] _GEN_4 = {{63'd0}, shsrc1}; // @[src/main/scala/nutcore/backend/fu/ALU.scala 99:33]
  wire [126:0] _res_T_1 = _GEN_4 << shamt; // @[src/main/scala/nutcore/backend/fu/ALU.scala 99:33]
  wire [63:0] _res_T_3 = {63'h0,slt}; // @[src/main/scala/utils/BitUtils.scala 49:41]
  wire [63:0] _res_T_4 = {63'h0,sltu}; // @[src/main/scala/utils/BitUtils.scala 49:41]
  wire [63:0] _res_T_5 = shsrc1 >> shamt; // @[src/main/scala/nutcore/backend/fu/ALU.scala 103:32]
  wire [63:0] _res_T_6 = io_in_bits_src1 | io_in_bits_src2; // @[src/main/scala/nutcore/backend/fu/ALU.scala 104:30]
  wire [63:0] _res_T_7 = io_in_bits_src1 & io_in_bits_src2; // @[src/main/scala/nutcore/backend/fu/ALU.scala 105:30]
  wire [63:0] _res_T_8 = 7'h2d == io_in_bits_func ? _shsrc1_T_6 : _shsrc1_T_8; // @[src/main/scala/nutcore/backend/fu/ALU.scala 106:32]
  wire [63:0] _res_T_10 = $signed(_res_T_8) >>> shamt; // @[src/main/scala/nutcore/backend/fu/ALU.scala 106:49]
  wire [64:0] _res_T_12 = 4'h1 == io_in_bits_func[3:0] ? {{1'd0}, _res_T_1[63:0]} : adderRes; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [64:0] _res_T_14 = 4'h2 == io_in_bits_func[3:0] ? {{1'd0}, _res_T_3} : _res_T_12; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [64:0] _res_T_16 = 4'h3 == io_in_bits_func[3:0] ? {{1'd0}, _res_T_4} : _res_T_14; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [64:0] _res_T_18 = 4'h4 == io_in_bits_func[3:0] ? {{1'd0}, xorRes} : _res_T_16; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [64:0] _res_T_20 = 4'h5 == io_in_bits_func[3:0] ? {{1'd0}, _res_T_5} : _res_T_18; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [64:0] _res_T_22 = 4'h6 == io_in_bits_func[3:0] ? {{1'd0}, _res_T_6} : _res_T_20; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [64:0] _res_T_24 = 4'h7 == io_in_bits_func[3:0] ? {{1'd0}, _res_T_7} : _res_T_22; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [64:0] res = 4'hd == io_in_bits_func[3:0] ? {{1'd0}, _res_T_10} : _res_T_24; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  aluRes_signBit = res[31]; // @[src/main/scala/utils/BitUtils.scala 41:20]
  wire [31:0] _aluRes_T_3 = aluRes_signBit ? 32'hffffffff : 32'h0; // @[src/main/scala/utils/BitUtils.scala 42:46]
  wire [63:0] _aluRes_T_4 = {_aluRes_T_3,res[31:0]}; // @[src/main/scala/utils/BitUtils.scala 42:41]
  wire [64:0] aluRes = io_in_bits_func[5] ? {{1'd0}, _aluRes_T_4} : res; // @[src/main/scala/nutcore/backend/fu/ALU.scala 108:19]
  wire  _T_1 = ~(|xorRes); // @[src/main/scala/nutcore/backend/fu/ALU.scala 111:48]
  wire  isBranch = ~io_in_bits_func[3]; // @[src/main/scala/nutcore/backend/fu/ALU.scala 63:30]
  wire  isBru = io_in_bits_func[4]; // @[src/main/scala/nutcore/backend/fu/ALU.scala 62:31]
  wire  _taken_T_1 = 2'h0 == io_in_bits_func[2:1]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _taken_T_2 = 2'h2 == io_in_bits_func[2:1]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _taken_T_3 = 2'h3 == io_in_bits_func[2:1]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _taken_T_8 = _taken_T_1 & _T_1 | _taken_T_2 & slt | _taken_T_3 & sltu; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  taken = _taken_T_8 ^ io_in_bits_func[0]; // @[src/main/scala/nutcore/backend/fu/ALU.scala 118:72]
  wire [63:0] _GEN_1 = {{25'd0}, io_cfIn_pc}; // @[src/main/scala/nutcore/backend/fu/ALU.scala 119:41]
  wire [63:0] _target_T_1 = _GEN_1 + io_offset; // @[src/main/scala/nutcore/backend/fu/ALU.scala 119:41]
  wire [64:0] _target_T_2 = isBranch ? {{1'd0}, _target_T_1} : adderRes; // @[src/main/scala/nutcore/backend/fu/ALU.scala 119:19]
  wire [38:0] target = _target_T_2[38:0]; // @[src/main/scala/nutcore/backend/fu/ALU.scala 119:63]
  wire  _predictWrong_T_1 = ~taken & isBranch; // @[src/main/scala/nutcore/backend/fu/ALU.scala 120:33]
  wire  predictWrong = ~taken & isBranch ? io_cfIn_brIdx[0] : ~io_cfIn_brIdx[0] | io_redirect_target != io_cfIn_pnpc; // @[src/main/scala/nutcore/backend/fu/ALU.scala 120:25]
  wire  isRVC = io_cfIn_instr[1:0] != 2'h3; // @[src/main/scala/nutcore/backend/fu/ALU.scala 121:35]
  wire  _T_3 = io_cfIn_instr[1:0] == 2'h3; // @[src/main/scala/nutcore/backend/fu/ALU.scala 122:29]
  wire  _T_8 = ~reset; // @[src/main/scala/nutcore/backend/fu/ALU.scala 122:9]
  wire  _T_12 = ~isRVC; // @[src/main/scala/nutcore/backend/fu/ALU.scala 123:55]
  wire  _T_14 = io_in_valid & _T_3 != ~isRVC; // @[src/main/scala/nutcore/backend/fu/ALU.scala 123:15]
  reg [63:0] c; // @[src/main/scala/utils/GTimer.scala 24:20]
  wire [63:0] _c_T_1 = c + 64'h1; // @[src/main/scala/utils/GTimer.scala 25:12]
  wire  _T_15 = _T_14 & DISPLAY_ENABLE; // @[src/main/scala/utils/Debug.scala 55:16]
  wire [38:0] _io_redirect_target_T_3 = io_cfIn_pc + 39'h2; // @[src/main/scala/nutcore/backend/fu/ALU.scala 124:71]
  wire [38:0] _io_redirect_target_T_5 = io_cfIn_pc + 39'h4; // @[src/main/scala/nutcore/backend/fu/ALU.scala 124:89]
  wire [38:0] _io_redirect_target_T_6 = isRVC ? _io_redirect_target_T_3 : _io_redirect_target_T_5; // @[src/main/scala/nutcore/backend/fu/ALU.scala 124:52]
  wire  _io_redirect_valid_T = io_in_valid & isBru; // @[src/main/scala/nutcore/backend/fu/ALU.scala 126:30]
  wire  _io_redirect_valid_T_1 = io_in_valid & isBru & predictWrong; // @[src/main/scala/nutcore/backend/fu/ALU.scala 126:39]
  wire  io_out_bits_signBit = io_cfIn_pc[38]; // @[src/main/scala/utils/BitUtils.scala 41:20]
  wire [24:0] _io_out_bits_T_2 = io_out_bits_signBit ? 25'h1ffffff : 25'h0; // @[src/main/scala/utils/BitUtils.scala 42:46]
  wire [63:0] _io_out_bits_T_3 = {_io_out_bits_T_2,io_cfIn_pc}; // @[src/main/scala/utils/BitUtils.scala 42:41]
  wire [63:0] _io_out_bits_T_5 = _io_out_bits_T_3 + 64'h4; // @[src/main/scala/nutcore/backend/fu/ALU.scala 132:71]
  wire [63:0] _io_out_bits_T_10 = _io_out_bits_T_3 + 64'h2; // @[src/main/scala/nutcore/backend/fu/ALU.scala 132:108]
  wire [63:0] _io_out_bits_T_11 = _T_12 ? _io_out_bits_T_5 : _io_out_bits_T_10; // @[src/main/scala/nutcore/backend/fu/ALU.scala 132:32]
  wire [64:0] _io_out_bits_T_12 = isBru ? {{1'd0}, _io_out_bits_T_11} : aluRes; // @[src/main/scala/nutcore/backend/fu/ALU.scala 132:21]
  reg [63:0] c_1; // @[src/main/scala/utils/GTimer.scala 24:20]
  wire [63:0] _c_T_3 = c_1 + 64'h1; // @[src/main/scala/utils/GTimer.scala 25:12]
  wire  _T_21 = _io_redirect_valid_T & DISPLAY_ENABLE; // @[src/main/scala/utils/Debug.scala 55:16]
  reg [63:0] c_2; // @[src/main/scala/utils/GTimer.scala 24:20]
  wire [63:0] _c_T_5 = c_2 + 64'h1; // @[src/main/scala/utils/GTimer.scala 25:12]
  wire  _T_35 = io_in_bits_func == 7'h58 | io_in_bits_func == 7'h5c; // @[src/main/scala/nutcore/backend/fu/ALU.scala 136:180]
  wire  _T_36 = io_in_bits_func == 7'h5a; // @[src/main/scala/nutcore/backend/fu/ALU.scala 136:214]
  wire  _T_37 = io_in_bits_func == 7'h5e; // @[src/main/scala/nutcore/backend/fu/ALU.scala 136:239]
  reg [63:0] c_3; // @[src/main/scala/utils/GTimer.scala 24:20]
  wire [63:0] _c_T_7 = c_3 + 64'h1; // @[src/main/scala/utils/GTimer.scala 25:12]
  reg [63:0] c_4; // @[src/main/scala/utils/GTimer.scala 24:20]
  wire [63:0] _c_T_9 = c_4 + 64'h1; // @[src/main/scala/utils/GTimer.scala 25:12]
  wire  _T_56 = 7'h5c == io_in_bits_func; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _T_57 = 7'h5e == io_in_bits_func; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _T_58 = 7'h58 == io_in_bits_func; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _T_59 = 7'h5a == io_in_bits_func; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [1:0] _T_67 = _T_57 ? 2'h3 : 2'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [1:0] _T_69 = _T_59 ? 2'h2 : 2'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [1:0] _GEN_2 = {{1'd0}, _T_56}; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [1:0] _T_76 = _GEN_2 | _T_67; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [1:0] _GEN_3 = {{1'd0}, _T_58}; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [1:0] _T_77 = _T_76 | _GEN_3; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [1:0] _T_78 = _T_77 | _T_69; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  reg [63:0] c_5; // @[src/main/scala/utils/GTimer.scala 24:20]
  wire [63:0] _c_T_11 = c_5 + 64'h1; // @[src/main/scala/utils/GTimer.scala 25:12]
  reg  REG_valid; // @[src/main/scala/nutcore/backend/fu/ALU.scala 159:34]
  reg [38:0] REG_pc; // @[src/main/scala/nutcore/backend/fu/ALU.scala 159:34]
  reg  REG_isMissPredict; // @[src/main/scala/nutcore/backend/fu/ALU.scala 159:34]
  reg [38:0] REG_actualTarget; // @[src/main/scala/nutcore/backend/fu/ALU.scala 159:34]
  reg  REG_actualTaken; // @[src/main/scala/nutcore/backend/fu/ALU.scala 159:34]
  reg [6:0] REG_fuOpType; // @[src/main/scala/nutcore/backend/fu/ALU.scala 159:34]
  reg [1:0] REG_btbType; // @[src/main/scala/nutcore/backend/fu/ALU.scala 159:34]
  reg  REG_isRVC; // @[src/main/scala/nutcore/backend/fu/ALU.scala 159:34]
  wire  right = _io_redirect_valid_T & ~predictWrong; // @[src/main/scala/nutcore/backend/fu/ALU.scala 161:32]
  wire  _T_85 = _io_redirect_valid_T_1 & isBranch; // @[src/main/scala/nutcore/backend/fu/ALU.scala 164:42]
  wire  _T_89 = _T_85 & io_cfIn_pc[2:0] == 3'h0; // @[src/main/scala/nutcore/backend/fu/ALU.scala 165:54]
  wire  _T_100 = _T_85 & io_cfIn_pc[2:0] == 3'h2; // @[src/main/scala/nutcore/backend/fu/ALU.scala 167:54]
  wire  _T_111 = _T_85 & io_cfIn_pc[2:0] == 3'h4; // @[src/main/scala/nutcore/backend/fu/ALU.scala 169:54]
  wire  _T_122 = _T_85 & io_cfIn_pc[2:0] == 3'h6; // @[src/main/scala/nutcore/backend/fu/ALU.scala 171:54]
  wire  _WIRE_1 = right & isBranch; // @[src/main/scala/nutcore/backend/fu/ALU.scala 163:42]
  wire  _WIRE_2 = _io_redirect_valid_T_1 & isBranch; // @[src/main/scala/nutcore/backend/fu/ALU.scala 164:42]
  wire  _WIRE_3 = _T_85 & io_cfIn_pc[2:0] == 3'h0 & isRVC; // @[src/main/scala/nutcore/backend/fu/ALU.scala 165:82]
  wire  _WIRE_4 = _T_89 & _T_12; // @[src/main/scala/nutcore/backend/fu/ALU.scala 166:82]
  wire  _WIRE_5 = _T_85 & io_cfIn_pc[2:0] == 3'h2 & isRVC; // @[src/main/scala/nutcore/backend/fu/ALU.scala 167:82]
  wire  _WIRE_6 = _T_100 & _T_12; // @[src/main/scala/nutcore/backend/fu/ALU.scala 168:82]
  wire  _WIRE_7 = _T_85 & io_cfIn_pc[2:0] == 3'h4 & isRVC; // @[src/main/scala/nutcore/backend/fu/ALU.scala 169:82]
  wire  _WIRE_8 = _T_111 & _T_12; // @[src/main/scala/nutcore/backend/fu/ALU.scala 170:82]
  wire  _WIRE_9 = _T_85 & io_cfIn_pc[2:0] == 3'h6 & isRVC; // @[src/main/scala/nutcore/backend/fu/ALU.scala 171:82]
  wire  _WIRE_10 = _T_122 & _T_12; // @[src/main/scala/nutcore/backend/fu/ALU.scala 172:82]
  wire  _WIRE_11 = right & _T_35; // @[src/main/scala/nutcore/backend/fu/ALU.scala 173:42]
  wire  _WIRE_12 = _io_redirect_valid_T_1 & _T_35; // @[src/main/scala/nutcore/backend/fu/ALU.scala 174:42]
  wire  _WIRE_13 = right & _T_36; // @[src/main/scala/nutcore/backend/fu/ALU.scala 175:42]
  wire  _WIRE_14 = _io_redirect_valid_T_1 & _T_36; // @[src/main/scala/nutcore/backend/fu/ALU.scala 176:42]
  wire  _WIRE_15 = right & _T_37; // @[src/main/scala/nutcore/backend/fu/ALU.scala 177:42]
  wire  _WIRE_16 = _io_redirect_valid_T_1 & _T_37; // @[src/main/scala/nutcore/backend/fu/ALU.scala 178:42]
  assign io_out_valid = io_in_valid; // @[src/main/scala/nutcore/backend/fu/ALU.scala 146:16]
  assign io_out_bits = _io_out_bits_T_12[63:0]; // @[src/main/scala/nutcore/backend/fu/ALU.scala 132:15]
  assign io_redirect_target = _predictWrong_T_1 ? _io_redirect_target_T_6 : target; // @[src/main/scala/nutcore/backend/fu/ALU.scala 124:28]
  assign io_redirect_valid = io_in_valid & isBru & predictWrong; // @[src/main/scala/nutcore/backend/fu/ALU.scala 126:39]
  assign _WIRE_2_0 = _WIRE_2;
  assign REG_0_valid = REG_valid;
  assign REG_0_pc = REG_pc;
  assign REG_0_isMissPredict = REG_isMissPredict;
  assign REG_0_actualTarget = REG_actualTarget;
  assign REG_0_actualTaken = REG_actualTaken;
  assign REG_0_fuOpType = REG_fuOpType;
  assign REG_0_btbType = REG_btbType;
  assign REG_0_isRVC = REG_isRVC;
  assign _WIRE_15_0 = _WIRE_15;
  assign _WIRE_13_0 = _WIRE_13;
  assign _WIRE_6_0 = _WIRE_6;
  assign _WIRE_5_0 = _WIRE_5;
  assign _WIRE_4_1 = _WIRE_4;
  assign _WIRE_3_0 = _WIRE_3;
  assign _WIRE_10_0 = _WIRE_10;
  assign _WIRE_9_0 = _WIRE_9;
  assign _WIRE_8_0 = _WIRE_8;
  assign _WIRE_7_0 = _WIRE_7;
  assign _WIRE_1_2 = _WIRE_1;
  assign _WIRE_12_0 = _WIRE_12;
  assign _WIRE_14_0 = _WIRE_14;
  assign _WIRE_11_0 = _WIRE_11;
  assign _WIRE_16_0 = _WIRE_16;
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/utils/GTimer.scala 24:20]
      c <= 64'h0; // @[src/main/scala/utils/GTimer.scala 24:20]
    end else begin
      c <= _c_T_1; // @[src/main/scala/utils/GTimer.scala 25:7]
    end
    if (reset) begin // @[src/main/scala/utils/GTimer.scala 24:20]
      c_1 <= 64'h0; // @[src/main/scala/utils/GTimer.scala 24:20]
    end else begin
      c_1 <= _c_T_3; // @[src/main/scala/utils/GTimer.scala 25:7]
    end
    if (reset) begin // @[src/main/scala/utils/GTimer.scala 24:20]
      c_2 <= 64'h0; // @[src/main/scala/utils/GTimer.scala 24:20]
    end else begin
      c_2 <= _c_T_5; // @[src/main/scala/utils/GTimer.scala 25:7]
    end
    if (reset) begin // @[src/main/scala/utils/GTimer.scala 24:20]
      c_3 <= 64'h0; // @[src/main/scala/utils/GTimer.scala 24:20]
    end else begin
      c_3 <= _c_T_7; // @[src/main/scala/utils/GTimer.scala 25:7]
    end
    if (reset) begin // @[src/main/scala/utils/GTimer.scala 24:20]
      c_4 <= 64'h0; // @[src/main/scala/utils/GTimer.scala 24:20]
    end else begin
      c_4 <= _c_T_9; // @[src/main/scala/utils/GTimer.scala 25:7]
    end
    if (reset) begin // @[src/main/scala/utils/GTimer.scala 24:20]
      c_5 <= 64'h0; // @[src/main/scala/utils/GTimer.scala 24:20]
    end else begin
      c_5 <= _c_T_11; // @[src/main/scala/utils/GTimer.scala 25:7]
    end
    REG_valid <= io_in_valid & isBru; // @[src/main/scala/nutcore/backend/fu/ALU.scala 149:31]
    REG_pc <= io_cfIn_pc; // @[src/main/scala/nutcore/backend/fu/ALU.scala 148:30 150:19]
    if (~taken & isBranch) begin // @[src/main/scala/nutcore/backend/fu/ALU.scala 120:25]
      REG_isMissPredict <= io_cfIn_brIdx[0];
    end else begin
      REG_isMissPredict <= ~io_cfIn_brIdx[0] | io_redirect_target != io_cfIn_pnpc;
    end
    REG_actualTarget <= _target_T_2[38:0]; // @[src/main/scala/nutcore/backend/fu/ALU.scala 119:63]
    REG_actualTaken <= _taken_T_8 ^ io_in_bits_func[0]; // @[src/main/scala/nutcore/backend/fu/ALU.scala 118:72]
    REG_fuOpType <= io_in_bits_func; // @[src/main/scala/nutcore/backend/fu/ALU.scala 148:30 154:25]
    REG_btbType <= _T_77 | _T_69; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
    REG_isRVC <= io_cfIn_instr[1:0] != 2'h3; // @[src/main/scala/nutcore/backend/fu/ALU.scala 121:35]
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_cfIn_instr[1:0] == 2'h3 | isRVC | ~io_in_valid)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ALU.scala:122 assert(io.cfIn.instr(1,0) === \"b11\".U || isRVC || !valid)\n"); // @[src/main/scala/nutcore/backend/fu/ALU.scala 122:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(io_cfIn_instr[1:0] == 2'h3 | isRVC | ~io_in_valid) & ~reset) begin
          $fatal; // @[src/main/scala/nutcore/backend/fu/ALU.scala 122:9]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_15 & _T_8) begin
          $fwrite(32'h80000002,"[%d] ALU: ",c); // @[src/main/scala/utils/Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_15 & _T_8) begin
          $fwrite(32'h80000002,"[ERROR] pc %x inst %x rvc %x\n",io_cfIn_pc,io_cfIn_instr,isRVC); // @[src/main/scala/utils/Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_21 & _T_8) begin
          $fwrite(32'h80000002,"[%d] ALU: ",c_1); // @[src/main/scala/utils/Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_21 & _T_8) begin
          $fwrite(32'h80000002,"tgt %x, valid:%d, npc: %x, pdwrong: %x\n",io_redirect_target,io_redirect_valid,
            io_cfIn_pnpc,predictWrong); // @[src/main/scala/utils/Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_21 & _T_8) begin
          $fwrite(32'h80000002,"[%d] ALU: ",c_2); // @[src/main/scala/utils/Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_21 & _T_8) begin
          $fwrite(32'h80000002,"taken:%d addrRes:%x src1:%x src2:%x func:%x\n",taken,adderRes,io_in_bits_src1,
            io_in_bits_src2,io_in_bits_func); // @[src/main/scala/utils/Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_21 & _T_8) begin
          $fwrite(32'h80000002,"[%d] ALU: ",c_3); // @[src/main/scala/utils/Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_21 & _T_8) begin
          $fwrite(32'h80000002,"[BPW] pc %x tgt %x, npc: %x, pdwrong: %x type: %x%x%x%x\n",io_cfIn_pc,io_redirect_target
            ,io_cfIn_pnpc,predictWrong,isBranch,_T_35,_T_36,_T_37); // @[src/main/scala/utils/Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_8) begin
          $fwrite(32'h80000002,"[%d] ALU: ",c_4); // @[src/main/scala/utils/Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_8) begin
          $fwrite(32'h80000002,"valid:%d isBru:%d isBranch:%d \n",io_in_valid,isBru,isBranch); // @[src/main/scala/utils/Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_21 & _T_8) begin
          $fwrite(32'h80000002,"[%d] ALU: ",c_5); // @[src/main/scala/utils/Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_21 & _T_8) begin
          $fwrite(32'h80000002,
            " bpuUpdateReq: valid:%d pc:%x isMissPredict:%d actualTarget:%x actualTaken:%x fuOpType:%x btbType:%x isRVC:%d \n"
            ,_io_redirect_valid_T,io_cfIn_pc,predictWrong,target,taken,io_in_bits_func,_T_78,isRVC); // @[src/main/scala/utils/Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  c = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  c_1 = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  c_2 = _RAND_2[63:0];
  _RAND_3 = {2{`RANDOM}};
  c_3 = _RAND_3[63:0];
  _RAND_4 = {2{`RANDOM}};
  c_4 = _RAND_4[63:0];
  _RAND_5 = {2{`RANDOM}};
  c_5 = _RAND_5[63:0];
  _RAND_6 = {1{`RANDOM}};
  REG_valid = _RAND_6[0:0];
  _RAND_7 = {2{`RANDOM}};
  REG_pc = _RAND_7[38:0];
  _RAND_8 = {1{`RANDOM}};
  REG_isMissPredict = _RAND_8[0:0];
  _RAND_9 = {2{`RANDOM}};
  REG_actualTarget = _RAND_9[38:0];
  _RAND_10 = {1{`RANDOM}};
  REG_actualTaken = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  REG_fuOpType = _RAND_11[6:0];
  _RAND_12 = {1{`RANDOM}};
  REG_btbType = _RAND_12[1:0];
  _RAND_13 = {1{`RANDOM}};
  REG_isRVC = _RAND_13[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module LSExecUnit(
  input         clock,
  input         reset,
  input         io__in_valid, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 290:14]
  input  [63:0] io__in_bits_src1, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 290:14]
  input  [6:0]  io__in_bits_func, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 290:14]
  input         io__out_ready, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 290:14]
  output        io__out_valid, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 290:14]
  output [63:0] io__out_bits, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 290:14]
  input  [63:0] io__wdata, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 290:14]
  input         io__dmem_req_ready, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 290:14]
  output        io__dmem_req_valid, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 290:14]
  output [38:0] io__dmem_req_bits_addr, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 290:14]
  output [2:0]  io__dmem_req_bits_size, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 290:14]
  output [3:0]  io__dmem_req_bits_cmd, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 290:14]
  output [7:0]  io__dmem_req_bits_wmask, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 290:14]
  output [63:0] io__dmem_req_bits_wdata, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 290:14]
  output        io__dmem_resp_ready, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 290:14]
  input         io__dmem_resp_valid, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 290:14]
  input  [63:0] io__dmem_resp_bits_rdata, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 290:14]
  output        io__isMMIO, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 290:14]
  output        io__dtlbPF, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 290:14]
  output        io__loadAddrMisaligned, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 290:14]
  output        io__storeAddrMisaligned, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 290:14]
  output        io_isMMIO,
  input         DISPLAY_ENABLE,
  input         DTLBPF,
  output        r_0,
  output [63:0] io_in_bits_src1,
  input         DTLBENABLE,
  input         ISAMO2,
  input         DTLBFINISH,
  output        r_1_0,
  output        _WIRE_17
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
`endif // RANDOMIZE_REG_INIT
  reg [63:0] addrLatch; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 333:26]
  wire  isStore = io__in_valid & io__in_bits_func[3]; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 334:23]
  wire  _partialLoad_T = ~isStore; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 335:21]
  wire  partialLoad = ~isStore & io__in_bits_func != 7'h3; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 335:30]
  reg [1:0] state; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 338:22]
  wire  _T_1 = io__dmem_req_ready & io__dmem_req_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  wire [1:0] _GEN_2 = DTLBFINISH & DTLBPF ? 2'h0 : state; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 338:22 358:{36,44}]
  wire  _T_11 = io__dmem_resp_ready & io__dmem_resp_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  wire [1:0] _state_T = partialLoad ? 2'h3 : 2'h0; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 361:60]
  wire [1:0] _GEN_4 = _T_11 ? _state_T : state; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 338:22 361:{46,54}]
  wire [1:0] _GEN_5 = 2'h3 == state ? 2'h0 : state; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 351:18 338:22 362:32]
  reg [63:0] c; // @[src/main/scala/utils/GTimer.scala 24:20]
  wire [63:0] _c_T_1 = c + 64'h1; // @[src/main/scala/utils/GTimer.scala 25:12]
  wire  _T_15 = _T_1 & DISPLAY_ENABLE; // @[src/main/scala/utils/Debug.scala 55:16]
  wire  _T_17 = ~reset; // @[src/main/scala/utils/Debug.scala 56:24]
  reg [63:0] c_1; // @[src/main/scala/utils/GTimer.scala 24:20]
  wire [63:0] _c_T_3 = c_1 + 64'h1; // @[src/main/scala/utils/GTimer.scala 25:12]
  wire  _T_28 = DTLBFINISH & DTLBENABLE; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 367:20]
  reg [63:0] c_2; // @[src/main/scala/utils/GTimer.scala 24:20]
  wire [63:0] _c_T_5 = c_2 + 64'h1; // @[src/main/scala/utils/GTimer.scala 25:12]
  wire  _T_31 = _T_28 & DISPLAY_ENABLE; // @[src/main/scala/utils/Debug.scala 55:16]
  wire [63:0] _reqWdata_T_3 = {io__wdata[7:0],io__wdata[7:0],io__wdata[7:0],io__wdata[7:0],io__wdata[7:0],io__wdata[7:0]
    ,io__wdata[7:0],io__wdata[7:0]}; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 310:22]
  wire [63:0] _reqWdata_T_6 = {io__wdata[15:0],io__wdata[15:0],io__wdata[15:0],io__wdata[15:0]}; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 311:22]
  wire [63:0] _reqWdata_T_8 = {io__wdata[31:0],io__wdata[31:0]}; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 312:22]
  wire  _reqWdata_T_9 = 2'h0 == io__in_bits_func[1:0]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _reqWdata_T_10 = 2'h1 == io__in_bits_func[1:0]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _reqWdata_T_11 = 2'h2 == io__in_bits_func[1:0]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _reqWdata_T_12 = 2'h3 == io__in_bits_func[1:0]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _reqWdata_T_13 = _reqWdata_T_9 ? _reqWdata_T_3 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _reqWdata_T_14 = _reqWdata_T_10 ? _reqWdata_T_6 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _reqWdata_T_15 = _reqWdata_T_11 ? _reqWdata_T_8 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _reqWdata_T_16 = _reqWdata_T_12 ? io__wdata : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _reqWdata_T_17 = _reqWdata_T_13 | _reqWdata_T_14; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _reqWdata_T_18 = _reqWdata_T_17 | _reqWdata_T_15; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [1:0] _reqWmask_T_5 = _reqWdata_T_10 ? 2'h3 : 2'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [3:0] _reqWmask_T_6 = _reqWdata_T_11 ? 4'hf : 4'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [7:0] _reqWmask_T_7 = _reqWdata_T_12 ? 8'hff : 8'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [1:0] _GEN_13 = {{1'd0}, _reqWdata_T_9}; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [1:0] _reqWmask_T_8 = _GEN_13 | _reqWmask_T_5; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [3:0] _GEN_14 = {{2'd0}, _reqWmask_T_8}; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [3:0] _reqWmask_T_9 = _GEN_14 | _reqWmask_T_6; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [7:0] _GEN_15 = {{4'd0}, _reqWmask_T_9}; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [7:0] _reqWmask_T_10 = _GEN_15 | _reqWmask_T_7; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [14:0] _GEN_23 = {{7'd0}, _reqWmask_T_10}; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 306:8]
  wire [14:0] reqWmask = _GEN_23 << io__in_bits_src1[2:0]; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 306:8]
  wire  _io_out_valid_T_8 = partialLoad ? state == 2'h3 : _T_11 & state == 2'h2; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 382:114]
  wire  _T_36 = io__out_ready & io__out_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  reg [63:0] c_3; // @[src/main/scala/utils/GTimer.scala 24:20]
  wire [63:0] _c_T_7 = c_3 + 64'h1; // @[src/main/scala/utils/GTimer.scala 25:12]
  wire  _T_38 = _T_36 & DISPLAY_ENABLE; // @[src/main/scala/utils/Debug.scala 55:16]
  reg [63:0] rdataLatch; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 388:27]
  wire  _rdataSel64_T_9 = 3'h0 == addrLatch[2:0]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _rdataSel64_T_10 = 3'h1 == addrLatch[2:0]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _rdataSel64_T_11 = 3'h2 == addrLatch[2:0]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _rdataSel64_T_12 = 3'h3 == addrLatch[2:0]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _rdataSel64_T_13 = 3'h4 == addrLatch[2:0]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _rdataSel64_T_14 = 3'h5 == addrLatch[2:0]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _rdataSel64_T_15 = 3'h6 == addrLatch[2:0]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _rdataSel64_T_16 = 3'h7 == addrLatch[2:0]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdataSel64_T_17 = _rdataSel64_T_9 ? rdataLatch : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [55:0] _rdataSel64_T_18 = _rdataSel64_T_10 ? rdataLatch[63:8] : 56'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [47:0] _rdataSel64_T_19 = _rdataSel64_T_11 ? rdataLatch[63:16] : 48'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [39:0] _rdataSel64_T_20 = _rdataSel64_T_12 ? rdataLatch[63:24] : 40'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] _rdataSel64_T_21 = _rdataSel64_T_13 ? rdataLatch[63:32] : 32'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [23:0] _rdataSel64_T_22 = _rdataSel64_T_14 ? rdataLatch[63:40] : 24'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [15:0] _rdataSel64_T_23 = _rdataSel64_T_15 ? rdataLatch[63:48] : 16'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [7:0] _rdataSel64_T_24 = _rdataSel64_T_16 ? rdataLatch[63:56] : 8'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _GEN_16 = {{8'd0}, _rdataSel64_T_18}; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdataSel64_T_25 = _rdataSel64_T_17 | _GEN_16; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _GEN_17 = {{16'd0}, _rdataSel64_T_19}; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdataSel64_T_26 = _rdataSel64_T_25 | _GEN_17; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _GEN_18 = {{24'd0}, _rdataSel64_T_20}; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdataSel64_T_27 = _rdataSel64_T_26 | _GEN_18; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _GEN_19 = {{32'd0}, _rdataSel64_T_21}; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdataSel64_T_28 = _rdataSel64_T_27 | _GEN_19; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _GEN_20 = {{40'd0}, _rdataSel64_T_22}; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdataSel64_T_29 = _rdataSel64_T_28 | _GEN_20; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _GEN_21 = {{48'd0}, _rdataSel64_T_23}; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdataSel64_T_30 = _rdataSel64_T_29 | _GEN_21; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _GEN_22 = {{56'd0}, _rdataSel64_T_24}; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] rdataSel64 = _rdataSel64_T_30 | _GEN_22; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  rdataPartialLoad_signBit = rdataSel64[7]; // @[src/main/scala/utils/BitUtils.scala 41:20]
  wire [55:0] _rdataPartialLoad_T_2 = rdataPartialLoad_signBit ? 56'hffffffffffffff : 56'h0; // @[src/main/scala/utils/BitUtils.scala 42:46]
  wire [63:0] _rdataPartialLoad_T_3 = {_rdataPartialLoad_T_2,rdataSel64[7:0]}; // @[src/main/scala/utils/BitUtils.scala 42:41]
  wire  rdataPartialLoad_signBit_1 = rdataSel64[15]; // @[src/main/scala/utils/BitUtils.scala 41:20]
  wire [47:0] _rdataPartialLoad_T_6 = rdataPartialLoad_signBit_1 ? 48'hffffffffffff : 48'h0; // @[src/main/scala/utils/BitUtils.scala 42:46]
  wire [63:0] _rdataPartialLoad_T_7 = {_rdataPartialLoad_T_6,rdataSel64[15:0]}; // @[src/main/scala/utils/BitUtils.scala 42:41]
  wire  rdataPartialLoad_signBit_2 = rdataSel64[31]; // @[src/main/scala/utils/BitUtils.scala 41:20]
  wire [31:0] _rdataPartialLoad_T_10 = rdataPartialLoad_signBit_2 ? 32'hffffffff : 32'h0; // @[src/main/scala/utils/BitUtils.scala 42:46]
  wire [63:0] _rdataPartialLoad_T_11 = {_rdataPartialLoad_T_10,rdataSel64[31:0]}; // @[src/main/scala/utils/BitUtils.scala 42:41]
  wire [63:0] _rdataPartialLoad_T_13 = {56'h0,rdataSel64[7:0]}; // @[src/main/scala/utils/BitUtils.scala 49:41]
  wire [63:0] _rdataPartialLoad_T_15 = {48'h0,rdataSel64[15:0]}; // @[src/main/scala/utils/BitUtils.scala 49:41]
  wire [63:0] _rdataPartialLoad_T_17 = {32'h0,rdataSel64[31:0]}; // @[src/main/scala/utils/BitUtils.scala 49:41]
  wire  _rdataPartialLoad_T_18 = 7'h0 == io__in_bits_func; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _rdataPartialLoad_T_19 = 7'h1 == io__in_bits_func; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _rdataPartialLoad_T_20 = 7'h2 == io__in_bits_func; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _rdataPartialLoad_T_21 = 7'h4 == io__in_bits_func; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _rdataPartialLoad_T_22 = 7'h5 == io__in_bits_func; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _rdataPartialLoad_T_23 = 7'h6 == io__in_bits_func; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdataPartialLoad_T_24 = _rdataPartialLoad_T_18 ? _rdataPartialLoad_T_3 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdataPartialLoad_T_25 = _rdataPartialLoad_T_19 ? _rdataPartialLoad_T_7 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdataPartialLoad_T_26 = _rdataPartialLoad_T_20 ? _rdataPartialLoad_T_11 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdataPartialLoad_T_27 = _rdataPartialLoad_T_21 ? _rdataPartialLoad_T_13 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdataPartialLoad_T_28 = _rdataPartialLoad_T_22 ? _rdataPartialLoad_T_15 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdataPartialLoad_T_29 = _rdataPartialLoad_T_23 ? _rdataPartialLoad_T_17 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdataPartialLoad_T_30 = _rdataPartialLoad_T_24 | _rdataPartialLoad_T_25; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdataPartialLoad_T_31 = _rdataPartialLoad_T_30 | _rdataPartialLoad_T_26; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdataPartialLoad_T_32 = _rdataPartialLoad_T_31 | _rdataPartialLoad_T_27; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdataPartialLoad_T_33 = _rdataPartialLoad_T_32 | _rdataPartialLoad_T_28; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] rdataPartialLoad = _rdataPartialLoad_T_33 | _rdataPartialLoad_T_29; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _addrAligned_T_2 = ~io__in_bits_src1[0]; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 416:27]
  wire  _addrAligned_T_4 = io__in_bits_src1[1:0] == 2'h0; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 417:29]
  wire  _addrAligned_T_6 = io__in_bits_src1[2:0] == 3'h0; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 418:29]
  wire  addrAligned = _reqWdata_T_9 | _reqWdata_T_10 & _addrAligned_T_2 | _reqWdata_T_11 & _addrAligned_T_4 |
    _reqWdata_T_12 & _addrAligned_T_6; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _io_loadAddrMisaligned_T_4 = ~addrAligned; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 429:60]
  wire  _T_43 = io__loadAddrMisaligned | io__storeAddrMisaligned; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 432:31]
  reg [63:0] c_4; // @[src/main/scala/utils/GTimer.scala 24:20]
  wire [63:0] _c_T_9 = c_4 + 64'h1; // @[src/main/scala/utils/GTimer.scala 25:12]
  wire  _T_44 = _T_43 & DISPLAY_ENABLE; // @[src/main/scala/utils/Debug.scala 55:16]
  wire  _T_53 = ~io__dmem_req_bits_cmd[0] & ~io__dmem_req_bits_cmd[3]; // @[src/main/scala/bus/simplebus/SimpleBus.scala 73:26]
  wire  _T_54 = io__dmem_req_valid & _T_53; // @[src/main/scala/bus/simplebus/SimpleBus.scala 104:27]
  reg  r; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  _GEN_9 = _T_54 | r; // @[src/main/scala/utils/StopWatch.scala 24:20 30:{20,24}]
  wire  _T_65 = io__dmem_req_valid & io__dmem_req_bits_cmd[0]; // @[src/main/scala/bus/simplebus/SimpleBus.scala 103:27]
  reg  r_1; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  _GEN_11 = _T_65 | r_1; // @[src/main/scala/utils/StopWatch.scala 24:20 30:{20,24}]
  wire  _WIRE = _T_54 & _T_1; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 434:46]
  assign io__out_valid = DTLBPF & state != 2'h0 | io__loadAddrMisaligned | io__storeAddrMisaligned | _io_out_valid_T_8; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 382:22]
  assign io__out_bits = partialLoad ? rdataPartialLoad : io__dmem_resp_bits_rdata; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 421:21]
  assign io__dmem_req_valid = io__in_valid & state == 2'h0 & ~io__loadAddrMisaligned & ~io__storeAddrMisaligned; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 379:75]
  assign io__dmem_req_bits_addr = io__in_bits_src1[38:0]; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 370:68]
  assign io__dmem_req_bits_size = {{1'd0}, io__in_bits_func[1:0]}; // @[src/main/scala/bus/simplebus/SimpleBus.scala 66:15]
  assign io__dmem_req_bits_cmd = {{3'd0}, isStore}; // @[src/main/scala/bus/simplebus/SimpleBus.scala 65:14]
  assign io__dmem_req_bits_wmask = reqWmask[7:0]; // @[src/main/scala/bus/simplebus/SimpleBus.scala 68:16]
  assign io__dmem_req_bits_wdata = _reqWdata_T_18 | _reqWdata_T_16; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign io__dmem_resp_ready = 1'h1; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 380:19]
  assign io__isMMIO = 1'h0;
  assign io__dtlbPF = DTLBPF; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 341:24]
  assign io__loadAddrMisaligned = io__in_valid & _partialLoad_T & ~ISAMO2 & ~addrAligned; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 429:57]
  assign io__storeAddrMisaligned = io__in_valid & (isStore | ISAMO2) & _io_loadAddrMisaligned_T_4; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 430:57]
  assign io_isMMIO = io__isMMIO;
  assign r_0 = r;
  assign io_in_bits_src1 = io__in_bits_src1;
  assign r_1_0 = r_1;
  assign _WIRE_17 = _WIRE;
  always @(posedge clock) begin
    addrLatch <= io__in_bits_src1; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 333:26]
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 338:22]
      state <= 2'h0; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 338:22]
    end else if (2'h0 == state) begin // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 351:18]
      if (_T_1 & ~DTLBENABLE) begin // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 354:43]
        state <= 2'h2; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 354:51]
      end else if (_T_1 & DTLBENABLE) begin // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 353:43]
        state <= 2'h1; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 353:51]
      end
    end else if (2'h1 == state) begin // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 351:18]
      if (DTLBFINISH & ~DTLBPF) begin // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 359:36]
        state <= 2'h2; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 359:44]
      end else begin
        state <= _GEN_2;
      end
    end else if (2'h2 == state) begin // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 351:18]
      state <= _GEN_4;
    end else begin
      state <= _GEN_5;
    end
    if (reset) begin // @[src/main/scala/utils/GTimer.scala 24:20]
      c <= 64'h0; // @[src/main/scala/utils/GTimer.scala 24:20]
    end else begin
      c <= _c_T_1; // @[src/main/scala/utils/GTimer.scala 25:7]
    end
    if (reset) begin // @[src/main/scala/utils/GTimer.scala 24:20]
      c_1 <= 64'h0; // @[src/main/scala/utils/GTimer.scala 24:20]
    end else begin
      c_1 <= _c_T_3; // @[src/main/scala/utils/GTimer.scala 25:7]
    end
    if (reset) begin // @[src/main/scala/utils/GTimer.scala 24:20]
      c_2 <= 64'h0; // @[src/main/scala/utils/GTimer.scala 24:20]
    end else begin
      c_2 <= _c_T_5; // @[src/main/scala/utils/GTimer.scala 25:7]
    end
    if (reset) begin // @[src/main/scala/utils/GTimer.scala 24:20]
      c_3 <= 64'h0; // @[src/main/scala/utils/GTimer.scala 24:20]
    end else begin
      c_3 <= _c_T_7; // @[src/main/scala/utils/GTimer.scala 25:7]
    end
    rdataLatch <= io__dmem_resp_bits_rdata; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 388:27]
    if (reset) begin // @[src/main/scala/utils/GTimer.scala 24:20]
      c_4 <= 64'h0; // @[src/main/scala/utils/GTimer.scala 24:20]
    end else begin
      c_4 <= _c_T_9; // @[src/main/scala/utils/GTimer.scala 25:7]
    end
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      r <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else if (_T_11) begin // @[src/main/scala/utils/StopWatch.scala 31:19]
      r <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 31:23]
    end else begin
      r <= _GEN_9;
    end
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      r_1 <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else if (_T_11) begin // @[src/main/scala/utils/StopWatch.scala 31:19]
      r_1 <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 31:23]
    end else begin
      r_1 <= _GEN_11;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_15 & ~reset) begin
          $fwrite(32'h80000002,"[%d] LSExecUnit: ",c); // @[src/main/scala/utils/Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_15 & _T_17) begin
          $fwrite(32'h80000002,"[LSU] %x, size %x, wdata_raw %x, isStore %x\n",io__in_bits_src1,io__in_bits_func[1:0],
            io__wdata,isStore); // @[src/main/scala/utils/Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_15 & ~reset) begin
          $fwrite(32'h80000002,"[%d] LSExecUnit: ",c_1); // @[src/main/scala/utils/Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_15 & _T_17) begin
          $fwrite(32'h80000002,
            "[LSU] dtlbFinish:%d dtlbEnable:%d dtlbPF:%d state:%d addr:%x dmemReqFire:%d dmemRespFire:%d dmemRdata:%x\n"
            ,DTLBFINISH,DTLBENABLE,DTLBPF,state,io__dmem_req_bits_addr,_T_1,_T_11,io__dmem_resp_bits_rdata); // @[src/main/scala/utils/Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_31 & ~reset) begin
          $fwrite(32'h80000002,"[%d] LSExecUnit: ",c_2); // @[src/main/scala/utils/Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_31 & _T_17) begin
          $fwrite(32'h80000002,
            "[LSU] dtlbFinish:%d dtlbEnable:%d dtlbPF:%d state:%d addr:%x dmemReqFire:%d dmemRespFire:%d dmemRdata:%x\n"
            ,DTLBFINISH,DTLBENABLE,DTLBPF,state,io__dmem_req_bits_addr,_T_1,_T_11,io__dmem_resp_bits_rdata); // @[src/main/scala/utils/Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_38 & ~reset) begin
          $fwrite(32'h80000002,"[%d] LSExecUnit: ",c_3); // @[src/main/scala/utils/Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_38 & _T_17) begin
          $fwrite(32'h80000002,"[LSU-EXECUNIT] state %x dresp %x dpf %x lm %x sm %x\n",state,_T_11,DTLBPF,
            io__loadAddrMisaligned,io__storeAddrMisaligned); // @[src/main/scala/utils/Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_44 & ~reset) begin
          $fwrite(32'h80000002,"[%d] LSExecUnit: ",c_4); // @[src/main/scala/utils/Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_44 & _T_17) begin
          $fwrite(32'h80000002,"misaligned addr detected\n"); // @[src/main/scala/utils/Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  addrLatch = _RAND_0[63:0];
  _RAND_1 = {1{`RANDOM}};
  state = _RAND_1[1:0];
  _RAND_2 = {2{`RANDOM}};
  c = _RAND_2[63:0];
  _RAND_3 = {2{`RANDOM}};
  c_1 = _RAND_3[63:0];
  _RAND_4 = {2{`RANDOM}};
  c_2 = _RAND_4[63:0];
  _RAND_5 = {2{`RANDOM}};
  c_3 = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  rdataLatch = _RAND_6[63:0];
  _RAND_7 = {2{`RANDOM}};
  c_4 = _RAND_7[63:0];
  _RAND_8 = {1{`RANDOM}};
  r = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  r_1 = _RAND_9[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module AtomALU(
  input  [63:0] io_src1, // @[src/main/scala/nutcore/backend/fu/LSU.scala 171:14]
  input  [63:0] io_src2, // @[src/main/scala/nutcore/backend/fu/LSU.scala 171:14]
  input  [6:0]  io_func, // @[src/main/scala/nutcore/backend/fu/LSU.scala 171:14]
  input         io_isWordOp, // @[src/main/scala/nutcore/backend/fu/LSU.scala 171:14]
  output [63:0] io_result // @[src/main/scala/nutcore/backend/fu/LSU.scala 171:14]
);
  wire  isAdderSub = ~io_func[6]; // @[src/main/scala/nutcore/backend/fu/LSU.scala 184:20]
  wire [63:0] _adderRes_T_1 = isAdderSub ? 64'hffffffffffffffff : 64'h0; // @[src/main/scala/nutcore/backend/fu/LSU.scala 185:39]
  wire [63:0] _adderRes_T_2 = io_src2 ^ _adderRes_T_1; // @[src/main/scala/nutcore/backend/fu/LSU.scala 185:33]
  wire [64:0] _adderRes_T_3 = io_src1 + _adderRes_T_2; // @[src/main/scala/nutcore/backend/fu/LSU.scala 185:24]
  wire [64:0] _GEN_0 = {{64'd0}, isAdderSub}; // @[src/main/scala/nutcore/backend/fu/LSU.scala 185:60]
  wire [64:0] adderRes = _adderRes_T_3 + _GEN_0; // @[src/main/scala/nutcore/backend/fu/LSU.scala 185:60]
  wire [63:0] xorRes = io_src1 ^ io_src2; // @[src/main/scala/nutcore/backend/fu/LSU.scala 186:21]
  wire  sltu = ~adderRes[64]; // @[src/main/scala/nutcore/backend/fu/LSU.scala 187:14]
  wire  slt = xorRes[63] ^ sltu; // @[src/main/scala/nutcore/backend/fu/LSU.scala 188:28]
  wire [63:0] _res_T_1 = io_src1 & io_src2; // @[src/main/scala/nutcore/backend/fu/LSU.scala 194:32]
  wire [63:0] _res_T_2 = io_src1 | io_src2; // @[src/main/scala/nutcore/backend/fu/LSU.scala 195:32]
  wire [63:0] _res_T_4 = slt ? io_src1 : io_src2; // @[src/main/scala/nutcore/backend/fu/LSU.scala 196:29]
  wire [63:0] _res_T_6 = slt ? io_src2 : io_src1; // @[src/main/scala/nutcore/backend/fu/LSU.scala 197:29]
  wire [63:0] _res_T_8 = sltu ? io_src1 : io_src2; // @[src/main/scala/nutcore/backend/fu/LSU.scala 198:29]
  wire [63:0] _res_T_10 = sltu ? io_src2 : io_src1; // @[src/main/scala/nutcore/backend/fu/LSU.scala 199:29]
  wire [64:0] _res_T_12 = 6'h22 == io_func[5:0] ? {{1'd0}, io_src2} : adderRes; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [64:0] _res_T_14 = 6'h24 == io_func[5:0] ? {{1'd0}, xorRes} : _res_T_12; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [64:0] _res_T_16 = 6'h25 == io_func[5:0] ? {{1'd0}, _res_T_1} : _res_T_14; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [64:0] _res_T_18 = 6'h26 == io_func[5:0] ? {{1'd0}, _res_T_2} : _res_T_16; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [64:0] _res_T_20 = 6'h37 == io_func[5:0] ? {{1'd0}, _res_T_4} : _res_T_18; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [64:0] _res_T_22 = 6'h30 == io_func[5:0] ? {{1'd0}, _res_T_6} : _res_T_20; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [64:0] _res_T_24 = 6'h31 == io_func[5:0] ? {{1'd0}, _res_T_8} : _res_T_22; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [64:0] res = 6'h32 == io_func[5:0] ? {{1'd0}, _res_T_10} : _res_T_24; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  io_result_signBit = res[31]; // @[src/main/scala/utils/BitUtils.scala 41:20]
  wire [31:0] _io_result_T_2 = io_result_signBit ? 32'hffffffff : 32'h0; // @[src/main/scala/utils/BitUtils.scala 42:46]
  wire [63:0] _io_result_T_3 = {_io_result_T_2,res[31:0]}; // @[src/main/scala/utils/BitUtils.scala 42:41]
  assign io_result = io_isWordOp ? _io_result_T_3 : res[63:0]; // @[src/main/scala/nutcore/backend/fu/LSU.scala 202:20]
endmodule
module UnpipelinedLSU(
  input         clock,
  input         reset,
  output        io__in_ready, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 37:14]
  input         io__in_valid, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 37:14]
  input  [63:0] io__in_bits_src1, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 37:14]
  input  [63:0] io__in_bits_src2, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 37:14]
  input  [6:0]  io__in_bits_func, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 37:14]
  input         io__out_ready, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 37:14]
  output        io__out_valid, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 37:14]
  output [63:0] io__out_bits, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 37:14]
  input  [63:0] io__wdata, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 37:14]
  input  [31:0] io__instr, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 37:14]
  input         io__dmem_req_ready, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 37:14]
  output        io__dmem_req_valid, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 37:14]
  output [38:0] io__dmem_req_bits_addr, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 37:14]
  output [2:0]  io__dmem_req_bits_size, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 37:14]
  output [3:0]  io__dmem_req_bits_cmd, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 37:14]
  output [7:0]  io__dmem_req_bits_wmask, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 37:14]
  output [63:0] io__dmem_req_bits_wdata, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 37:14]
  input         io__dmem_resp_valid, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 37:14]
  input  [63:0] io__dmem_resp_bits_rdata, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 37:14]
  output        io__isMMIO, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 37:14]
  output        io__dtlbPF, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 37:14]
  output        io__loadAddrMisaligned, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 37:14]
  output        io__storeAddrMisaligned, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 37:14]
  output        setLr_0,
  input         lr_0,
  output        _WIRE_4,
  input  [63:0] lr_addr,
  output        io_isMMIO,
  input         DISPLAY_ENABLE,
  input         DTLBPF,
  output        r,
  output        setLrVal_0,
  output [63:0] io_in_bits_src1,
  input         DTLBENABLE,
  input         DTLBFINISH,
  output        r_1,
  input         lsuMMIO_0,
  output        _WIRE_16,
  output [63:0] setLrAddr_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [31:0] _RAND_9;
`endif // RANDOMIZE_REG_INIT
  wire  lsExecUnit_clock; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 47:28]
  wire  lsExecUnit_reset; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 47:28]
  wire  lsExecUnit_io__in_valid; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 47:28]
  wire [63:0] lsExecUnit_io__in_bits_src1; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 47:28]
  wire [6:0] lsExecUnit_io__in_bits_func; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 47:28]
  wire  lsExecUnit_io__out_ready; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 47:28]
  wire  lsExecUnit_io__out_valid; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 47:28]
  wire [63:0] lsExecUnit_io__out_bits; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 47:28]
  wire [63:0] lsExecUnit_io__wdata; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 47:28]
  wire  lsExecUnit_io__dmem_req_ready; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 47:28]
  wire  lsExecUnit_io__dmem_req_valid; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 47:28]
  wire [38:0] lsExecUnit_io__dmem_req_bits_addr; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 47:28]
  wire [2:0] lsExecUnit_io__dmem_req_bits_size; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 47:28]
  wire [3:0] lsExecUnit_io__dmem_req_bits_cmd; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 47:28]
  wire [7:0] lsExecUnit_io__dmem_req_bits_wmask; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 47:28]
  wire [63:0] lsExecUnit_io__dmem_req_bits_wdata; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 47:28]
  wire  lsExecUnit_io__dmem_resp_ready; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 47:28]
  wire  lsExecUnit_io__dmem_resp_valid; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 47:28]
  wire [63:0] lsExecUnit_io__dmem_resp_bits_rdata; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 47:28]
  wire  lsExecUnit_io__isMMIO; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 47:28]
  wire  lsExecUnit_io__dtlbPF; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 47:28]
  wire  lsExecUnit_io__loadAddrMisaligned; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 47:28]
  wire  lsExecUnit_io__storeAddrMisaligned; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 47:28]
  wire  lsExecUnit_io_isMMIO; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 47:28]
  wire  lsExecUnit_DISPLAY_ENABLE; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 47:28]
  wire  lsExecUnit_DTLBPF; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 47:28]
  wire  lsExecUnit_r_0; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 47:28]
  wire [63:0] lsExecUnit_io_in_bits_src1; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 47:28]
  wire  lsExecUnit_DTLBENABLE; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 47:28]
  wire  lsExecUnit_ISAMO2; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 47:28]
  wire  lsExecUnit_DTLBFINISH; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 47:28]
  wire  lsExecUnit_r_1_0; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 47:28]
  wire  lsExecUnit__WIRE_17; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 47:28]
  wire [63:0] atomALU_io_src1; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 98:25]
  wire [63:0] atomALU_io_src2; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 98:25]
  wire [6:0] atomALU_io_func; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 98:25]
  wire  atomALU_io_isWordOp; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 98:25]
  wire [63:0] atomALU_io_result; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 98:25]
  wire  atomReq = io__in_valid & io__in_bits_func[5]; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 53:26]
  wire  _amoReq_T_1 = io__in_bits_func == 7'h20; // @[src/main/scala/nutcore/backend/fu/LSU.scala 57:37]
  wire  _amoReq_T_4 = io__in_bits_func == 7'h21; // @[src/main/scala/nutcore/backend/fu/LSU.scala 58:37]
  wire  _amoReq_T_6 = io__in_bits_func[5] & ~_amoReq_T_1 & ~_amoReq_T_4; // @[src/main/scala/nutcore/backend/fu/LSU.scala 59:61]
  wire  amoReq = io__in_valid & _amoReq_T_6; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 54:26]
  wire  lrReq = io__in_valid & _amoReq_T_1; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 55:25]
  wire  scReq = io__in_valid & _amoReq_T_4; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 56:25]
  wire [2:0] funct3 = io__instr[14:12]; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 64:26]
  wire  scInvalid = (io__in_bits_src1 != lr_addr | ~lr_0) & scReq; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 81:46]
  reg [2:0] state; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 95:24]
  reg [63:0] atomMemReg; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 96:25]
  reg [63:0] atomRegReg; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 97:25]
  wire  _T = 3'h0 == state; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 128:20]
  wire  _lsExecUnit_io_in_valid_T = ~atomReq; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 141:56]
  wire [63:0] _lsExecUnit_io_in_bits_src1_T_1 = io__in_bits_src1 + io__in_bits_src2; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 143:46]
  wire  _io_in_ready_T_1 = lsExecUnit_io__out_ready & lsExecUnit_io__out_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  wire [2:0] _GEN_1 = amoReq ? 3'h5 : 3'h0; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 149:17 152:{21,28}]
  wire [2:0] _GEN_2 = lrReq ? 3'h3 : _GEN_1; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 153:{20,27}]
  wire [2:0] _state_T = scInvalid ? 3'h0 : 3'h4; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 154:33]
  wire  _T_1 = 3'h1 == state; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 128:20]
  wire  _T_10 = ~reset; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 167:15]
  wire [2:0] _GEN_4 = io__out_valid ? 3'h0 : state; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 168:{26,33} 95:24]
  wire  _T_13 = 3'h5 == state; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 128:20]
  wire [1:0] _lsExecUnit_io_in_bits_func_T = funct3[0] ? 2'h3 : 2'h2; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 188:42]
  reg [63:0] c; // @[src/main/scala/utils/GTimer.scala 24:20]
  wire [63:0] _c_T_1 = c + 64'h1; // @[src/main/scala/utils/GTimer.scala 25:12]
  wire [2:0] _GEN_5 = _io_in_ready_T_1 ? 3'h6 : state; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 192:37 193:17 95:24]
  wire  _T_20 = 3'h6 == state; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 128:20]
  reg [63:0] c_1; // @[src/main/scala/utils/GTimer.scala 24:20]
  wire [63:0] _c_T_3 = c_1 + 64'h1; // @[src/main/scala/utils/GTimer.scala 25:12]
  wire  _T_26 = 3'h7 == state; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 128:20]
  wire [3:0] _lsExecUnit_io_in_bits_func_T_1 = funct3[0] ? 4'hb : 4'ha; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 219:42]
  reg [63:0] c_2; // @[src/main/scala/utils/GTimer.scala 24:20]
  wire [63:0] _c_T_5 = c_2 + 64'h1; // @[src/main/scala/utils/GTimer.scala 25:12]
  wire [2:0] _GEN_6 = _io_in_ready_T_1 ? 3'h0 : state; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 223:37 224:17 95:24]
  wire  _T_33 = 3'h3 == state; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 128:20]
  reg [63:0] c_3; // @[src/main/scala/utils/GTimer.scala 24:20]
  wire [63:0] _c_T_7 = c_3 + 64'h1; // @[src/main/scala/utils/GTimer.scala 25:12]
  wire  _T_40 = 3'h4 == state; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 128:20]
  reg [63:0] c_4; // @[src/main/scala/utils/GTimer.scala 24:20]
  wire [63:0] _c_T_9 = c_4 + 64'h1; // @[src/main/scala/utils/GTimer.scala 25:12]
  wire [63:0] _GEN_11 = io__in_bits_src1; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 128:20 245:36]
  wire  _GEN_14 = 3'h4 == state & _io_in_ready_T_1; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 128:20 126:32 249:36]
  wire [2:0] _GEN_16 = 3'h4 == state ? _GEN_6 : state; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 128:20 95:24]
  wire  _GEN_17 = 3'h3 == state | 3'h4 == state; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 128:20 229:36]
  wire [3:0] _GEN_20 = 3'h3 == state ? {{2'd0}, _lsExecUnit_io_in_bits_func_T} : _lsExecUnit_io_in_bits_func_T_1; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 128:20 233:36]
  wire  _GEN_22 = 3'h3 == state ? _io_in_ready_T_1 : _GEN_14; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 128:20 235:36]
  wire [2:0] _GEN_24 = 3'h3 == state ? _GEN_6 : _GEN_16; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 128:20]
  wire  _GEN_25 = 3'h7 == state | _GEN_17; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 128:20 215:36]
  wire [3:0] _GEN_28 = 3'h7 == state ? _lsExecUnit_io_in_bits_func_T_1 : _GEN_20; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 128:20 219:36]
  wire [63:0] _GEN_29 = 3'h7 == state ? atomMemReg : io__wdata; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 128:20 220:36]
  wire  _GEN_30 = 3'h7 == state ? _io_in_ready_T_1 : _GEN_22; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 128:20 221:36]
  wire [2:0] _GEN_32 = 3'h7 == state ? _GEN_6 : _GEN_24; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 128:20]
  wire  _GEN_33 = 3'h6 == state ? 1'h0 : _GEN_25; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 128:20 201:36]
  wire  _GEN_34 = 3'h6 == state ? 1'h0 : 1'h1; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 128:20 202:36]
  wire  _GEN_38 = 3'h6 == state ? 1'h0 : _GEN_30; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 128:20 207:36]
  wire [2:0] _GEN_40 = 3'h6 == state ? 3'h7 : _GEN_32; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 128:20 209:15]
  wire  _GEN_42 = 3'h5 == state | _GEN_33; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 128:20 184:36]
  wire  _GEN_43 = 3'h5 == state | _GEN_34; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 128:20 185:36]
  wire [3:0] _GEN_45 = 3'h5 == state ? {{2'd0}, _lsExecUnit_io_in_bits_func_T} : _GEN_28; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 128:20 188:36]
  wire  _GEN_47 = 3'h5 == state ? 1'h0 : _GEN_38; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 128:20 190:36]
  wire [2:0] _GEN_49 = 3'h5 == state ? _GEN_5 : _GEN_40; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 128:20]
  wire  _GEN_52 = 3'h1 == state | _GEN_42; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 128:20 159:36]
  wire  _GEN_53 = 3'h1 == state | _GEN_43; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 128:20 160:36]
  wire [6:0] _GEN_55 = 3'h1 == state ? io__in_bits_func : {{3'd0}, _GEN_45}; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 128:20 163:36]
  wire [63:0] _GEN_56 = 3'h1 == state ? io__wdata : _GEN_29; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 128:20 164:36]
  wire  _GEN_57 = 3'h1 == state ? _io_in_ready_T_1 : _GEN_47; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 128:20 165:36]
  wire  _GEN_58 = 3'h1 == state ? lsExecUnit_io__out_valid : _GEN_47; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 128:20 166:36]
  wire  _GEN_67 = 3'h0 == state ? _io_in_ready_T_1 | scInvalid : _GEN_57; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 128:20 147:38]
  wire  _GEN_68 = 3'h0 == state ? lsExecUnit_io__out_valid | scInvalid : _GEN_58; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 128:20 148:38]
  reg [63:0] c_5; // @[src/main/scala/utils/GTimer.scala 24:20]
  wire [63:0] _c_T_11 = c_5 + 64'h1; // @[src/main/scala/utils/GTimer.scala 25:12]
  wire  _T_50 = io__out_valid & DISPLAY_ENABLE; // @[src/main/scala/utils/Debug.scala 55:16]
  wire [63:0] _io_out_bits_T_1 = state == 3'h7 ? atomRegReg : lsExecUnit_io__out_bits; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 275:45]
  reg  mmioReg; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 280:26]
  wire  _WIRE_1 = amoReq; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 54:26]
  wire  _WIRE = amoReq; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 54:26]
  wire  setLr = io__out_valid & (lrReq | scReq); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 270:26]
  wire  setLrVal = lrReq; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 55:25]
  wire [63:0] setLrAddr = io__in_bits_src1; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 272:15 72:25]
  wire  _GEN_77 = ~_T; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 167:15]
  wire  _GEN_89 = _GEN_77 & ~_T_1 & _T_13 & _io_in_ready_T_1 & DISPLAY_ENABLE; // @[src/main/scala/utils/Debug.scala 56:24]
  wire  _GEN_102 = _GEN_77 & ~_T_1 & ~_T_13 & _T_20 & DISPLAY_ENABLE; // @[src/main/scala/utils/Debug.scala 56:24]
  wire  _GEN_119 = _GEN_77 & ~_T_1 & ~_T_13 & ~_T_20 & _T_26 & _io_in_ready_T_1 & DISPLAY_ENABLE; // @[src/main/scala/utils/Debug.scala 56:24]
  wire  _GEN_141 = _GEN_77 & ~_T_1 & ~_T_13 & ~_T_20 & ~_T_26 & _T_33 & _io_in_ready_T_1 & DISPLAY_ENABLE; // @[src/main/scala/utils/Debug.scala 56:24]
  wire  _GEN_167 = _GEN_77 & ~_T_1 & ~_T_13 & ~_T_20 & ~_T_26 & ~_T_33 & _T_40 & _io_in_ready_T_1 & DISPLAY_ENABLE; // @[src/main/scala/utils/Debug.scala 56:24]
  LSExecUnit lsExecUnit ( // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 47:28]
    .clock(lsExecUnit_clock),
    .reset(lsExecUnit_reset),
    .io__in_valid(lsExecUnit_io__in_valid),
    .io__in_bits_src1(lsExecUnit_io__in_bits_src1),
    .io__in_bits_func(lsExecUnit_io__in_bits_func),
    .io__out_ready(lsExecUnit_io__out_ready),
    .io__out_valid(lsExecUnit_io__out_valid),
    .io__out_bits(lsExecUnit_io__out_bits),
    .io__wdata(lsExecUnit_io__wdata),
    .io__dmem_req_ready(lsExecUnit_io__dmem_req_ready),
    .io__dmem_req_valid(lsExecUnit_io__dmem_req_valid),
    .io__dmem_req_bits_addr(lsExecUnit_io__dmem_req_bits_addr),
    .io__dmem_req_bits_size(lsExecUnit_io__dmem_req_bits_size),
    .io__dmem_req_bits_cmd(lsExecUnit_io__dmem_req_bits_cmd),
    .io__dmem_req_bits_wmask(lsExecUnit_io__dmem_req_bits_wmask),
    .io__dmem_req_bits_wdata(lsExecUnit_io__dmem_req_bits_wdata),
    .io__dmem_resp_ready(lsExecUnit_io__dmem_resp_ready),
    .io__dmem_resp_valid(lsExecUnit_io__dmem_resp_valid),
    .io__dmem_resp_bits_rdata(lsExecUnit_io__dmem_resp_bits_rdata),
    .io__isMMIO(lsExecUnit_io__isMMIO),
    .io__dtlbPF(lsExecUnit_io__dtlbPF),
    .io__loadAddrMisaligned(lsExecUnit_io__loadAddrMisaligned),
    .io__storeAddrMisaligned(lsExecUnit_io__storeAddrMisaligned),
    .io_isMMIO(lsExecUnit_io_isMMIO),
    .DISPLAY_ENABLE(lsExecUnit_DISPLAY_ENABLE),
    .DTLBPF(lsExecUnit_DTLBPF),
    .r_0(lsExecUnit_r_0),
    .io_in_bits_src1(lsExecUnit_io_in_bits_src1),
    .DTLBENABLE(lsExecUnit_DTLBENABLE),
    .ISAMO2(lsExecUnit_ISAMO2),
    .DTLBFINISH(lsExecUnit_DTLBFINISH),
    .r_1_0(lsExecUnit_r_1_0),
    ._WIRE_17(lsExecUnit__WIRE_17)
  );
  AtomALU atomALU ( // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 98:25]
    .io_src1(atomALU_io_src1),
    .io_src2(atomALU_io_src2),
    .io_func(atomALU_io_func),
    .io_isWordOp(atomALU_io_isWordOp),
    .io_result(atomALU_io_result)
  );
  assign io__in_ready = DTLBPF | io__loadAddrMisaligned | io__storeAddrMisaligned | _GEN_67; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 257:68 260:19]
  assign io__out_valid = DTLBPF | io__loadAddrMisaligned | io__storeAddrMisaligned | _GEN_68; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 257:68 259:20]
  assign io__out_bits = scReq ? {{63'd0}, scInvalid} : _io_out_bits_T_1; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 275:23]
  assign io__dmem_req_valid = lsExecUnit_io__dmem_req_valid; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 274:13]
  assign io__dmem_req_bits_addr = lsExecUnit_io__dmem_req_bits_addr; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 274:13]
  assign io__dmem_req_bits_size = lsExecUnit_io__dmem_req_bits_size; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 274:13]
  assign io__dmem_req_bits_cmd = lsExecUnit_io__dmem_req_bits_cmd; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 274:13]
  assign io__dmem_req_bits_wmask = lsExecUnit_io__dmem_req_bits_wmask; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 274:13]
  assign io__dmem_req_bits_wdata = lsExecUnit_io__dmem_req_bits_wdata; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 274:13]
  assign io__isMMIO = mmioReg & io__out_valid; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 283:26]
  assign io__dtlbPF = lsExecUnit_io__dtlbPF; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 49:15]
  assign io__loadAddrMisaligned = lsExecUnit_io__loadAddrMisaligned; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 285:27]
  assign io__storeAddrMisaligned = lsExecUnit_io__storeAddrMisaligned; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 286:28]
  assign setLr_0 = setLr;
  assign _WIRE_4 = _WIRE_1;
  assign io_isMMIO = lsExecUnit_io_isMMIO;
  assign r = lsExecUnit_r_0;
  assign setLrVal_0 = setLrVal;
  assign io_in_bits_src1 = lsExecUnit_io_in_bits_src1;
  assign r_1 = lsExecUnit_r_1_0;
  assign _WIRE_16 = lsExecUnit__WIRE_17;
  assign setLrAddr_0 = _GEN_11;
  assign lsExecUnit_clock = clock;
  assign lsExecUnit_reset = reset;
  assign lsExecUnit_io__in_valid = 3'h0 == state ? io__in_valid & ~atomReq : _GEN_52; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 128:20 141:38]
  assign lsExecUnit_io__in_bits_src1 = 3'h0 == state ? _lsExecUnit_io_in_bits_src1_T_1 : io__in_bits_src1; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 128:20 143:38]
  assign lsExecUnit_io__in_bits_func = 3'h0 == state ? io__in_bits_func : _GEN_55; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 128:20 145:38]
  assign lsExecUnit_io__out_ready = 3'h0 == state | _GEN_53; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 128:20 142:38]
  assign lsExecUnit_io__wdata = 3'h0 == state ? io__wdata : _GEN_56; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 128:20 146:38]
  assign lsExecUnit_io__dmem_req_ready = io__dmem_req_ready; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 274:13]
  assign lsExecUnit_io__dmem_resp_valid = io__dmem_resp_valid; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 274:13]
  assign lsExecUnit_io__dmem_resp_bits_rdata = io__dmem_resp_bits_rdata; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 274:13]
  assign lsExecUnit_DISPLAY_ENABLE = DISPLAY_ENABLE;
  assign lsExecUnit_DTLBPF = DTLBPF;
  assign lsExecUnit_DTLBENABLE = DTLBENABLE;
  assign lsExecUnit_ISAMO2 = _WIRE_1;
  assign lsExecUnit_DTLBFINISH = DTLBFINISH;
  assign atomALU_io_src1 = atomMemReg; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 99:21]
  assign atomALU_io_src2 = io__wdata; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 100:21]
  assign atomALU_io_func = io__in_bits_func; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 101:21]
  assign atomALU_io_isWordOp = ~funct3[0]; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 66:22]
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 95:24]
      state <= 3'h0; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 95:24]
    end else if (DTLBPF | io__loadAddrMisaligned | io__storeAddrMisaligned) begin // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 257:68]
      state <= 3'h0; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 258:13]
    end else if (3'h0 == state) begin // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 128:20]
      if (scReq) begin // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 154:20]
        state <= _state_T; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 154:27]
      end else begin
        state <= _GEN_2;
      end
    end else if (3'h1 == state) begin // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 128:20]
      state <= _GEN_4;
    end else begin
      state <= _GEN_49;
    end
    if (!(3'h0 == state)) begin // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 128:20]
      if (!(3'h1 == state)) begin // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 128:20]
        if (3'h5 == state) begin // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 128:20]
          atomMemReg <= lsExecUnit_io__out_bits; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 196:20]
        end else if (3'h6 == state) begin // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 128:20]
          atomMemReg <= atomALU_io_result; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 210:20]
        end
      end
    end
    if (!(3'h0 == state)) begin // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 128:20]
      if (!(3'h1 == state)) begin // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 128:20]
        if (3'h5 == state) begin // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 128:20]
          atomRegReg <= lsExecUnit_io__out_bits; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 197:20]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/GTimer.scala 24:20]
      c <= 64'h0; // @[src/main/scala/utils/GTimer.scala 24:20]
    end else begin
      c <= _c_T_1; // @[src/main/scala/utils/GTimer.scala 25:7]
    end
    if (reset) begin // @[src/main/scala/utils/GTimer.scala 24:20]
      c_1 <= 64'h0; // @[src/main/scala/utils/GTimer.scala 24:20]
    end else begin
      c_1 <= _c_T_3; // @[src/main/scala/utils/GTimer.scala 25:7]
    end
    if (reset) begin // @[src/main/scala/utils/GTimer.scala 24:20]
      c_2 <= 64'h0; // @[src/main/scala/utils/GTimer.scala 24:20]
    end else begin
      c_2 <= _c_T_5; // @[src/main/scala/utils/GTimer.scala 25:7]
    end
    if (reset) begin // @[src/main/scala/utils/GTimer.scala 24:20]
      c_3 <= 64'h0; // @[src/main/scala/utils/GTimer.scala 24:20]
    end else begin
      c_3 <= _c_T_7; // @[src/main/scala/utils/GTimer.scala 25:7]
    end
    if (reset) begin // @[src/main/scala/utils/GTimer.scala 24:20]
      c_4 <= 64'h0; // @[src/main/scala/utils/GTimer.scala 24:20]
    end else begin
      c_4 <= _c_T_9; // @[src/main/scala/utils/GTimer.scala 25:7]
    end
    if (reset) begin // @[src/main/scala/utils/GTimer.scala 24:20]
      c_5 <= 64'h0; // @[src/main/scala/utils/GTimer.scala 24:20]
    end else begin
      c_5 <= _c_T_11; // @[src/main/scala/utils/GTimer.scala 25:7]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 280:26]
      mmioReg <= 1'h0; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 280:26]
    end else if (io__out_valid) begin // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 282:25]
      mmioReg <= 1'h0; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 282:35]
    end else if (~mmioReg) begin // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 281:21]
      mmioReg <= lsuMMIO_0; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 281:31]
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~_T & _T_1 & ~reset & ~(_lsExecUnit_io_in_valid_T | ~amoReq | ~lrReq | ~scReq)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at UnpipelinedLSU.scala:167 assert(!atomReq || !amoReq || !lrReq || !scReq)\n"); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 167:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(_lsExecUnit_io_in_valid_T | ~amoReq | ~lrReq | ~scReq) & (~_T & _T_1 & ~reset)) begin
          $fatal; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 167:15]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_77 & ~_T_1 & _T_13 & _io_in_ready_T_1 & DISPLAY_ENABLE & _T_10) begin
          $fwrite(32'h80000002,"[%d] UnpipelinedLSU: ",c); // @[src/main/scala/utils/Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_89 & _T_10) begin
          $fwrite(32'h80000002,"[AMO-L] lsExecUnit.io.out.bits %x addr %x src2 %x\n",lsExecUnit_io__out_bits,
            lsExecUnit_io__in_bits_src1,io__wdata); // @[src/main/scala/utils/Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_77 & ~_T_1 & ~_T_13 & _T_20 & DISPLAY_ENABLE & _T_10) begin
          $fwrite(32'h80000002,"[%d] UnpipelinedLSU: ",c_1); // @[src/main/scala/utils/Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_102 & _T_10) begin
          $fwrite(32'h80000002,"[AMO-A] src1 %x src2 %x res %x\n",atomMemReg,io__wdata,atomALU_io_result); // @[src/main/scala/utils/Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_77 & ~_T_1 & ~_T_13 & ~_T_20 & _T_26 & _io_in_ready_T_1 & DISPLAY_ENABLE & _T_10) begin
          $fwrite(32'h80000002,"[%d] UnpipelinedLSU: ",c_2); // @[src/main/scala/utils/Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_119 & _T_10) begin
          $fwrite(32'h80000002,"[AMO-S] atomRegReg %x addr %x\n",atomRegReg,lsExecUnit_io__in_bits_src1); // @[src/main/scala/utils/Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_77 & ~_T_1 & ~_T_13 & ~_T_20 & ~_T_26 & _T_33 & _io_in_ready_T_1 & DISPLAY_ENABLE & _T_10) begin
          $fwrite(32'h80000002,"[%d] UnpipelinedLSU: ",c_3); // @[src/main/scala/utils/Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_141 & _T_10) begin
          $fwrite(32'h80000002,"[LR]\n"); // @[src/main/scala/utils/Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_77 & ~_T_1 & ~_T_13 & ~_T_20 & ~_T_26 & ~_T_33 & _T_40 & _io_in_ready_T_1 & DISPLAY_ENABLE & _T_10
          ) begin
          $fwrite(32'h80000002,"[%d] UnpipelinedLSU: ",c_4); // @[src/main/scala/utils/Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_167 & _T_10) begin
          $fwrite(32'h80000002,"[SC] \n"); // @[src/main/scala/utils/Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_50 & _T_10) begin
          $fwrite(32'h80000002,"[%d] UnpipelinedLSU: ",c_5); // @[src/main/scala/utils/Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_50 & _T_10) begin
          $fwrite(32'h80000002,"[LSU-AGU] state %x inv %x inr %x\n",state,io__in_valid,io__in_ready); // @[src/main/scala/utils/Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[2:0];
  _RAND_1 = {2{`RANDOM}};
  atomMemReg = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  atomRegReg = _RAND_2[63:0];
  _RAND_3 = {2{`RANDOM}};
  c = _RAND_3[63:0];
  _RAND_4 = {2{`RANDOM}};
  c_1 = _RAND_4[63:0];
  _RAND_5 = {2{`RANDOM}};
  c_2 = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  c_3 = _RAND_6[63:0];
  _RAND_7 = {2{`RANDOM}};
  c_4 = _RAND_7[63:0];
  _RAND_8 = {2{`RANDOM}};
  c_5 = _RAND_8[63:0];
  _RAND_9 = {1{`RANDOM}};
  mmioReg = _RAND_9[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Multiplier(
  input          clock,
  input          reset,
  output         io_in_ready, // @[src/main/scala/nutcore/backend/fu/MDU.scala 53:14]
  input          io_in_valid, // @[src/main/scala/nutcore/backend/fu/MDU.scala 53:14]
  input  [64:0]  io_in_bits_0, // @[src/main/scala/nutcore/backend/fu/MDU.scala 53:14]
  input  [64:0]  io_in_bits_1, // @[src/main/scala/nutcore/backend/fu/MDU.scala 53:14]
  input          io_out_ready, // @[src/main/scala/nutcore/backend/fu/MDU.scala 53:14]
  output         io_out_valid, // @[src/main/scala/nutcore/backend/fu/MDU.scala 53:14]
  output [129:0] io_out_bits // @[src/main/scala/nutcore/backend/fu/MDU.scala 53:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [95:0] _RAND_0;
  reg [95:0] _RAND_1;
  reg [159:0] _RAND_2;
  reg [159:0] _RAND_3;
  reg [159:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
`endif // RANDOMIZE_REG_INIT
  reg [64:0] mulRes_REG; // @[src/main/scala/nutcore/backend/fu/MDU.scala 56:43]
  reg [64:0] mulRes_REG_1; // @[src/main/scala/nutcore/backend/fu/MDU.scala 56:43]
  reg [129:0] io_out_bits_REG; // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:60]
  reg [129:0] io_out_bits_REG_1; // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:52]
  reg [129:0] io_out_bits_REG_2; // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:44]
  reg  io_out_valid_REG; // @[src/main/scala/nutcore/backend/fu/MDU.scala 56:43]
  reg  io_out_valid_REG_1; // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:60]
  reg  io_out_valid_REG_2; // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:52]
  reg  io_out_valid_REG_3; // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:44]
  reg  busy; // @[src/main/scala/nutcore/backend/fu/MDU.scala 62:21]
  wire  _GEN_0 = io_in_valid & ~busy | busy; // @[src/main/scala/nutcore/backend/fu/MDU.scala 62:21 63:{31,38}]
  assign io_in_ready = ~busy; // @[src/main/scala/nutcore/backend/fu/MDU.scala 65:49]
  assign io_out_valid = io_out_valid_REG_3; // @[src/main/scala/nutcore/backend/fu/MDU.scala 60:16]
  assign io_out_bits = io_out_bits_REG_2; // @[src/main/scala/nutcore/backend/fu/MDU.scala 59:37]
  always @(posedge clock) begin
    mulRes_REG <= io_in_bits_0; // @[src/main/scala/nutcore/backend/fu/MDU.scala 56:43]
    mulRes_REG_1 <= io_in_bits_1; // @[src/main/scala/nutcore/backend/fu/MDU.scala 56:43]
    io_out_bits_REG <= $signed(mulRes_REG) * $signed(mulRes_REG_1); // @[src/main/scala/nutcore/backend/fu/MDU.scala 58:49]
    io_out_bits_REG_1 <= io_out_bits_REG; // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:52]
    io_out_bits_REG_2 <= io_out_bits_REG_1; // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:44]
    io_out_valid_REG <= io_in_ready & io_in_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
    io_out_valid_REG_1 <= io_out_valid_REG; // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:60]
    io_out_valid_REG_2 <= io_out_valid_REG_1; // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:52]
    io_out_valid_REG_3 <= io_out_valid_REG_2; // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:44]
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/MDU.scala 62:21]
      busy <= 1'h0; // @[src/main/scala/nutcore/backend/fu/MDU.scala 62:21]
    end else if (io_out_valid) begin // @[src/main/scala/nutcore/backend/fu/MDU.scala 64:23]
      busy <= 1'h0; // @[src/main/scala/nutcore/backend/fu/MDU.scala 64:30]
    end else begin
      busy <= _GEN_0;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {3{`RANDOM}};
  mulRes_REG = _RAND_0[64:0];
  _RAND_1 = {3{`RANDOM}};
  mulRes_REG_1 = _RAND_1[64:0];
  _RAND_2 = {5{`RANDOM}};
  io_out_bits_REG = _RAND_2[129:0];
  _RAND_3 = {5{`RANDOM}};
  io_out_bits_REG_1 = _RAND_3[129:0];
  _RAND_4 = {5{`RANDOM}};
  io_out_bits_REG_2 = _RAND_4[129:0];
  _RAND_5 = {1{`RANDOM}};
  io_out_valid_REG = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  io_out_valid_REG_1 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  io_out_valid_REG_2 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  io_out_valid_REG_3 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  busy = _RAND_9[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Divider(
  input          clock,
  input          reset,
  output         io_in_ready, // @[src/main/scala/nutcore/backend/fu/MDU.scala 69:14]
  input          io_in_valid, // @[src/main/scala/nutcore/backend/fu/MDU.scala 69:14]
  input  [63:0]  io_in_bits_0, // @[src/main/scala/nutcore/backend/fu/MDU.scala 69:14]
  input  [63:0]  io_in_bits_1, // @[src/main/scala/nutcore/backend/fu/MDU.scala 69:14]
  input          io_sign, // @[src/main/scala/nutcore/backend/fu/MDU.scala 69:14]
  output         io_out_valid, // @[src/main/scala/nutcore/backend/fu/MDU.scala 69:14]
  output [127:0] io_out_bits // @[src/main/scala/nutcore/backend/fu/MDU.scala 69:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [159:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [95:0] _RAND_5;
  reg [31:0] _RAND_6;
`endif // RANDOMIZE_REG_INIT
  reg [2:0] state; // @[src/main/scala/nutcore/backend/fu/MDU.scala 77:22]
  wire  _newReq_T_1 = io_in_ready & io_in_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  wire  newReq = state == 3'h0 & _newReq_T_1; // @[src/main/scala/nutcore/backend/fu/MDU.scala 78:35]
  wire  divBy0 = io_in_bits_1 == 64'h0; // @[src/main/scala/nutcore/backend/fu/MDU.scala 81:18]
  reg [128:0] shiftReg; // @[src/main/scala/nutcore/backend/fu/MDU.scala 83:21]
  wire [64:0] hi = shiftReg[128:64]; // @[src/main/scala/nutcore/backend/fu/MDU.scala 84:20]
  wire [63:0] lo = shiftReg[63:0]; // @[src/main/scala/nutcore/backend/fu/MDU.scala 85:20]
  wire  aSign = io_in_bits_0[63] & io_sign; // @[src/main/scala/nutcore/backend/fu/MDU.scala 72:24]
  wire [63:0] _T_1 = 64'h0 - io_in_bits_0; // @[src/main/scala/nutcore/backend/fu/MDU.scala 73:16]
  wire [63:0] aVal = aSign ? _T_1 : io_in_bits_0; // @[src/main/scala/nutcore/backend/fu/MDU.scala 73:12]
  wire  bSign = io_in_bits_1[63] & io_sign; // @[src/main/scala/nutcore/backend/fu/MDU.scala 72:24]
  wire [63:0] _T_3 = 64'h0 - io_in_bits_1; // @[src/main/scala/nutcore/backend/fu/MDU.scala 73:16]
  reg  aSignReg; // @[src/main/scala/nutcore/backend/fu/MDU.scala 89:27]
  reg  qSignReg; // @[src/main/scala/nutcore/backend/fu/MDU.scala 90:27]
  reg [63:0] bReg; // @[src/main/scala/nutcore/backend/fu/MDU.scala 91:23]
  wire [64:0] _aValx2Reg_T = {aVal,1'h0}; // @[src/main/scala/nutcore/backend/fu/MDU.scala 92:32]
  reg [64:0] aValx2Reg; // @[src/main/scala/nutcore/backend/fu/MDU.scala 92:28]
  reg [5:0] cnt_value; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
  wire [31:0] canSkipShift_hi = bReg[63:32]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [31:0] canSkipShift_lo = bReg[31:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  canSkipShift_useHi = |canSkipShift_hi; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [15:0] canSkipShift_hi_1 = canSkipShift_hi[31:16]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [15:0] canSkipShift_lo_1 = canSkipShift_hi[15:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  canSkipShift_useHi_1 = |canSkipShift_hi_1; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [7:0] canSkipShift_hi_2 = canSkipShift_hi_1[15:8]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [7:0] canSkipShift_lo_2 = canSkipShift_hi_1[7:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  canSkipShift_useHi_2 = |canSkipShift_hi_2; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [3:0] canSkipShift_hi_3 = canSkipShift_hi_2[7:4]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [3:0] canSkipShift_lo_3 = canSkipShift_hi_2[3:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  canSkipShift_useHi_3 = |canSkipShift_hi_3; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [1:0] _canSkipShift_T_3 = canSkipShift_hi_3[2] ? 2'h2 : {{1'd0}, canSkipShift_hi_3[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_4 = canSkipShift_hi_3[3] ? 2'h3 : _canSkipShift_T_3; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_8 = canSkipShift_lo_3[2] ? 2'h2 : {{1'd0}, canSkipShift_lo_3[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_9 = canSkipShift_lo_3[3] ? 2'h3 : _canSkipShift_T_8; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_10 = canSkipShift_useHi_3 ? _canSkipShift_T_4 : _canSkipShift_T_9; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [2:0] _canSkipShift_T_11 = {canSkipShift_useHi_3,_canSkipShift_T_10}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [3:0] canSkipShift_hi_4 = canSkipShift_lo_2[7:4]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [3:0] canSkipShift_lo_4 = canSkipShift_lo_2[3:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  canSkipShift_useHi_4 = |canSkipShift_hi_4; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [1:0] _canSkipShift_T_15 = canSkipShift_hi_4[2] ? 2'h2 : {{1'd0}, canSkipShift_hi_4[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_16 = canSkipShift_hi_4[3] ? 2'h3 : _canSkipShift_T_15; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_20 = canSkipShift_lo_4[2] ? 2'h2 : {{1'd0}, canSkipShift_lo_4[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_21 = canSkipShift_lo_4[3] ? 2'h3 : _canSkipShift_T_20; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_22 = canSkipShift_useHi_4 ? _canSkipShift_T_16 : _canSkipShift_T_21; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [2:0] _canSkipShift_T_23 = {canSkipShift_useHi_4,_canSkipShift_T_22}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [2:0] _canSkipShift_T_24 = canSkipShift_useHi_2 ? _canSkipShift_T_11 : _canSkipShift_T_23; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [3:0] _canSkipShift_T_25 = {canSkipShift_useHi_2,_canSkipShift_T_24}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [7:0] canSkipShift_hi_5 = canSkipShift_lo_1[15:8]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [7:0] canSkipShift_lo_5 = canSkipShift_lo_1[7:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  canSkipShift_useHi_5 = |canSkipShift_hi_5; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [3:0] canSkipShift_hi_6 = canSkipShift_hi_5[7:4]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [3:0] canSkipShift_lo_6 = canSkipShift_hi_5[3:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  canSkipShift_useHi_6 = |canSkipShift_hi_6; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [1:0] _canSkipShift_T_29 = canSkipShift_hi_6[2] ? 2'h2 : {{1'd0}, canSkipShift_hi_6[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_30 = canSkipShift_hi_6[3] ? 2'h3 : _canSkipShift_T_29; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_34 = canSkipShift_lo_6[2] ? 2'h2 : {{1'd0}, canSkipShift_lo_6[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_35 = canSkipShift_lo_6[3] ? 2'h3 : _canSkipShift_T_34; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_36 = canSkipShift_useHi_6 ? _canSkipShift_T_30 : _canSkipShift_T_35; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [2:0] _canSkipShift_T_37 = {canSkipShift_useHi_6,_canSkipShift_T_36}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [3:0] canSkipShift_hi_7 = canSkipShift_lo_5[7:4]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [3:0] canSkipShift_lo_7 = canSkipShift_lo_5[3:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  canSkipShift_useHi_7 = |canSkipShift_hi_7; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [1:0] _canSkipShift_T_41 = canSkipShift_hi_7[2] ? 2'h2 : {{1'd0}, canSkipShift_hi_7[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_42 = canSkipShift_hi_7[3] ? 2'h3 : _canSkipShift_T_41; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_46 = canSkipShift_lo_7[2] ? 2'h2 : {{1'd0}, canSkipShift_lo_7[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_47 = canSkipShift_lo_7[3] ? 2'h3 : _canSkipShift_T_46; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_48 = canSkipShift_useHi_7 ? _canSkipShift_T_42 : _canSkipShift_T_47; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [2:0] _canSkipShift_T_49 = {canSkipShift_useHi_7,_canSkipShift_T_48}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [2:0] _canSkipShift_T_50 = canSkipShift_useHi_5 ? _canSkipShift_T_37 : _canSkipShift_T_49; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [3:0] _canSkipShift_T_51 = {canSkipShift_useHi_5,_canSkipShift_T_50}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [3:0] _canSkipShift_T_52 = canSkipShift_useHi_1 ? _canSkipShift_T_25 : _canSkipShift_T_51; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [4:0] _canSkipShift_T_53 = {canSkipShift_useHi_1,_canSkipShift_T_52}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [15:0] canSkipShift_hi_8 = canSkipShift_lo[31:16]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [15:0] canSkipShift_lo_8 = canSkipShift_lo[15:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  canSkipShift_useHi_8 = |canSkipShift_hi_8; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [7:0] canSkipShift_hi_9 = canSkipShift_hi_8[15:8]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [7:0] canSkipShift_lo_9 = canSkipShift_hi_8[7:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  canSkipShift_useHi_9 = |canSkipShift_hi_9; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [3:0] canSkipShift_hi_10 = canSkipShift_hi_9[7:4]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [3:0] canSkipShift_lo_10 = canSkipShift_hi_9[3:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  canSkipShift_useHi_10 = |canSkipShift_hi_10; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [1:0] _canSkipShift_T_57 = canSkipShift_hi_10[2] ? 2'h2 : {{1'd0}, canSkipShift_hi_10[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_58 = canSkipShift_hi_10[3] ? 2'h3 : _canSkipShift_T_57; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_62 = canSkipShift_lo_10[2] ? 2'h2 : {{1'd0}, canSkipShift_lo_10[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_63 = canSkipShift_lo_10[3] ? 2'h3 : _canSkipShift_T_62; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_64 = canSkipShift_useHi_10 ? _canSkipShift_T_58 : _canSkipShift_T_63; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [2:0] _canSkipShift_T_65 = {canSkipShift_useHi_10,_canSkipShift_T_64}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [3:0] canSkipShift_hi_11 = canSkipShift_lo_9[7:4]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [3:0] canSkipShift_lo_11 = canSkipShift_lo_9[3:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  canSkipShift_useHi_11 = |canSkipShift_hi_11; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [1:0] _canSkipShift_T_69 = canSkipShift_hi_11[2] ? 2'h2 : {{1'd0}, canSkipShift_hi_11[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_70 = canSkipShift_hi_11[3] ? 2'h3 : _canSkipShift_T_69; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_74 = canSkipShift_lo_11[2] ? 2'h2 : {{1'd0}, canSkipShift_lo_11[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_75 = canSkipShift_lo_11[3] ? 2'h3 : _canSkipShift_T_74; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_76 = canSkipShift_useHi_11 ? _canSkipShift_T_70 : _canSkipShift_T_75; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [2:0] _canSkipShift_T_77 = {canSkipShift_useHi_11,_canSkipShift_T_76}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [2:0] _canSkipShift_T_78 = canSkipShift_useHi_9 ? _canSkipShift_T_65 : _canSkipShift_T_77; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [3:0] _canSkipShift_T_79 = {canSkipShift_useHi_9,_canSkipShift_T_78}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [7:0] canSkipShift_hi_12 = canSkipShift_lo_8[15:8]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [7:0] canSkipShift_lo_12 = canSkipShift_lo_8[7:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  canSkipShift_useHi_12 = |canSkipShift_hi_12; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [3:0] canSkipShift_hi_13 = canSkipShift_hi_12[7:4]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [3:0] canSkipShift_lo_13 = canSkipShift_hi_12[3:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  canSkipShift_useHi_13 = |canSkipShift_hi_13; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [1:0] _canSkipShift_T_83 = canSkipShift_hi_13[2] ? 2'h2 : {{1'd0}, canSkipShift_hi_13[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_84 = canSkipShift_hi_13[3] ? 2'h3 : _canSkipShift_T_83; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_88 = canSkipShift_lo_13[2] ? 2'h2 : {{1'd0}, canSkipShift_lo_13[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_89 = canSkipShift_lo_13[3] ? 2'h3 : _canSkipShift_T_88; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_90 = canSkipShift_useHi_13 ? _canSkipShift_T_84 : _canSkipShift_T_89; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [2:0] _canSkipShift_T_91 = {canSkipShift_useHi_13,_canSkipShift_T_90}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [3:0] canSkipShift_hi_14 = canSkipShift_lo_12[7:4]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [3:0] canSkipShift_lo_14 = canSkipShift_lo_12[3:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  canSkipShift_useHi_14 = |canSkipShift_hi_14; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [1:0] _canSkipShift_T_95 = canSkipShift_hi_14[2] ? 2'h2 : {{1'd0}, canSkipShift_hi_14[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_96 = canSkipShift_hi_14[3] ? 2'h3 : _canSkipShift_T_95; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_100 = canSkipShift_lo_14[2] ? 2'h2 : {{1'd0}, canSkipShift_lo_14[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_101 = canSkipShift_lo_14[3] ? 2'h3 : _canSkipShift_T_100; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_102 = canSkipShift_useHi_14 ? _canSkipShift_T_96 : _canSkipShift_T_101; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [2:0] _canSkipShift_T_103 = {canSkipShift_useHi_14,_canSkipShift_T_102}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [2:0] _canSkipShift_T_104 = canSkipShift_useHi_12 ? _canSkipShift_T_91 : _canSkipShift_T_103; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [3:0] _canSkipShift_T_105 = {canSkipShift_useHi_12,_canSkipShift_T_104}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [3:0] _canSkipShift_T_106 = canSkipShift_useHi_8 ? _canSkipShift_T_79 : _canSkipShift_T_105; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [4:0] _canSkipShift_T_107 = {canSkipShift_useHi_8,_canSkipShift_T_106}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [4:0] _canSkipShift_T_108 = canSkipShift_useHi ? _canSkipShift_T_53 : _canSkipShift_T_107; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [5:0] _canSkipShift_T_109 = {canSkipShift_useHi,_canSkipShift_T_108}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [6:0] _GEN_18 = {{1'd0}, _canSkipShift_T_109}; // @[src/main/scala/nutcore/backend/fu/MDU.scala 105:31]
  wire [6:0] _canSkipShift_T_110 = 7'h40 | _GEN_18; // @[src/main/scala/nutcore/backend/fu/MDU.scala 105:31]
  wire  canSkipShift_hi_15 = aValx2Reg[64]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [63:0] canSkipShift_lo_15 = aValx2Reg[63:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  canSkipShift_useHi_15 = |canSkipShift_hi_15; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [31:0] canSkipShift_hi_16 = canSkipShift_lo_15[63:32]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [31:0] canSkipShift_lo_16 = canSkipShift_lo_15[31:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  canSkipShift_useHi_16 = |canSkipShift_hi_16; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [15:0] canSkipShift_hi_17 = canSkipShift_hi_16[31:16]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [15:0] canSkipShift_lo_17 = canSkipShift_hi_16[15:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  canSkipShift_useHi_17 = |canSkipShift_hi_17; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [7:0] canSkipShift_hi_18 = canSkipShift_hi_17[15:8]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [7:0] canSkipShift_lo_18 = canSkipShift_hi_17[7:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  canSkipShift_useHi_18 = |canSkipShift_hi_18; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [3:0] canSkipShift_hi_19 = canSkipShift_hi_18[7:4]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [3:0] canSkipShift_lo_19 = canSkipShift_hi_18[3:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  canSkipShift_useHi_19 = |canSkipShift_hi_19; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [1:0] _canSkipShift_T_114 = canSkipShift_hi_19[2] ? 2'h2 : {{1'd0}, canSkipShift_hi_19[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_115 = canSkipShift_hi_19[3] ? 2'h3 : _canSkipShift_T_114; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_119 = canSkipShift_lo_19[2] ? 2'h2 : {{1'd0}, canSkipShift_lo_19[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_120 = canSkipShift_lo_19[3] ? 2'h3 : _canSkipShift_T_119; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_121 = canSkipShift_useHi_19 ? _canSkipShift_T_115 : _canSkipShift_T_120; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [2:0] _canSkipShift_T_122 = {canSkipShift_useHi_19,_canSkipShift_T_121}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [3:0] canSkipShift_hi_20 = canSkipShift_lo_18[7:4]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [3:0] canSkipShift_lo_20 = canSkipShift_lo_18[3:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  canSkipShift_useHi_20 = |canSkipShift_hi_20; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [1:0] _canSkipShift_T_126 = canSkipShift_hi_20[2] ? 2'h2 : {{1'd0}, canSkipShift_hi_20[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_127 = canSkipShift_hi_20[3] ? 2'h3 : _canSkipShift_T_126; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_131 = canSkipShift_lo_20[2] ? 2'h2 : {{1'd0}, canSkipShift_lo_20[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_132 = canSkipShift_lo_20[3] ? 2'h3 : _canSkipShift_T_131; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_133 = canSkipShift_useHi_20 ? _canSkipShift_T_127 : _canSkipShift_T_132; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [2:0] _canSkipShift_T_134 = {canSkipShift_useHi_20,_canSkipShift_T_133}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [2:0] _canSkipShift_T_135 = canSkipShift_useHi_18 ? _canSkipShift_T_122 : _canSkipShift_T_134; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [3:0] _canSkipShift_T_136 = {canSkipShift_useHi_18,_canSkipShift_T_135}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [7:0] canSkipShift_hi_21 = canSkipShift_lo_17[15:8]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [7:0] canSkipShift_lo_21 = canSkipShift_lo_17[7:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  canSkipShift_useHi_21 = |canSkipShift_hi_21; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [3:0] canSkipShift_hi_22 = canSkipShift_hi_21[7:4]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [3:0] canSkipShift_lo_22 = canSkipShift_hi_21[3:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  canSkipShift_useHi_22 = |canSkipShift_hi_22; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [1:0] _canSkipShift_T_140 = canSkipShift_hi_22[2] ? 2'h2 : {{1'd0}, canSkipShift_hi_22[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_141 = canSkipShift_hi_22[3] ? 2'h3 : _canSkipShift_T_140; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_145 = canSkipShift_lo_22[2] ? 2'h2 : {{1'd0}, canSkipShift_lo_22[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_146 = canSkipShift_lo_22[3] ? 2'h3 : _canSkipShift_T_145; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_147 = canSkipShift_useHi_22 ? _canSkipShift_T_141 : _canSkipShift_T_146; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [2:0] _canSkipShift_T_148 = {canSkipShift_useHi_22,_canSkipShift_T_147}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [3:0] canSkipShift_hi_23 = canSkipShift_lo_21[7:4]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [3:0] canSkipShift_lo_23 = canSkipShift_lo_21[3:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  canSkipShift_useHi_23 = |canSkipShift_hi_23; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [1:0] _canSkipShift_T_152 = canSkipShift_hi_23[2] ? 2'h2 : {{1'd0}, canSkipShift_hi_23[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_153 = canSkipShift_hi_23[3] ? 2'h3 : _canSkipShift_T_152; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_157 = canSkipShift_lo_23[2] ? 2'h2 : {{1'd0}, canSkipShift_lo_23[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_158 = canSkipShift_lo_23[3] ? 2'h3 : _canSkipShift_T_157; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_159 = canSkipShift_useHi_23 ? _canSkipShift_T_153 : _canSkipShift_T_158; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [2:0] _canSkipShift_T_160 = {canSkipShift_useHi_23,_canSkipShift_T_159}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [2:0] _canSkipShift_T_161 = canSkipShift_useHi_21 ? _canSkipShift_T_148 : _canSkipShift_T_160; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [3:0] _canSkipShift_T_162 = {canSkipShift_useHi_21,_canSkipShift_T_161}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [3:0] _canSkipShift_T_163 = canSkipShift_useHi_17 ? _canSkipShift_T_136 : _canSkipShift_T_162; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [4:0] _canSkipShift_T_164 = {canSkipShift_useHi_17,_canSkipShift_T_163}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [15:0] canSkipShift_hi_24 = canSkipShift_lo_16[31:16]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [15:0] canSkipShift_lo_24 = canSkipShift_lo_16[15:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  canSkipShift_useHi_24 = |canSkipShift_hi_24; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [7:0] canSkipShift_hi_25 = canSkipShift_hi_24[15:8]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [7:0] canSkipShift_lo_25 = canSkipShift_hi_24[7:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  canSkipShift_useHi_25 = |canSkipShift_hi_25; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [3:0] canSkipShift_hi_26 = canSkipShift_hi_25[7:4]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [3:0] canSkipShift_lo_26 = canSkipShift_hi_25[3:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  canSkipShift_useHi_26 = |canSkipShift_hi_26; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [1:0] _canSkipShift_T_168 = canSkipShift_hi_26[2] ? 2'h2 : {{1'd0}, canSkipShift_hi_26[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_169 = canSkipShift_hi_26[3] ? 2'h3 : _canSkipShift_T_168; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_173 = canSkipShift_lo_26[2] ? 2'h2 : {{1'd0}, canSkipShift_lo_26[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_174 = canSkipShift_lo_26[3] ? 2'h3 : _canSkipShift_T_173; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_175 = canSkipShift_useHi_26 ? _canSkipShift_T_169 : _canSkipShift_T_174; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [2:0] _canSkipShift_T_176 = {canSkipShift_useHi_26,_canSkipShift_T_175}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [3:0] canSkipShift_hi_27 = canSkipShift_lo_25[7:4]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [3:0] canSkipShift_lo_27 = canSkipShift_lo_25[3:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  canSkipShift_useHi_27 = |canSkipShift_hi_27; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [1:0] _canSkipShift_T_180 = canSkipShift_hi_27[2] ? 2'h2 : {{1'd0}, canSkipShift_hi_27[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_181 = canSkipShift_hi_27[3] ? 2'h3 : _canSkipShift_T_180; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_185 = canSkipShift_lo_27[2] ? 2'h2 : {{1'd0}, canSkipShift_lo_27[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_186 = canSkipShift_lo_27[3] ? 2'h3 : _canSkipShift_T_185; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_187 = canSkipShift_useHi_27 ? _canSkipShift_T_181 : _canSkipShift_T_186; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [2:0] _canSkipShift_T_188 = {canSkipShift_useHi_27,_canSkipShift_T_187}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [2:0] _canSkipShift_T_189 = canSkipShift_useHi_25 ? _canSkipShift_T_176 : _canSkipShift_T_188; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [3:0] _canSkipShift_T_190 = {canSkipShift_useHi_25,_canSkipShift_T_189}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [7:0] canSkipShift_hi_28 = canSkipShift_lo_24[15:8]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [7:0] canSkipShift_lo_28 = canSkipShift_lo_24[7:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  canSkipShift_useHi_28 = |canSkipShift_hi_28; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [3:0] canSkipShift_hi_29 = canSkipShift_hi_28[7:4]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [3:0] canSkipShift_lo_29 = canSkipShift_hi_28[3:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  canSkipShift_useHi_29 = |canSkipShift_hi_29; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [1:0] _canSkipShift_T_194 = canSkipShift_hi_29[2] ? 2'h2 : {{1'd0}, canSkipShift_hi_29[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_195 = canSkipShift_hi_29[3] ? 2'h3 : _canSkipShift_T_194; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_199 = canSkipShift_lo_29[2] ? 2'h2 : {{1'd0}, canSkipShift_lo_29[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_200 = canSkipShift_lo_29[3] ? 2'h3 : _canSkipShift_T_199; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_201 = canSkipShift_useHi_29 ? _canSkipShift_T_195 : _canSkipShift_T_200; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [2:0] _canSkipShift_T_202 = {canSkipShift_useHi_29,_canSkipShift_T_201}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [3:0] canSkipShift_hi_30 = canSkipShift_lo_28[7:4]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [3:0] canSkipShift_lo_30 = canSkipShift_lo_28[3:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  canSkipShift_useHi_30 = |canSkipShift_hi_30; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [1:0] _canSkipShift_T_206 = canSkipShift_hi_30[2] ? 2'h2 : {{1'd0}, canSkipShift_hi_30[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_207 = canSkipShift_hi_30[3] ? 2'h3 : _canSkipShift_T_206; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_211 = canSkipShift_lo_30[2] ? 2'h2 : {{1'd0}, canSkipShift_lo_30[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_212 = canSkipShift_lo_30[3] ? 2'h3 : _canSkipShift_T_211; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_213 = canSkipShift_useHi_30 ? _canSkipShift_T_207 : _canSkipShift_T_212; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [2:0] _canSkipShift_T_214 = {canSkipShift_useHi_30,_canSkipShift_T_213}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [2:0] _canSkipShift_T_215 = canSkipShift_useHi_28 ? _canSkipShift_T_202 : _canSkipShift_T_214; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [3:0] _canSkipShift_T_216 = {canSkipShift_useHi_28,_canSkipShift_T_215}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [3:0] _canSkipShift_T_217 = canSkipShift_useHi_24 ? _canSkipShift_T_190 : _canSkipShift_T_216; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [4:0] _canSkipShift_T_218 = {canSkipShift_useHi_24,_canSkipShift_T_217}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [4:0] _canSkipShift_T_219 = canSkipShift_useHi_16 ? _canSkipShift_T_164 : _canSkipShift_T_218; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [5:0] _canSkipShift_T_220 = {canSkipShift_useHi_16,_canSkipShift_T_219}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [5:0] _canSkipShift_T_221 = canSkipShift_useHi_15 ? 6'h0 : _canSkipShift_T_220; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [6:0] _canSkipShift_T_222 = {canSkipShift_useHi_15,_canSkipShift_T_221}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [6:0] canSkipShift = _canSkipShift_T_110 - _canSkipShift_T_222; // @[src/main/scala/nutcore/backend/fu/MDU.scala 105:45]
  wire [6:0] _value_T_1 = canSkipShift >= 7'h3f ? 7'h3f : canSkipShift; // @[src/main/scala/nutcore/backend/fu/MDU.scala 109:38]
  wire [6:0] _value_T_2 = divBy0 ? 7'h0 : _value_T_1; // @[src/main/scala/nutcore/backend/fu/MDU.scala 109:21]
  wire [127:0] _GEN_0 = {{63'd0}, aValx2Reg}; // @[src/main/scala/nutcore/backend/fu/MDU.scala 112:27]
  wire [127:0] _shiftReg_T = _GEN_0 << cnt_value; // @[src/main/scala/nutcore/backend/fu/MDU.scala 112:27]
  wire [64:0] _GEN_19 = {{1'd0}, bReg}; // @[src/main/scala/nutcore/backend/fu/MDU.scala 115:28]
  wire  enough = hi >= _GEN_19; // @[src/main/scala/nutcore/backend/fu/MDU.scala 115:28]
  wire [64:0] _shiftReg_T_2 = hi - _GEN_19; // @[src/main/scala/nutcore/backend/fu/MDU.scala 116:36]
  wire [64:0] _shiftReg_T_3 = enough ? _shiftReg_T_2 : hi; // @[src/main/scala/nutcore/backend/fu/MDU.scala 116:24]
  wire [128:0] _shiftReg_T_5 = {_shiftReg_T_3[63:0],lo,enough}; // @[src/main/scala/nutcore/backend/fu/MDU.scala 116:20]
  wire  wrap = cnt_value == 6'h3f; // @[src/main/scala/chisel3/util/Counter.scala 73:24]
  wire [5:0] _value_T_4 = cnt_value + 6'h1; // @[src/main/scala/chisel3/util/Counter.scala 77:24]
  wire [2:0] _GEN_4 = wrap ? 3'h4 : state; // @[src/main/scala/nutcore/backend/fu/MDU.scala 118:{36,44} 77:22]
  wire [2:0] _GEN_5 = state == 3'h4 ? 3'h0 : state; // @[src/main/scala/nutcore/backend/fu/MDU.scala 119:36 120:11 77:22]
  wire [5:0] _GEN_7 = state == 3'h3 ? _value_T_4 : cnt_value; // @[src/main/scala/nutcore/backend/fu/MDU.scala 114:37 src/main/scala/chisel3/util/Counter.scala 77:15 61:40]
  wire [2:0] _GEN_8 = state == 3'h3 ? _GEN_4 : _GEN_5; // @[src/main/scala/nutcore/backend/fu/MDU.scala 114:37]
  wire [5:0] _GEN_11 = state == 3'h2 ? cnt_value : _GEN_7; // @[src/main/scala/nutcore/backend/fu/MDU.scala 111:35 src/main/scala/chisel3/util/Counter.scala 61:40]
  wire [6:0] _GEN_12 = state == 3'h1 ? _value_T_2 : {{1'd0}, _GEN_11}; // @[src/main/scala/nutcore/backend/fu/MDU.scala 109:15 97:34]
  wire [6:0] _GEN_16 = newReq ? {{1'd0}, cnt_value} : _GEN_12; // @[src/main/scala/nutcore/backend/fu/MDU.scala 95:17 src/main/scala/chisel3/util/Counter.scala 61:40]
  wire [63:0] r = hi[64:1]; // @[src/main/scala/nutcore/backend/fu/MDU.scala 123:13]
  wire [63:0] _resQ_T_1 = 64'h0 - lo; // @[src/main/scala/nutcore/backend/fu/MDU.scala 124:28]
  wire [63:0] resQ = qSignReg ? _resQ_T_1 : lo; // @[src/main/scala/nutcore/backend/fu/MDU.scala 124:17]
  wire [63:0] _resR_T_1 = 64'h0 - r; // @[src/main/scala/nutcore/backend/fu/MDU.scala 125:28]
  wire [63:0] resR = aSignReg ? _resR_T_1 : r; // @[src/main/scala/nutcore/backend/fu/MDU.scala 125:17]
  wire [6:0] _GEN_21 = reset ? 7'h0 : _GEN_16; // @[src/main/scala/chisel3/util/Counter.scala 61:{40,40}]
  assign io_in_ready = state == 3'h0; // @[src/main/scala/nutcore/backend/fu/MDU.scala 129:25]
  assign io_out_valid = state == 3'h4; // @[src/main/scala/nutcore/backend/fu/MDU.scala 128:39]
  assign io_out_bits = {resR,resQ}; // @[src/main/scala/nutcore/backend/fu/MDU.scala 126:21]
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/MDU.scala 77:22]
      state <= 3'h0; // @[src/main/scala/nutcore/backend/fu/MDU.scala 77:22]
    end else if (newReq) begin // @[src/main/scala/nutcore/backend/fu/MDU.scala 95:17]
      state <= 3'h1; // @[src/main/scala/nutcore/backend/fu/MDU.scala 96:11]
    end else if (state == 3'h1) begin // @[src/main/scala/nutcore/backend/fu/MDU.scala 97:34]
      state <= 3'h2; // @[src/main/scala/nutcore/backend/fu/MDU.scala 110:11]
    end else if (state == 3'h2) begin // @[src/main/scala/nutcore/backend/fu/MDU.scala 111:35]
      state <= 3'h3; // @[src/main/scala/nutcore/backend/fu/MDU.scala 113:11]
    end else begin
      state <= _GEN_8;
    end
    if (!(newReq)) begin // @[src/main/scala/nutcore/backend/fu/MDU.scala 95:17]
      if (!(state == 3'h1)) begin // @[src/main/scala/nutcore/backend/fu/MDU.scala 97:34]
        if (state == 3'h2) begin // @[src/main/scala/nutcore/backend/fu/MDU.scala 111:35]
          shiftReg <= {{1'd0}, _shiftReg_T}; // @[src/main/scala/nutcore/backend/fu/MDU.scala 112:14]
        end else if (state == 3'h3) begin // @[src/main/scala/nutcore/backend/fu/MDU.scala 114:37]
          shiftReg <= _shiftReg_T_5; // @[src/main/scala/nutcore/backend/fu/MDU.scala 116:14]
        end
      end
    end
    if (newReq) begin // @[src/main/scala/nutcore/backend/fu/MDU.scala 89:27]
      aSignReg <= aSign; // @[src/main/scala/nutcore/backend/fu/MDU.scala 89:27]
    end
    if (newReq) begin // @[src/main/scala/nutcore/backend/fu/MDU.scala 90:27]
      qSignReg <= (aSign ^ bSign) & ~divBy0; // @[src/main/scala/nutcore/backend/fu/MDU.scala 90:27]
    end
    if (newReq) begin // @[src/main/scala/nutcore/backend/fu/MDU.scala 91:23]
      if (bSign) begin // @[src/main/scala/nutcore/backend/fu/MDU.scala 73:12]
        bReg <= _T_3;
      end else begin
        bReg <= io_in_bits_1;
      end
    end
    if (newReq) begin // @[src/main/scala/nutcore/backend/fu/MDU.scala 92:28]
      aValx2Reg <= _aValx2Reg_T; // @[src/main/scala/nutcore/backend/fu/MDU.scala 92:28]
    end
    cnt_value <= _GEN_21[5:0]; // @[src/main/scala/chisel3/util/Counter.scala 61:{40,40}]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[2:0];
  _RAND_1 = {5{`RANDOM}};
  shiftReg = _RAND_1[128:0];
  _RAND_2 = {1{`RANDOM}};
  aSignReg = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  qSignReg = _RAND_3[0:0];
  _RAND_4 = {2{`RANDOM}};
  bReg = _RAND_4[63:0];
  _RAND_5 = {3{`RANDOM}};
  aValx2Reg = _RAND_5[64:0];
  _RAND_6 = {1{`RANDOM}};
  cnt_value = _RAND_6[5:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module MDU(
  input         clock,
  input         reset,
  output        io_in_ready, // @[src/main/scala/nutcore/backend/fu/MDU.scala 136:14]
  input         io_in_valid, // @[src/main/scala/nutcore/backend/fu/MDU.scala 136:14]
  input  [63:0] io_in_bits_src1, // @[src/main/scala/nutcore/backend/fu/MDU.scala 136:14]
  input  [63:0] io_in_bits_src2, // @[src/main/scala/nutcore/backend/fu/MDU.scala 136:14]
  input  [6:0]  io_in_bits_func, // @[src/main/scala/nutcore/backend/fu/MDU.scala 136:14]
  input         io_out_ready, // @[src/main/scala/nutcore/backend/fu/MDU.scala 136:14]
  output        io_out_valid, // @[src/main/scala/nutcore/backend/fu/MDU.scala 136:14]
  output [63:0] io_out_bits, // @[src/main/scala/nutcore/backend/fu/MDU.scala 136:14]
  output        _WIRE_0,
  input         DISPLAY_ENABLE
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  wire  mul_clock; // @[src/main/scala/nutcore/backend/fu/MDU.scala 151:19]
  wire  mul_reset; // @[src/main/scala/nutcore/backend/fu/MDU.scala 151:19]
  wire  mul_io_in_ready; // @[src/main/scala/nutcore/backend/fu/MDU.scala 151:19]
  wire  mul_io_in_valid; // @[src/main/scala/nutcore/backend/fu/MDU.scala 151:19]
  wire [64:0] mul_io_in_bits_0; // @[src/main/scala/nutcore/backend/fu/MDU.scala 151:19]
  wire [64:0] mul_io_in_bits_1; // @[src/main/scala/nutcore/backend/fu/MDU.scala 151:19]
  wire  mul_io_out_ready; // @[src/main/scala/nutcore/backend/fu/MDU.scala 151:19]
  wire  mul_io_out_valid; // @[src/main/scala/nutcore/backend/fu/MDU.scala 151:19]
  wire [129:0] mul_io_out_bits; // @[src/main/scala/nutcore/backend/fu/MDU.scala 151:19]
  wire  div_clock; // @[src/main/scala/nutcore/backend/fu/MDU.scala 152:19]
  wire  div_reset; // @[src/main/scala/nutcore/backend/fu/MDU.scala 152:19]
  wire  div_io_in_ready; // @[src/main/scala/nutcore/backend/fu/MDU.scala 152:19]
  wire  div_io_in_valid; // @[src/main/scala/nutcore/backend/fu/MDU.scala 152:19]
  wire [63:0] div_io_in_bits_0; // @[src/main/scala/nutcore/backend/fu/MDU.scala 152:19]
  wire [63:0] div_io_in_bits_1; // @[src/main/scala/nutcore/backend/fu/MDU.scala 152:19]
  wire  div_io_sign; // @[src/main/scala/nutcore/backend/fu/MDU.scala 152:19]
  wire  div_io_out_valid; // @[src/main/scala/nutcore/backend/fu/MDU.scala 152:19]
  wire [127:0] div_io_out_bits; // @[src/main/scala/nutcore/backend/fu/MDU.scala 152:19]
  wire  isDiv = io_in_bits_func[2]; // @[src/main/scala/nutcore/backend/fu/MDU.scala 41:27]
  wire  isDivSign = isDiv & ~io_in_bits_func[0]; // @[src/main/scala/nutcore/backend/fu/MDU.scala 42:39]
  wire  isW = io_in_bits_func[3]; // @[src/main/scala/nutcore/backend/fu/MDU.scala 43:25]
  wire [64:0] _mul_io_in_bits_0_T_1 = {1'h0,io_in_bits_src1}; // @[src/main/scala/utils/BitUtils.scala 49:41]
  wire  mul_io_in_bits_0_signBit = io_in_bits_src1[63]; // @[src/main/scala/utils/BitUtils.scala 41:20]
  wire [64:0] _mul_io_in_bits_0_T_2 = {mul_io_in_bits_0_signBit,io_in_bits_src1}; // @[src/main/scala/utils/BitUtils.scala 42:41]
  wire  _mul_io_in_bits_0_T_5 = 2'h0 == io_in_bits_func[1:0]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _mul_io_in_bits_0_T_6 = 2'h1 == io_in_bits_func[1:0]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _mul_io_in_bits_0_T_7 = 2'h2 == io_in_bits_func[1:0]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _mul_io_in_bits_0_T_8 = 2'h3 == io_in_bits_func[1:0]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [64:0] _mul_io_in_bits_0_T_9 = _mul_io_in_bits_0_T_5 ? _mul_io_in_bits_0_T_1 : 65'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [64:0] _mul_io_in_bits_0_T_10 = _mul_io_in_bits_0_T_6 ? _mul_io_in_bits_0_T_2 : 65'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [64:0] _mul_io_in_bits_0_T_11 = _mul_io_in_bits_0_T_7 ? _mul_io_in_bits_0_T_2 : 65'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [64:0] _mul_io_in_bits_0_T_12 = _mul_io_in_bits_0_T_8 ? _mul_io_in_bits_0_T_1 : 65'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [64:0] _mul_io_in_bits_0_T_13 = _mul_io_in_bits_0_T_9 | _mul_io_in_bits_0_T_10; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [64:0] _mul_io_in_bits_0_T_14 = _mul_io_in_bits_0_T_13 | _mul_io_in_bits_0_T_11; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [64:0] _mul_io_in_bits_1_T_1 = {1'h0,io_in_bits_src2}; // @[src/main/scala/utils/BitUtils.scala 49:41]
  wire  mul_io_in_bits_1_signBit = io_in_bits_src2[63]; // @[src/main/scala/utils/BitUtils.scala 41:20]
  wire [64:0] _mul_io_in_bits_1_T_2 = {mul_io_in_bits_1_signBit,io_in_bits_src2}; // @[src/main/scala/utils/BitUtils.scala 42:41]
  wire [64:0] _mul_io_in_bits_1_T_9 = _mul_io_in_bits_0_T_5 ? _mul_io_in_bits_1_T_1 : 65'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [64:0] _mul_io_in_bits_1_T_10 = _mul_io_in_bits_0_T_6 ? _mul_io_in_bits_1_T_2 : 65'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [64:0] _mul_io_in_bits_1_T_11 = _mul_io_in_bits_0_T_7 ? _mul_io_in_bits_1_T_1 : 65'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [64:0] _mul_io_in_bits_1_T_12 = _mul_io_in_bits_0_T_8 ? _mul_io_in_bits_1_T_1 : 65'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [64:0] _mul_io_in_bits_1_T_13 = _mul_io_in_bits_1_T_9 | _mul_io_in_bits_1_T_10; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [64:0] _mul_io_in_bits_1_T_14 = _mul_io_in_bits_1_T_13 | _mul_io_in_bits_1_T_11; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  div_io_in_bits_0_signBit = io_in_bits_src1[31]; // @[src/main/scala/utils/BitUtils.scala 41:20]
  wire [31:0] _div_io_in_bits_0_T_2 = div_io_in_bits_0_signBit ? 32'hffffffff : 32'h0; // @[src/main/scala/utils/BitUtils.scala 42:46]
  wire [63:0] _div_io_in_bits_0_T_3 = {_div_io_in_bits_0_T_2,io_in_bits_src1[31:0]}; // @[src/main/scala/utils/BitUtils.scala 42:41]
  wire [63:0] _div_io_in_bits_0_T_5 = {32'h0,io_in_bits_src1[31:0]}; // @[src/main/scala/utils/BitUtils.scala 49:41]
  wire [63:0] _div_io_in_bits_0_T_6 = isDivSign ? _div_io_in_bits_0_T_3 : _div_io_in_bits_0_T_5; // @[src/main/scala/nutcore/backend/fu/MDU.scala 169:47]
  wire  div_io_in_bits_1_signBit = io_in_bits_src2[31]; // @[src/main/scala/utils/BitUtils.scala 41:20]
  wire [31:0] _div_io_in_bits_1_T_2 = div_io_in_bits_1_signBit ? 32'hffffffff : 32'h0; // @[src/main/scala/utils/BitUtils.scala 42:46]
  wire [63:0] _div_io_in_bits_1_T_3 = {_div_io_in_bits_1_T_2,io_in_bits_src2[31:0]}; // @[src/main/scala/utils/BitUtils.scala 42:41]
  wire [63:0] _div_io_in_bits_1_T_5 = {32'h0,io_in_bits_src2[31:0]}; // @[src/main/scala/utils/BitUtils.scala 49:41]
  wire [63:0] _div_io_in_bits_1_T_6 = isDivSign ? _div_io_in_bits_1_T_3 : _div_io_in_bits_1_T_5; // @[src/main/scala/nutcore/backend/fu/MDU.scala 169:47]
  wire [63:0] mulRes = io_in_bits_func[1:0] == 2'h0 ? mul_io_out_bits[63:0] : mul_io_out_bits[127:64]; // @[src/main/scala/nutcore/backend/fu/MDU.scala 176:19]
  wire [63:0] divRes = io_in_bits_func[1] ? div_io_out_bits[127:64] : div_io_out_bits[63:0]; // @[src/main/scala/nutcore/backend/fu/MDU.scala 177:19]
  wire [63:0] res = isDiv ? divRes : mulRes; // @[src/main/scala/nutcore/backend/fu/MDU.scala 178:16]
  wire  io_out_bits_signBit = res[31]; // @[src/main/scala/utils/BitUtils.scala 41:20]
  wire [31:0] _io_out_bits_T_2 = io_out_bits_signBit ? 32'hffffffff : 32'h0; // @[src/main/scala/utils/BitUtils.scala 42:46]
  wire [63:0] _io_out_bits_T_3 = {_io_out_bits_T_2,res[31:0]}; // @[src/main/scala/utils/BitUtils.scala 42:41]
  wire  _isDivReg_T = io_in_ready & io_in_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  reg  isDivReg_REG; // @[src/main/scala/nutcore/backend/fu/MDU.scala 181:48]
  wire  isDivReg = _isDivReg_T ? isDiv : isDivReg_REG; // @[src/main/scala/nutcore/backend/fu/MDU.scala 181:21]
  reg [63:0] c; // @[src/main/scala/utils/GTimer.scala 24:20]
  wire [63:0] _c_T_1 = c + 64'h1; // @[src/main/scala/utils/GTimer.scala 25:12]
  wire  _T_2 = ~reset; // @[src/main/scala/utils/Debug.scala 56:24]
  wire  _WIRE = mul_io_out_ready & mul_io_out_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  Multiplier mul ( // @[src/main/scala/nutcore/backend/fu/MDU.scala 151:19]
    .clock(mul_clock),
    .reset(mul_reset),
    .io_in_ready(mul_io_in_ready),
    .io_in_valid(mul_io_in_valid),
    .io_in_bits_0(mul_io_in_bits_0),
    .io_in_bits_1(mul_io_in_bits_1),
    .io_out_ready(mul_io_out_ready),
    .io_out_valid(mul_io_out_valid),
    .io_out_bits(mul_io_out_bits)
  );
  Divider div ( // @[src/main/scala/nutcore/backend/fu/MDU.scala 152:19]
    .clock(div_clock),
    .reset(div_reset),
    .io_in_ready(div_io_in_ready),
    .io_in_valid(div_io_in_valid),
    .io_in_bits_0(div_io_in_bits_0),
    .io_in_bits_1(div_io_in_bits_1),
    .io_sign(div_io_sign),
    .io_out_valid(div_io_out_valid),
    .io_out_bits(div_io_out_bits)
  );
  assign io_in_ready = isDiv ? div_io_in_ready : mul_io_in_ready; // @[src/main/scala/nutcore/backend/fu/MDU.scala 182:21]
  assign io_out_valid = isDivReg ? div_io_out_valid : mul_io_out_valid; // @[src/main/scala/nutcore/backend/fu/MDU.scala 183:22]
  assign io_out_bits = isW ? _io_out_bits_T_3 : res; // @[src/main/scala/nutcore/backend/fu/MDU.scala 179:21]
  assign _WIRE_0 = _WIRE;
  assign mul_clock = clock;
  assign mul_reset = reset;
  assign mul_io_in_valid = io_in_valid & ~isDiv; // @[src/main/scala/nutcore/backend/fu/MDU.scala 173:34]
  assign mul_io_in_bits_0 = _mul_io_in_bits_0_T_14 | _mul_io_in_bits_0_T_12; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign mul_io_in_bits_1 = _mul_io_in_bits_1_T_14 | _mul_io_in_bits_1_T_12; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign mul_io_out_ready = 1'h1; // @[src/main/scala/nutcore/backend/fu/MDU.scala 155:17]
  assign div_clock = clock;
  assign div_reset = reset;
  assign div_io_in_valid = io_in_valid & isDiv; // @[src/main/scala/nutcore/backend/fu/MDU.scala 174:34]
  assign div_io_in_bits_0 = isW ? _div_io_in_bits_0_T_6 : io_in_bits_src1; // @[src/main/scala/nutcore/backend/fu/MDU.scala 169:38]
  assign div_io_in_bits_1 = isW ? _div_io_in_bits_1_T_6 : io_in_bits_src2; // @[src/main/scala/nutcore/backend/fu/MDU.scala 169:38]
  assign div_io_sign = isDiv & ~io_in_bits_func[0]; // @[src/main/scala/nutcore/backend/fu/MDU.scala 42:39]
  always @(posedge clock) begin
    isDivReg_REG <= io_in_bits_func[2]; // @[src/main/scala/nutcore/backend/fu/MDU.scala 41:27]
    if (reset) begin // @[src/main/scala/utils/GTimer.scala 24:20]
      c <= 64'h0; // @[src/main/scala/utils/GTimer.scala 24:20]
    end else begin
      c <= _c_T_1; // @[src/main/scala/utils/GTimer.scala 25:7]
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & ~reset) begin
          $fwrite(32'h80000002,"[%d] MDU: ",c); // @[src/main/scala/utils/Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_2) begin
          $fwrite(32'h80000002,"[FU-MDU] irv-orv %d %d - %d %d\n",io_in_ready,io_in_valid,1'h1,io_out_valid); // @[src/main/scala/utils/Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  isDivReg_REG = _RAND_0[0:0];
  _RAND_1 = {2{`RANDOM}};
  c = _RAND_1[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module CSR(
  input         clock,
  input         reset,
  input         io_in_valid, // @[src/main/scala/nutcore/backend/fu/CSR.scala 193:14]
  input  [63:0] io_in_bits_src1, // @[src/main/scala/nutcore/backend/fu/CSR.scala 193:14]
  input  [63:0] io_in_bits_src2, // @[src/main/scala/nutcore/backend/fu/CSR.scala 193:14]
  input  [6:0]  io_in_bits_func, // @[src/main/scala/nutcore/backend/fu/CSR.scala 193:14]
  input         io_out_ready, // @[src/main/scala/nutcore/backend/fu/CSR.scala 193:14]
  output        io_out_valid, // @[src/main/scala/nutcore/backend/fu/CSR.scala 193:14]
  output [63:0] io_out_bits, // @[src/main/scala/nutcore/backend/fu/CSR.scala 193:14]
  input  [63:0] io_cfIn_instr, // @[src/main/scala/nutcore/backend/fu/CSR.scala 193:14]
  input  [38:0] io_cfIn_pc, // @[src/main/scala/nutcore/backend/fu/CSR.scala 193:14]
  input         io_cfIn_exceptionVec_1, // @[src/main/scala/nutcore/backend/fu/CSR.scala 193:14]
  input         io_cfIn_exceptionVec_2, // @[src/main/scala/nutcore/backend/fu/CSR.scala 193:14]
  input         io_cfIn_exceptionVec_4, // @[src/main/scala/nutcore/backend/fu/CSR.scala 193:14]
  input         io_cfIn_exceptionVec_6, // @[src/main/scala/nutcore/backend/fu/CSR.scala 193:14]
  input         io_cfIn_exceptionVec_12, // @[src/main/scala/nutcore/backend/fu/CSR.scala 193:14]
  input         io_cfIn_intrVec_0, // @[src/main/scala/nutcore/backend/fu/CSR.scala 193:14]
  input         io_cfIn_intrVec_1, // @[src/main/scala/nutcore/backend/fu/CSR.scala 193:14]
  input         io_cfIn_intrVec_2, // @[src/main/scala/nutcore/backend/fu/CSR.scala 193:14]
  input         io_cfIn_intrVec_3, // @[src/main/scala/nutcore/backend/fu/CSR.scala 193:14]
  input         io_cfIn_intrVec_4, // @[src/main/scala/nutcore/backend/fu/CSR.scala 193:14]
  input         io_cfIn_intrVec_5, // @[src/main/scala/nutcore/backend/fu/CSR.scala 193:14]
  input         io_cfIn_intrVec_6, // @[src/main/scala/nutcore/backend/fu/CSR.scala 193:14]
  input         io_cfIn_intrVec_7, // @[src/main/scala/nutcore/backend/fu/CSR.scala 193:14]
  input         io_cfIn_intrVec_8, // @[src/main/scala/nutcore/backend/fu/CSR.scala 193:14]
  input         io_cfIn_intrVec_9, // @[src/main/scala/nutcore/backend/fu/CSR.scala 193:14]
  input         io_cfIn_intrVec_10, // @[src/main/scala/nutcore/backend/fu/CSR.scala 193:14]
  input         io_cfIn_intrVec_11, // @[src/main/scala/nutcore/backend/fu/CSR.scala 193:14]
  input         io_cfIn_crossPageIPFFix, // @[src/main/scala/nutcore/backend/fu/CSR.scala 193:14]
  output [38:0] io_redirect_target, // @[src/main/scala/nutcore/backend/fu/CSR.scala 193:14]
  output        io_redirect_valid, // @[src/main/scala/nutcore/backend/fu/CSR.scala 193:14]
  input         io_instrValid, // @[src/main/scala/nutcore/backend/fu/CSR.scala 193:14]
  output [63:0] io_intrNO, // @[src/main/scala/nutcore/backend/fu/CSR.scala 193:14]
  output [1:0]  io_imemMMU_priviledgeMode, // @[src/main/scala/nutcore/backend/fu/CSR.scala 193:14]
  output [1:0]  io_dmemMMU_priviledgeMode, // @[src/main/scala/nutcore/backend/fu/CSR.scala 193:14]
  output        io_dmemMMU_status_sum, // @[src/main/scala/nutcore/backend/fu/CSR.scala 193:14]
  output        io_dmemMMU_status_mxr, // @[src/main/scala/nutcore/backend/fu/CSR.scala 193:14]
  input         io_dmemMMU_loadPF, // @[src/main/scala/nutcore/backend/fu/CSR.scala 193:14]
  input         io_dmemMMU_storePF, // @[src/main/scala/nutcore/backend/fu/CSR.scala 193:14]
  input  [38:0] io_dmemMMU_addr, // @[src/main/scala/nutcore/backend/fu/CSR.scala 193:14]
  output        io_wenFix, // @[src/main/scala/nutcore/backend/fu/CSR.scala 193:14]
  input         set_lr,
  output        lr_0,
  input         MbpBWrong,
  input         perfCntCondMmulInstr,
  input         meip_0,
  input         perfCntCondMlsuInstr,
  output [63:0] lrAddr_0,
  input         perfCntCondMexuBusy,
  input         perfCntCondMmmioInstr,
  input         perfCntCondMaluInstr,
  input         MbpRRight,
  output [63:0] satp_0,
  input         DISPLAY_ENABLE,
  input         MbpIRight,
  input         perfCntCondMcsrInstr,
  input         Custom4,
  input         Custom3,
  input         perfCntCondMifuFlush,
  input         Custom2,
  input         Custom1,
  input         Custom8,
  input         Custom7,
  input         perfCntCondMrawStall,
  input         perfCntCondMloadStall,
  input         Custom6,
  input         Custom5,
  input         perfCntCondISUIssue,
  input         mtip_0,
  input         perfCntCondMultiCommit,
  input         MbpBRight,
  input         perfCntCondMbruInstr,
  input         set_lr_val,
  input         MbpJWrong,
  input         nutcoretrap_0,
  input  [63:0] LSUADDR,
  output [11:0] _WIRE_4,
  input         perfCntCondMstoreStall,
  input         MbpIWrong,
  input         MbpJRight,
  input         perfCntCondMloadInstr,
  input         perfCntCondMmduInstr,
  input  [63:0] set_lr_addr,
  input         perfCntCondMimemStall,
  input         MbpRWrong,
  input         msip_0,
  input         perfCntCondMinstret
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [63:0] _RAND_12;
  reg [63:0] _RAND_13;
  reg [63:0] _RAND_14;
  reg [63:0] _RAND_15;
  reg [63:0] _RAND_16;
  reg [63:0] _RAND_17;
  reg [63:0] _RAND_18;
  reg [63:0] _RAND_19;
  reg [63:0] _RAND_20;
  reg [63:0] _RAND_21;
  reg [63:0] _RAND_22;
  reg [63:0] _RAND_23;
  reg [63:0] _RAND_24;
  reg [63:0] _RAND_25;
  reg [63:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [63:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [63:0] _RAND_30;
  reg [63:0] _RAND_31;
  reg [63:0] _RAND_32;
  reg [63:0] _RAND_33;
  reg [63:0] _RAND_34;
  reg [63:0] _RAND_35;
  reg [63:0] _RAND_36;
  reg [63:0] _RAND_37;
  reg [63:0] _RAND_38;
  reg [63:0] _RAND_39;
  reg [63:0] _RAND_40;
  reg [63:0] _RAND_41;
  reg [63:0] _RAND_42;
  reg [63:0] _RAND_43;
  reg [63:0] _RAND_44;
  reg [63:0] _RAND_45;
  reg [63:0] _RAND_46;
  reg [63:0] _RAND_47;
  reg [63:0] _RAND_48;
  reg [63:0] _RAND_49;
  reg [63:0] _RAND_50;
  reg [63:0] _RAND_51;
  reg [63:0] _RAND_52;
  reg [63:0] _RAND_53;
  reg [63:0] _RAND_54;
  reg [63:0] _RAND_55;
  reg [63:0] _RAND_56;
  reg [63:0] _RAND_57;
  reg [63:0] _RAND_58;
  reg [63:0] _RAND_59;
  reg [63:0] _RAND_60;
  reg [63:0] _RAND_61;
  reg [63:0] _RAND_62;
  reg [63:0] _RAND_63;
  reg [63:0] _RAND_64;
  reg [63:0] _RAND_65;
  reg [63:0] _RAND_66;
  reg [63:0] _RAND_67;
  reg [63:0] _RAND_68;
  reg [63:0] _RAND_69;
  reg [63:0] _RAND_70;
  reg [63:0] _RAND_71;
  reg [63:0] _RAND_72;
  reg [63:0] _RAND_73;
  reg [63:0] _RAND_74;
  reg [63:0] _RAND_75;
  reg [63:0] _RAND_76;
  reg [63:0] _RAND_77;
  reg [63:0] _RAND_78;
  reg [63:0] _RAND_79;
  reg [63:0] _RAND_80;
  reg [63:0] _RAND_81;
  reg [63:0] _RAND_82;
  reg [63:0] _RAND_83;
  reg [63:0] _RAND_84;
  reg [63:0] _RAND_85;
  reg [63:0] _RAND_86;
  reg [63:0] _RAND_87;
  reg [63:0] _RAND_88;
  reg [63:0] _RAND_89;
  reg [63:0] _RAND_90;
  reg [63:0] _RAND_91;
  reg [63:0] _RAND_92;
  reg [63:0] _RAND_93;
  reg [63:0] _RAND_94;
  reg [63:0] _RAND_95;
  reg [63:0] _RAND_96;
  reg [63:0] _RAND_97;
  reg [63:0] _RAND_98;
  reg [63:0] _RAND_99;
  reg [63:0] _RAND_100;
  reg [63:0] _RAND_101;
  reg [63:0] _RAND_102;
  reg [63:0] _RAND_103;
  reg [63:0] _RAND_104;
  reg [63:0] _RAND_105;
  reg [63:0] _RAND_106;
  reg [63:0] _RAND_107;
  reg [63:0] _RAND_108;
  reg [63:0] _RAND_109;
  reg [63:0] _RAND_110;
  reg [63:0] _RAND_111;
  reg [63:0] _RAND_112;
  reg [63:0] _RAND_113;
  reg [63:0] _RAND_114;
  reg [63:0] _RAND_115;
  reg [63:0] _RAND_116;
  reg [63:0] _RAND_117;
  reg [63:0] _RAND_118;
  reg [63:0] _RAND_119;
  reg [63:0] _RAND_120;
  reg [63:0] _RAND_121;
  reg [63:0] _RAND_122;
  reg [63:0] _RAND_123;
  reg [63:0] _RAND_124;
  reg [63:0] _RAND_125;
  reg [63:0] _RAND_126;
  reg [63:0] _RAND_127;
  reg [63:0] _RAND_128;
  reg [63:0] _RAND_129;
  reg [63:0] _RAND_130;
  reg [63:0] _RAND_131;
  reg [63:0] _RAND_132;
  reg [63:0] _RAND_133;
  reg [63:0] _RAND_134;
  reg [63:0] _RAND_135;
  reg [63:0] _RAND_136;
  reg [63:0] _RAND_137;
  reg [63:0] _RAND_138;
  reg [63:0] _RAND_139;
  reg [63:0] _RAND_140;
  reg [63:0] _RAND_141;
  reg [63:0] _RAND_142;
  reg [63:0] _RAND_143;
  reg [63:0] _RAND_144;
  reg [63:0] _RAND_145;
  reg [63:0] _RAND_146;
  reg [63:0] _RAND_147;
  reg [63:0] _RAND_148;
  reg [63:0] _RAND_149;
  reg [63:0] _RAND_150;
  reg [63:0] _RAND_151;
  reg [63:0] _RAND_152;
  reg [63:0] _RAND_153;
  reg [63:0] _RAND_154;
  reg [63:0] _RAND_155;
  reg [63:0] _RAND_156;
  reg [63:0] _RAND_157;
  reg [63:0] _RAND_158;
  reg [63:0] _RAND_159;
  reg [63:0] _RAND_160;
  reg [63:0] _RAND_161;
  reg [63:0] _RAND_162;
  reg [63:0] _RAND_163;
  reg [63:0] _RAND_164;
  reg [63:0] _RAND_165;
  reg [63:0] _RAND_166;
  reg [63:0] _RAND_167;
  reg [63:0] _RAND_168;
  reg [63:0] _RAND_169;
  reg [63:0] _RAND_170;
`endif // RANDOMIZE_REG_INIT
  reg [63:0] mtvec; // @[src/main/scala/nutcore/backend/fu/CSR.scala 252:22]
  reg [63:0] mcounteren; // @[src/main/scala/nutcore/backend/fu/CSR.scala 253:27]
  reg [63:0] mcause; // @[src/main/scala/nutcore/backend/fu/CSR.scala 254:23]
  reg [63:0] mtval; // @[src/main/scala/nutcore/backend/fu/CSR.scala 255:22]
  reg [63:0] mepc; // @[src/main/scala/nutcore/backend/fu/CSR.scala 256:21]
  reg [63:0] mie; // @[src/main/scala/nutcore/backend/fu/CSR.scala 258:20]
  reg [63:0] mipReg; // @[src/main/scala/nutcore/backend/fu/CSR.scala 260:24]
  wire [11:0] _mip_T = {meip_0,1'h0,1'h0,1'h0,mtip_0,1'h0,2'h0,msip_0,3'h0}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 262:22]
  wire [63:0] _GEN_331 = {{52'd0}, _mip_T}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 262:29]
  wire [63:0] _mip_T_1 = _GEN_331 | mipReg; // @[src/main/scala/nutcore/backend/fu/CSR.scala 262:29]
  wire  mip_s_u = _mip_T_1[0]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 262:47]
  wire  mip_s_s = _mip_T_1[1]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 262:47]
  wire  mip_s_h = _mip_T_1[2]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 262:47]
  wire  mip_s_m = _mip_T_1[3]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 262:47]
  wire  mip_t_u = _mip_T_1[4]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 262:47]
  wire  mip_t_s = _mip_T_1[5]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 262:47]
  wire  mip_t_h = _mip_T_1[6]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 262:47]
  wire  mip_t_m = _mip_T_1[7]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 262:47]
  wire  mip_e_u = _mip_T_1[8]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 262:47]
  wire  mip_e_s = _mip_T_1[9]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 262:47]
  wire  mip_e_h = _mip_T_1[10]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 262:47]
  wire  mip_e_m = _mip_T_1[11]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 262:47]
  reg [63:0] misa; // @[src/main/scala/nutcore/backend/fu/CSR.scala 270:21]
  reg [63:0] mstatus; // @[src/main/scala/nutcore/backend/fu/CSR.scala 278:24]
  wire  mstatusStruct_ie_u = mstatus[0]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 299:39]
  wire  mstatusStruct_ie_s = mstatus[1]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 299:39]
  wire  mstatusStruct_ie_h = mstatus[2]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 299:39]
  wire  mstatusStruct_ie_m = mstatus[3]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 299:39]
  wire  mstatusStruct_pie_u = mstatus[4]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 299:39]
  wire  mstatusStruct_pie_s = mstatus[5]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 299:39]
  wire  mstatusStruct_pie_h = mstatus[6]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 299:39]
  wire  mstatusStruct_pie_m = mstatus[7]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 299:39]
  wire  mstatusStruct_spp = mstatus[8]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 299:39]
  wire [1:0] mstatusStruct_hpp = mstatus[10:9]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 299:39]
  wire [1:0] mstatusStruct_mpp = mstatus[12:11]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 299:39]
  wire [1:0] mstatusStruct_fs = mstatus[14:13]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 299:39]
  wire [1:0] mstatusStruct_xs = mstatus[16:15]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 299:39]
  wire  mstatusStruct_mprv = mstatus[17]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 299:39]
  wire  mstatusStruct_sum = mstatus[18]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 299:39]
  wire  mstatusStruct_mxr = mstatus[19]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 299:39]
  wire  mstatusStruct_tvm = mstatus[20]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 299:39]
  wire  mstatusStruct_tw = mstatus[21]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 299:39]
  wire  mstatusStruct_tsr = mstatus[22]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 299:39]
  wire [8:0] mstatusStruct_pad0 = mstatus[31:23]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 299:39]
  wire [1:0] mstatusStruct_uxl = mstatus[33:32]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 299:39]
  wire [1:0] mstatusStruct_sxl = mstatus[35:34]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 299:39]
  wire [26:0] mstatusStruct_pad1 = mstatus[62:36]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 299:39]
  wire  mstatusStruct_sd = mstatus[63]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 299:39]
  reg [63:0] medeleg; // @[src/main/scala/nutcore/backend/fu/CSR.scala 306:24]
  reg [63:0] mideleg; // @[src/main/scala/nutcore/backend/fu/CSR.scala 307:24]
  reg [63:0] mscratch; // @[src/main/scala/nutcore/backend/fu/CSR.scala 308:25]
  reg [63:0] pmpcfg0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 310:24]
  reg [63:0] pmpcfg1; // @[src/main/scala/nutcore/backend/fu/CSR.scala 311:24]
  reg [63:0] pmpcfg2; // @[src/main/scala/nutcore/backend/fu/CSR.scala 312:24]
  reg [63:0] pmpcfg3; // @[src/main/scala/nutcore/backend/fu/CSR.scala 313:24]
  reg [63:0] pmpaddr0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 314:25]
  reg [63:0] pmpaddr1; // @[src/main/scala/nutcore/backend/fu/CSR.scala 315:25]
  reg [63:0] pmpaddr2; // @[src/main/scala/nutcore/backend/fu/CSR.scala 316:25]
  reg [63:0] pmpaddr3; // @[src/main/scala/nutcore/backend/fu/CSR.scala 317:25]
  reg [63:0] stvec; // @[src/main/scala/nutcore/backend/fu/CSR.scala 332:22]
  wire [63:0] sieMask = 64'h222 & mideleg; // @[src/main/scala/nutcore/backend/fu/CSR.scala 334:32]
  reg [63:0] satp; // @[src/main/scala/nutcore/backend/fu/CSR.scala 337:21]
  reg [63:0] sepc; // @[src/main/scala/nutcore/backend/fu/CSR.scala 338:21]
  reg [63:0] scause; // @[src/main/scala/nutcore/backend/fu/CSR.scala 339:23]
  reg [63:0] stval; // @[src/main/scala/nutcore/backend/fu/CSR.scala 340:18]
  reg [63:0] sscratch; // @[src/main/scala/nutcore/backend/fu/CSR.scala 341:25]
  reg [63:0] scounteren; // @[src/main/scala/nutcore/backend/fu/CSR.scala 342:27]
  reg  lr; // @[src/main/scala/nutcore/backend/fu/CSR.scala 355:19]
  reg [63:0] lrAddr; // @[src/main/scala/nutcore/backend/fu/CSR.scala 356:23]
  reg [1:0] priviledgeMode; // @[src/main/scala/nutcore/backend/fu/CSR.scala 369:31]
  reg [63:0] perfCnts_0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
  reg [63:0] perfCnts_1; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
  reg [63:0] perfCnts_2; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
  reg [63:0] perfCnts_3; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
  reg [63:0] perfCnts_4; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
  reg [63:0] perfCnts_5; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
  reg [63:0] perfCnts_6; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
  reg [63:0] perfCnts_7; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
  reg [63:0] perfCnts_8; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
  reg [63:0] perfCnts_9; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
  reg [63:0] perfCnts_10; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
  reg [63:0] perfCnts_11; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
  reg [63:0] perfCnts_12; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
  reg [63:0] perfCnts_13; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
  reg [63:0] perfCnts_14; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
  reg [63:0] perfCnts_15; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
  reg [63:0] perfCnts_16; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
  reg [63:0] perfCnts_17; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
  reg [63:0] perfCnts_18; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
  reg [63:0] perfCnts_19; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
  reg [63:0] perfCnts_20; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
  reg [63:0] perfCnts_21; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
  reg [63:0] perfCnts_22; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
  reg [63:0] perfCnts_23; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
  reg [63:0] perfCnts_24; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
  reg [63:0] perfCnts_25; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
  reg [63:0] perfCnts_26; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
  reg [63:0] perfCnts_27; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
  reg [63:0] perfCnts_28; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
  reg [63:0] perfCnts_29; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
  reg [63:0] perfCnts_30; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
  reg [63:0] perfCnts_31; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
  reg [63:0] perfCnts_32; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
  reg [63:0] perfCnts_33; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
  reg [63:0] perfCnts_34; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
  reg [63:0] perfCnts_35; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
  reg [63:0] perfCnts_36; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
  reg [63:0] perfCnts_37; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
  reg [63:0] perfCnts_38; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
  reg [63:0] perfCnts_39; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
  reg [63:0] perfCnts_40; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
  reg [63:0] perfCnts_41; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
  reg [63:0] perfCnts_42; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
  reg [63:0] perfCnts_43; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
  reg [63:0] perfCnts_44; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
  reg [63:0] perfCnts_45; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
  reg [63:0] perfCnts_46; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
  reg [63:0] perfCnts_47; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
  reg [63:0] perfCnts_48; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
  reg [63:0] perfCnts_49; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
  reg [63:0] perfCnts_50; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
  reg [63:0] perfCnts_51; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
  reg [63:0] perfCnts_52; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
  reg [63:0] perfCnts_53; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
  reg [63:0] perfCnts_54; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
  reg [63:0] perfCnts_55; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
  reg [63:0] perfCnts_56; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
  reg [63:0] perfCnts_57; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
  reg [63:0] perfCnts_58; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
  reg [63:0] perfCnts_59; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
  reg [63:0] perfCnts_60; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
  reg [63:0] perfCnts_61; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
  reg [63:0] perfCnts_62; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
  reg [63:0] perfCnts_63; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
  reg [63:0] perfCnts_64; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
  reg [63:0] perfCnts_65; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
  reg [63:0] perfCnts_66; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
  reg [63:0] perfCnts_67; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
  reg [63:0] perfCnts_68; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
  reg [63:0] perfCnts_69; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
  reg [63:0] perfCnts_70; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
  reg [63:0] perfCnts_71; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
  reg [63:0] perfCnts_72; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
  reg [63:0] perfCnts_73; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
  reg [63:0] perfCnts_74; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
  reg [63:0] perfCnts_75; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
  reg [63:0] perfCnts_76; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
  reg [63:0] perfCnts_77; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
  reg [63:0] perfCnts_78; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
  reg [63:0] perfCnts_79; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
  reg [63:0] perfCnts_80; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
  reg [63:0] perfCnts_81; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
  reg [63:0] perfCnts_82; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
  reg [63:0] perfCnts_83; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
  reg [63:0] perfCnts_84; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
  reg [63:0] perfCnts_85; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
  reg [63:0] perfCnts_86; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
  reg [63:0] perfCnts_87; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
  reg [63:0] perfCnts_88; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
  reg [63:0] perfCnts_89; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
  reg [63:0] perfCnts_90; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
  reg [63:0] perfCnts_91; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
  reg [63:0] perfCnts_92; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
  reg [63:0] perfCnts_93; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
  reg [63:0] perfCnts_94; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
  reg [63:0] perfCnts_95; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
  reg [63:0] perfCnts_96; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
  reg [63:0] perfCnts_97; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
  reg [63:0] perfCnts_98; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
  reg [63:0] perfCnts_99; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
  reg [63:0] perfCnts_100; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
  reg [63:0] perfCnts_101; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
  reg [63:0] perfCnts_102; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
  reg [63:0] perfCnts_103; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
  reg [63:0] perfCnts_104; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
  reg [63:0] perfCnts_105; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
  reg [63:0] perfCnts_106; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
  reg [63:0] perfCnts_107; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
  reg [63:0] perfCnts_108; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
  reg [63:0] perfCnts_109; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
  reg [63:0] perfCnts_110; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
  reg [63:0] perfCnts_111; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
  reg [63:0] perfCnts_112; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
  reg [63:0] perfCnts_113; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
  reg [63:0] perfCnts_114; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
  reg [63:0] perfCnts_115; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
  reg [63:0] perfCnts_116; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
  reg [63:0] perfCnts_117; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
  reg [63:0] perfCnts_118; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
  reg [63:0] perfCnts_119; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
  reg [63:0] perfCnts_120; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
  reg [63:0] perfCnts_121; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
  reg [63:0] perfCnts_122; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
  reg [63:0] perfCnts_123; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
  reg [63:0] perfCnts_124; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
  reg [63:0] perfCnts_125; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
  reg [63:0] perfCnts_126; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
  reg [63:0] perfCnts_127; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
  wire [5:0] lo = {mip_t_s,mip_t_u,mip_s_m,mip_s_h,mip_s_s,mip_s_u}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 417:27]
  wire [11:0] _T_652 = {mip_e_m,mip_e_h,mip_e_s,mip_e_u,mip_t_m,mip_t_h,lo}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 417:27]
  wire [11:0] addr = io_in_bits_src2[11:0]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 457:18]
  wire [63:0] csri = {59'h0,io_cfIn_instr[19:15]}; // @[src/main/scala/utils/BitUtils.scala 49:41]
  wire  _rdata_T_162 = 12'hb06 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_324 = _rdata_T_162 ? perfCnts_6 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_163 = 12'hb49 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_325 = _rdata_T_163 ? perfCnts_73 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_486 = _rdata_T_324 | _rdata_T_325; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_164 = 12'hb3c == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_326 = _rdata_T_164 ? perfCnts_60 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_487 = _rdata_T_486 | _rdata_T_326; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_165 = 12'hb69 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_327 = _rdata_T_165 ? perfCnts_105 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_488 = _rdata_T_487 | _rdata_T_327; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_166 = 12'hb7c == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_328 = _rdata_T_166 ? perfCnts_124 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_489 = _rdata_T_488 | _rdata_T_328; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_167 = 12'hf12 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _rdata_T_168 = 12'hb5c == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_330 = _rdata_T_168 ? perfCnts_92 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_491 = _rdata_T_489 | _rdata_T_330; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_169 = 12'hb15 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_331 = _rdata_T_169 ? perfCnts_21 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_492 = _rdata_T_491 | _rdata_T_331; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_170 = 12'hb26 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_332 = _rdata_T_170 ? perfCnts_38 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_493 = _rdata_T_492 | _rdata_T_332; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_171 = 12'h180 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_333 = _rdata_T_171 ? satp : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_494 = _rdata_T_493 | _rdata_T_333; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_172 = 12'hb66 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_334 = _rdata_T_172 ? perfCnts_102 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_495 = _rdata_T_494 | _rdata_T_334; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_173 = 12'hb75 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_335 = _rdata_T_173 ? perfCnts_117 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_496 = _rdata_T_495 | _rdata_T_335; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_174 = 12'hb1c == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_336 = _rdata_T_174 ? perfCnts_28 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_497 = _rdata_T_496 | _rdata_T_336; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_175 = 12'h3a2 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_337 = _rdata_T_175 ? pmpcfg2 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_498 = _rdata_T_497 | _rdata_T_337; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_176 = 12'hb55 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_338 = _rdata_T_176 ? perfCnts_85 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_499 = _rdata_T_498 | _rdata_T_338; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_177 = 12'h3b1 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_339 = _rdata_T_177 ? pmpaddr1 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_500 = _rdata_T_499 | _rdata_T_339; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_178 = 12'hb46 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_340 = _rdata_T_178 ? perfCnts_70 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_501 = _rdata_T_500 | _rdata_T_340; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_179 = 12'h140 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_341 = _rdata_T_179 ? sscratch : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_502 = _rdata_T_501 | _rdata_T_341; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_180 = 12'hb09 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_342 = _rdata_T_180 ? perfCnts_9 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_503 = _rdata_T_502 | _rdata_T_342; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_181 = 12'hb03 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_343 = _rdata_T_181 ? perfCnts_3 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_504 = _rdata_T_503 | _rdata_T_343; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_182 = 12'hb35 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_344 = _rdata_T_182 ? perfCnts_53 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_505 = _rdata_T_504 | _rdata_T_344; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_183 = 12'hb64 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_345 = _rdata_T_183 ? perfCnts_100 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_506 = _rdata_T_505 | _rdata_T_345; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_184 = 12'hb51 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_346 = _rdata_T_184 ? perfCnts_81 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_507 = _rdata_T_506 | _rdata_T_346; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_185 = 12'hb29 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_347 = _rdata_T_185 ? perfCnts_41 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_508 = _rdata_T_507 | _rdata_T_347; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_186 = 12'h302 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_348 = _rdata_T_186 ? medeleg : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_509 = _rdata_T_508 | _rdata_T_348; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_187 = 12'hb71 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_349 = _rdata_T_187 ? perfCnts_113 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_510 = _rdata_T_509 | _rdata_T_349; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_188 = 12'hb24 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_350 = _rdata_T_188 ? perfCnts_36 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_511 = _rdata_T_510 | _rdata_T_350; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_189 = 12'h105 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_351 = _rdata_T_189 ? stvec : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_512 = _rdata_T_511 | _rdata_T_351; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_190 = 12'hb0d == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_352 = _rdata_T_190 ? perfCnts_13 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_513 = _rdata_T_512 | _rdata_T_352; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_191 = 12'hb6d == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_353 = _rdata_T_191 ? perfCnts_109 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_514 = _rdata_T_513 | _rdata_T_353; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_192 = 12'hb4d == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_354 = _rdata_T_192 ? perfCnts_77 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_515 = _rdata_T_514 | _rdata_T_354; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_193 = 12'h141 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_355 = _rdata_T_193 ? sepc : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_516 = _rdata_T_515 | _rdata_T_355; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_194 = 12'hb40 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_356 = _rdata_T_194 ? perfCnts_64 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_517 = _rdata_T_516 | _rdata_T_356; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_195 = 12'h342 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_357 = _rdata_T_195 ? mcause : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_518 = _rdata_T_517 | _rdata_T_357; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_196 = 12'hb11 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_358 = _rdata_T_196 ? perfCnts_17 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_519 = _rdata_T_518 | _rdata_T_358; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_197 = 12'hb2d == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_359 = _rdata_T_197 ? perfCnts_45 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_520 = _rdata_T_519 | _rdata_T_359; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_198 = 12'h306 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_360 = _rdata_T_198 ? mcounteren : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_521 = _rdata_T_520 | _rdata_T_360; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_199 = 12'hb44 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_361 = _rdata_T_199 ? perfCnts_68 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_522 = _rdata_T_521 | _rdata_T_361; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_200 = 12'hb6a == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_362 = _rdata_T_200 ? perfCnts_106 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_523 = _rdata_T_522 | _rdata_T_362; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_201 = 12'hf11 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _rdata_T_202 = 12'hb5e == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_364 = _rdata_T_202 ? perfCnts_94 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_525 = _rdata_T_523 | _rdata_T_364; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_203 = 12'hb59 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_365 = _rdata_T_203 ? perfCnts_89 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_526 = _rdata_T_525 | _rdata_T_365; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_204 = 12'h104 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_42 = mie & sieMask; // @[src/main/scala/utils/RegMap.scala 48:84]
  wire [63:0] _rdata_T_366 = _rdata_T_204 ? _rdata_T_42 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_527 = _rdata_T_526 | _rdata_T_366; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_205 = 12'hb79 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_367 = _rdata_T_205 ? perfCnts_121 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_528 = _rdata_T_527 | _rdata_T_367; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_206 = 12'hb4a == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_368 = _rdata_T_206 ? perfCnts_74 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_529 = _rdata_T_528 | _rdata_T_368; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_207 = 12'hb39 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_369 = _rdata_T_207 ? perfCnts_57 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_530 = _rdata_T_529 | _rdata_T_369; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_208 = 12'hb38 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_370 = _rdata_T_208 ? perfCnts_56 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_531 = _rdata_T_530 | _rdata_T_370; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_209 = 12'h144 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _GEN_332 = {{52'd0}, _T_652}; // @[src/main/scala/utils/RegMap.scala 48:84]
  wire [63:0] _rdata_T_47 = _GEN_332 & sieMask; // @[src/main/scala/utils/RegMap.scala 48:84]
  wire [63:0] _rdata_T_371 = _rdata_T_209 ? _rdata_T_47 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_532 = _rdata_T_531 | _rdata_T_371; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_210 = 12'hb0a == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_372 = _rdata_T_210 ? perfCnts_10 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_533 = _rdata_T_532 | _rdata_T_372; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_211 = 12'hb04 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_373 = _rdata_T_211 ? perfCnts_4 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_534 = _rdata_T_533 | _rdata_T_373; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_212 = 12'hb18 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_374 = _rdata_T_212 ? perfCnts_24 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_535 = _rdata_T_534 | _rdata_T_374; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_213 = 12'hb4f == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_375 = _rdata_T_213 ? perfCnts_79 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_536 = _rdata_T_535 | _rdata_T_375; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_214 = 12'hb19 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_376 = _rdata_T_214 ? perfCnts_25 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_537 = _rdata_T_536 | _rdata_T_376; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_215 = 12'hb2a == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_377 = _rdata_T_215 ? perfCnts_42 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_538 = _rdata_T_537 | _rdata_T_377; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_216 = 12'h100 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_54 = mstatus & 64'h80000003000de122; // @[src/main/scala/utils/RegMap.scala 48:84]
  wire [63:0] _rdata_T_378 = _rdata_T_216 ? _rdata_T_54 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_539 = _rdata_T_538 | _rdata_T_378; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_217 = 12'hb3d == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_379 = _rdata_T_217 ? perfCnts_61 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_540 = _rdata_T_539 | _rdata_T_379; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_218 = 12'hb0e == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_380 = _rdata_T_218 ? perfCnts_14 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_541 = _rdata_T_540 | _rdata_T_380; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_219 = 12'hb34 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_381 = _rdata_T_219 ? perfCnts_52 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_542 = _rdata_T_541 | _rdata_T_381; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_220 = 12'hb74 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_382 = _rdata_T_220 ? perfCnts_116 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_543 = _rdata_T_542 | _rdata_T_382; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_221 = 12'hb14 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_383 = _rdata_T_221 ? perfCnts_20 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_544 = _rdata_T_543 | _rdata_T_383; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_222 = 12'hb1d == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_384 = _rdata_T_222 ? perfCnts_29 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_545 = _rdata_T_544 | _rdata_T_384; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_223 = 12'hb54 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_385 = _rdata_T_223 ? perfCnts_84 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_546 = _rdata_T_545 | _rdata_T_385; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_224 = 12'hb23 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_386 = _rdata_T_224 ? perfCnts_35 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_547 = _rdata_T_546 | _rdata_T_386; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_225 = 12'hb2e == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_387 = _rdata_T_225 ? perfCnts_46 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_548 = _rdata_T_547 | _rdata_T_387; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_226 = 12'hb6e == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_388 = _rdata_T_226 ? perfCnts_110 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_549 = _rdata_T_548 | _rdata_T_388; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_227 = 12'hb43 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_389 = _rdata_T_227 ? perfCnts_67 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_550 = _rdata_T_549 | _rdata_T_389; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_228 = 12'hb63 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_390 = _rdata_T_228 ? perfCnts_99 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_551 = _rdata_T_550 | _rdata_T_390; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_229 = 12'h305 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_391 = _rdata_T_229 ? mtvec : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_552 = _rdata_T_551 | _rdata_T_391; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_230 = 12'hb5d == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_392 = _rdata_T_230 ? perfCnts_93 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_553 = _rdata_T_552 | _rdata_T_392; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_231 = 12'hb78 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_393 = _rdata_T_231 ? perfCnts_120 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_554 = _rdata_T_553 | _rdata_T_393; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_232 = 12'hb58 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_394 = _rdata_T_232 ? perfCnts_88 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_555 = _rdata_T_554 | _rdata_T_394; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_233 = 12'hb7d == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_395 = _rdata_T_233 ? perfCnts_125 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_556 = _rdata_T_555 | _rdata_T_395; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_234 = 12'hb4e == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_396 = _rdata_T_234 ? perfCnts_78 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_557 = _rdata_T_556 | _rdata_T_396; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_235 = 12'hb21 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_397 = _rdata_T_235 ? perfCnts_33 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_558 = _rdata_T_557 | _rdata_T_397; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_236 = 12'h304 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_398 = _rdata_T_236 ? mie : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_559 = _rdata_T_558 | _rdata_T_398; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_237 = 12'hb01 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_399 = _rdata_T_237 ? perfCnts_1 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_560 = _rdata_T_559 | _rdata_T_399; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_238 = 12'hb0b == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_400 = _rdata_T_238 ? perfCnts_11 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_561 = _rdata_T_560 | _rdata_T_400; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_239 = 12'hb2b == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_401 = _rdata_T_239 ? perfCnts_43 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_562 = _rdata_T_561 | _rdata_T_401; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_240 = 12'hb7a == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_402 = _rdata_T_240 ? perfCnts_122 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_563 = _rdata_T_562 | _rdata_T_402; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_241 = 12'hb4b == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_403 = _rdata_T_241 ? perfCnts_75 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_564 = _rdata_T_563 | _rdata_T_403; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_242 = 12'hb77 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_404 = _rdata_T_242 ? perfCnts_119 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_565 = _rdata_T_564 | _rdata_T_404; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_243 = 12'h3b3 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_405 = _rdata_T_243 ? pmpaddr3 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_566 = _rdata_T_565 | _rdata_T_405; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_244 = 12'hb5a == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_406 = _rdata_T_244 ? perfCnts_90 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_567 = _rdata_T_566 | _rdata_T_406; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_245 = 12'hb17 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_407 = _rdata_T_245 ? perfCnts_23 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_568 = _rdata_T_567 | _rdata_T_407; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_246 = 12'hb7f == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_408 = _rdata_T_246 ? perfCnts_127 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_569 = _rdata_T_568 | _rdata_T_408; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_247 = 12'hb28 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_409 = _rdata_T_247 ? perfCnts_40 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_570 = _rdata_T_569 | _rdata_T_409; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_248 = 12'hb50 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_410 = _rdata_T_248 ? perfCnts_80 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_571 = _rdata_T_570 | _rdata_T_410; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_249 = 12'hb37 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_411 = _rdata_T_249 ? perfCnts_55 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_572 = _rdata_T_571 | _rdata_T_411; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_250 = 12'hb08 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_412 = _rdata_T_250 ? perfCnts_8 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_573 = _rdata_T_572 | _rdata_T_412; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_251 = 12'h143 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_413 = _rdata_T_251 ? stval : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_574 = _rdata_T_573 | _rdata_T_413; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_252 = 12'hb6b == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_414 = _rdata_T_252 ? perfCnts_107 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_575 = _rdata_T_574 | _rdata_T_414; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_253 = 12'hb3a == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_415 = _rdata_T_253 ? perfCnts_58 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_576 = _rdata_T_575 | _rdata_T_415; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_254 = 12'h301 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_416 = _rdata_T_254 ? misa : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_577 = _rdata_T_576 | _rdata_T_416; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_255 = 12'hb70 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_417 = _rdata_T_255 ? perfCnts_112 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_578 = _rdata_T_577 | _rdata_T_417; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_256 = 12'hb1a == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_418 = _rdata_T_256 ? perfCnts_26 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_579 = _rdata_T_578 | _rdata_T_418; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_257 = 12'hb5f == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_419 = _rdata_T_257 ? perfCnts_95 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_580 = _rdata_T_579 | _rdata_T_419; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_258 = 12'hb73 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_420 = _rdata_T_258 ? perfCnts_115 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_581 = _rdata_T_580 | _rdata_T_420; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_259 = 12'hb33 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_421 = _rdata_T_259 ? perfCnts_51 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_582 = _rdata_T_581 | _rdata_T_421; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_260 = 12'h300 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_422 = _rdata_T_260 ? mstatus : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_583 = _rdata_T_582 | _rdata_T_422; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_261 = 12'hb13 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_423 = _rdata_T_261 ? perfCnts_19 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_584 = _rdata_T_583 | _rdata_T_423; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_262 = 12'h3b0 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_424 = _rdata_T_262 ? pmpaddr0 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_585 = _rdata_T_584 | _rdata_T_424; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_263 = 12'hb3e == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_425 = _rdata_T_263 ? perfCnts_62 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_586 = _rdata_T_585 | _rdata_T_425; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_264 = 12'hb6f == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_426 = _rdata_T_264 ? perfCnts_111 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_587 = _rdata_T_586 | _rdata_T_426; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_265 = 12'hb1e == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_427 = _rdata_T_265 ? perfCnts_30 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_588 = _rdata_T_587 | _rdata_T_427; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_266 = 12'hb53 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_428 = _rdata_T_266 ? perfCnts_83 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_589 = _rdata_T_588 | _rdata_T_428; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_267 = 12'h344 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_429 = _rdata_T_267 ? _GEN_332 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_590 = _rdata_T_589 | _rdata_T_429; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_268 = 12'hb62 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_430 = _rdata_T_268 ? perfCnts_98 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_591 = _rdata_T_590 | _rdata_T_430; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_269 = 12'hb00 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_431 = _rdata_T_269 ? perfCnts_0 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_592 = _rdata_T_591 | _rdata_T_431; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_270 = 12'hb7e == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_432 = _rdata_T_270 ? perfCnts_126 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_593 = _rdata_T_592 | _rdata_T_432; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_271 = 12'hb2f == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_433 = _rdata_T_271 ? perfCnts_47 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_594 = _rdata_T_593 | _rdata_T_433; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_272 = 12'hb05 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_434 = _rdata_T_272 ? perfCnts_5 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_595 = _rdata_T_594 | _rdata_T_434; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_273 = 12'hb22 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_435 = _rdata_T_273 ? perfCnts_34 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_596 = _rdata_T_595 | _rdata_T_435; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_274 = 12'hb48 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_436 = _rdata_T_274 ? perfCnts_72 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_597 = _rdata_T_596 | _rdata_T_436; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_275 = 12'hb42 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_437 = _rdata_T_275 ? perfCnts_66 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_598 = _rdata_T_597 | _rdata_T_437; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_276 = 12'hb0f == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_438 = _rdata_T_276 ? perfCnts_15 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_599 = _rdata_T_598 | _rdata_T_438; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_277 = 12'hb68 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_439 = _rdata_T_277 ? perfCnts_104 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_600 = _rdata_T_599 | _rdata_T_439; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_278 = 12'hb57 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_440 = _rdata_T_278 ? perfCnts_87 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_601 = _rdata_T_600 | _rdata_T_440; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_279 = 12'hb16 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_441 = _rdata_T_279 ? perfCnts_22 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_602 = _rdata_T_601 | _rdata_T_441; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_280 = 12'hb1b == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_442 = _rdata_T_280 ? perfCnts_27 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_603 = _rdata_T_602 | _rdata_T_442; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_281 = 12'hb2c == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_443 = _rdata_T_281 ? perfCnts_44 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_604 = _rdata_T_603 | _rdata_T_443; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_282 = 12'hb7b == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_444 = _rdata_T_282 ? perfCnts_123 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_605 = _rdata_T_604 | _rdata_T_444; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_283 = 12'hb4c == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_445 = _rdata_T_283 ? perfCnts_76 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_606 = _rdata_T_605 | _rdata_T_445; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_284 = 12'hb20 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_446 = _rdata_T_284 ? perfCnts_32 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_607 = _rdata_T_606 | _rdata_T_446; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_285 = 12'hb6c == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_447 = _rdata_T_285 ? perfCnts_108 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_608 = _rdata_T_607 | _rdata_T_447; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_286 = 12'hb02 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_448 = _rdata_T_286 ? perfCnts_2 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_609 = _rdata_T_608 | _rdata_T_448; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_287 = 12'hb67 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_449 = _rdata_T_287 ? perfCnts_103 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_610 = _rdata_T_609 | _rdata_T_449; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_288 = 12'hb31 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_450 = _rdata_T_288 ? perfCnts_49 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_611 = _rdata_T_610 | _rdata_T_450; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_289 = 12'hb3b == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_451 = _rdata_T_289 ? perfCnts_59 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_612 = _rdata_T_611 | _rdata_T_451; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_290 = 12'h3a3 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_452 = _rdata_T_290 ? pmpcfg3 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_613 = _rdata_T_612 | _rdata_T_452; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_291 = 12'hb45 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_453 = _rdata_T_291 ? perfCnts_69 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_614 = _rdata_T_613 | _rdata_T_453; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_292 = 12'hb36 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_454 = _rdata_T_292 ? perfCnts_54 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_615 = _rdata_T_614 | _rdata_T_454; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_293 = 12'hb0c == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_455 = _rdata_T_293 ? perfCnts_12 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_616 = _rdata_T_615 | _rdata_T_455; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_294 = 12'h303 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_456 = _rdata_T_294 ? mideleg : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_617 = _rdata_T_616 | _rdata_T_456; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_295 = 12'hb5b == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_457 = _rdata_T_295 ? perfCnts_91 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_618 = _rdata_T_617 | _rdata_T_457; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_296 = 12'hb27 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_458 = _rdata_T_296 ? perfCnts_39 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_619 = _rdata_T_618 | _rdata_T_458; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_297 = 12'hb25 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_459 = _rdata_T_297 ? perfCnts_37 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_620 = _rdata_T_619 | _rdata_T_459; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_298 = 12'h3b2 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_460 = _rdata_T_298 ? pmpaddr2 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_621 = _rdata_T_620 | _rdata_T_460; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_299 = 12'hb07 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_461 = _rdata_T_299 ? perfCnts_7 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_622 = _rdata_T_621 | _rdata_T_461; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_300 = 12'hf13 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _rdata_T_301 = 12'hb76 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_463 = _rdata_T_301 ? perfCnts_118 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_624 = _rdata_T_622 | _rdata_T_463; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_302 = 12'hb60 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_464 = _rdata_T_302 ? perfCnts_96 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_625 = _rdata_T_624 | _rdata_T_464; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_303 = 12'h3a1 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_465 = _rdata_T_303 ? pmpcfg1 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_626 = _rdata_T_625 | _rdata_T_465; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_304 = 12'hb56 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_466 = _rdata_T_304 ? perfCnts_86 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_627 = _rdata_T_626 | _rdata_T_466; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_305 = 12'h340 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_467 = _rdata_T_305 ? mscratch : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_628 = _rdata_T_627 | _rdata_T_467; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_306 = 12'hb65 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_468 = _rdata_T_306 ? perfCnts_101 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_629 = _rdata_T_628 | _rdata_T_468; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_307 = 12'hb72 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_469 = _rdata_T_307 ? perfCnts_114 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_630 = _rdata_T_629 | _rdata_T_469; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_308 = 12'hf14 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _rdata_T_309 = 12'h341 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_471 = _rdata_T_309 ? mepc : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_632 = _rdata_T_630 | _rdata_T_471; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_310 = 12'h343 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_472 = _rdata_T_310 ? mtval : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_633 = _rdata_T_632 | _rdata_T_472; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_311 = 12'h106 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_473 = _rdata_T_311 ? scounteren : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_634 = _rdata_T_633 | _rdata_T_473; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_312 = 12'hb61 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_474 = _rdata_T_312 ? perfCnts_97 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_635 = _rdata_T_634 | _rdata_T_474; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_313 = 12'h3a0 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_475 = _rdata_T_313 ? pmpcfg0 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_636 = _rdata_T_635 | _rdata_T_475; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_314 = 12'hb1f == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_476 = _rdata_T_314 ? perfCnts_31 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_637 = _rdata_T_636 | _rdata_T_476; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_315 = 12'hb52 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_477 = _rdata_T_315 ? perfCnts_82 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_638 = _rdata_T_637 | _rdata_T_477; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_316 = 12'hb30 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_478 = _rdata_T_316 ? perfCnts_48 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_639 = _rdata_T_638 | _rdata_T_478; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_317 = 12'h142 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_479 = _rdata_T_317 ? scause : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_640 = _rdata_T_639 | _rdata_T_479; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_318 = 12'hb3f == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_480 = _rdata_T_318 ? perfCnts_63 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_641 = _rdata_T_640 | _rdata_T_480; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_319 = 12'hb41 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_481 = _rdata_T_319 ? perfCnts_65 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_642 = _rdata_T_641 | _rdata_T_481; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_320 = 12'hb47 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_482 = _rdata_T_320 ? perfCnts_71 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_643 = _rdata_T_642 | _rdata_T_482; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_321 = 12'hb12 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_483 = _rdata_T_321 ? perfCnts_18 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_644 = _rdata_T_643 | _rdata_T_483; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_322 = 12'hb32 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_484 = _rdata_T_322 ? perfCnts_50 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_645 = _rdata_T_644 | _rdata_T_484; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_323 = 12'hb10 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_485 = _rdata_T_323 ? perfCnts_16 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] rdata = _rdata_T_645 | _rdata_T_485; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _wdata_T = rdata | io_in_bits_src1; // @[src/main/scala/nutcore/backend/fu/CSR.scala 462:30]
  wire [63:0] _wdata_T_1 = ~io_in_bits_src1; // @[src/main/scala/nutcore/backend/fu/CSR.scala 463:32]
  wire [63:0] _wdata_T_2 = rdata & _wdata_T_1; // @[src/main/scala/nutcore/backend/fu/CSR.scala 463:30]
  wire [63:0] _wdata_T_3 = rdata | csri; // @[src/main/scala/nutcore/backend/fu/CSR.scala 465:30]
  wire [63:0] _wdata_T_4 = ~csri; // @[src/main/scala/nutcore/backend/fu/CSR.scala 466:32]
  wire [63:0] _wdata_T_5 = rdata & _wdata_T_4; // @[src/main/scala/nutcore/backend/fu/CSR.scala 466:30]
  wire  _wdata_T_6 = 7'h1 == io_in_bits_func; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _wdata_T_7 = 7'h2 == io_in_bits_func; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _wdata_T_8 = 7'h3 == io_in_bits_func; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _wdata_T_9 = 7'h5 == io_in_bits_func; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _wdata_T_10 = 7'h6 == io_in_bits_func; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _wdata_T_11 = 7'h7 == io_in_bits_func; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _wdata_T_12 = _wdata_T_6 ? io_in_bits_src1 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _wdata_T_13 = _wdata_T_7 ? _wdata_T : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _wdata_T_14 = _wdata_T_8 ? _wdata_T_2 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _wdata_T_15 = _wdata_T_9 ? csri : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _wdata_T_16 = _wdata_T_10 ? _wdata_T_3 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _wdata_T_17 = _wdata_T_11 ? _wdata_T_5 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _wdata_T_18 = _wdata_T_12 | _wdata_T_13; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _wdata_T_19 = _wdata_T_18 | _wdata_T_14; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _wdata_T_20 = _wdata_T_19 | _wdata_T_15; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _wdata_T_21 = _wdata_T_20 | _wdata_T_16; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] wdata = _wdata_T_21 | _wdata_T_17; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  satpLegalMode = wdata[63:60] == 4'h0 | wdata[63:60] == 4'h8; // @[src/main/scala/nutcore/backend/fu/CSR.scala 470:69]
  wire  wen = io_in_valid & io_in_bits_func != 7'h0 & (addr != 12'h180 | satpLegalMode); // @[src/main/scala/nutcore/backend/fu/CSR.scala 473:47]
  wire  isIllegalMode = priviledgeMode < addr[9:8]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 474:39]
  wire  justRead = (io_in_bits_func == 7'h2 | io_in_bits_func == 7'h6) & io_in_bits_src1 == 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 475:70]
  wire  isIllegalWrite = wen & addr[11:10] == 2'h3 & ~justRead; // @[src/main/scala/nutcore/backend/fu/CSR.scala 476:58]
  wire  isIllegalAccess = isIllegalMode | isIllegalWrite; // @[src/main/scala/nutcore/backend/fu/CSR.scala 477:39]
  wire  _T_693 = wen & ~isIllegalAccess; // @[src/main/scala/nutcore/backend/fu/CSR.scala 479:51]
  wire  _T_710 = addr == 12'h180; // @[src/main/scala/utils/RegMap.scala 50:65]
  wire [63:0] _pmpaddr1_T = wdata & 64'h3fffffff; // @[src/main/scala/utils/BitUtils.scala 34:14]
  wire [63:0] _pmpaddr1_T_2 = pmpaddr1 & 64'hffffffffc0000000; // @[src/main/scala/utils/BitUtils.scala 34:37]
  wire [63:0] _pmpaddr1_T_3 = _pmpaddr1_T | _pmpaddr1_T_2; // @[src/main/scala/utils/BitUtils.scala 34:26]
  wire  _T_740 = addr == 12'h302; // @[src/main/scala/utils/RegMap.scala 50:65]
  wire [63:0] _medeleg_T = wdata & 64'hbbff; // @[src/main/scala/utils/BitUtils.scala 34:14]
  wire [63:0] _medeleg_T_2 = medeleg & 64'hffffffffffff4400; // @[src/main/scala/utils/BitUtils.scala 34:37]
  wire [63:0] _medeleg_T_3 = _medeleg_T | _medeleg_T_2; // @[src/main/scala/utils/BitUtils.scala 34:26]
  wire [63:0] _GEN_32 = _T_693 & addr == 12'h141 ? wdata : sepc; // @[src/main/scala/nutcore/backend/fu/CSR.scala 338:21 src/main/scala/utils/RegMap.scala 50:{72,76}]
  wire [63:0] _GEN_34 = _T_693 & addr == 12'h342 ? wdata : mcause; // @[src/main/scala/nutcore/backend/fu/CSR.scala 254:23 src/main/scala/utils/RegMap.scala 50:{72,76}]
  wire [63:0] _mie_T = wdata & sieMask; // @[src/main/scala/utils/BitUtils.scala 34:14]
  wire [63:0] _mie_T_1 = ~sieMask; // @[src/main/scala/utils/BitUtils.scala 34:39]
  wire [63:0] _mie_T_2 = mie & _mie_T_1; // @[src/main/scala/utils/BitUtils.scala 34:37]
  wire [63:0] _mie_T_3 = _mie_T | _mie_T_2; // @[src/main/scala/utils/BitUtils.scala 34:26]
  wire [63:0] _mstatus_T = wdata & 64'hc6122; // @[src/main/scala/utils/BitUtils.scala 34:14]
  wire [63:0] _mstatus_T_2 = mstatus & 64'hfffffffffff39edd; // @[src/main/scala/utils/BitUtils.scala 34:37]
  wire [63:0] _mstatus_T_3 = _mstatus_T | _mstatus_T_2; // @[src/main/scala/utils/BitUtils.scala 34:26]
  wire [1:0] mstatus_mstatusOld_fs = _mstatus_T_3[14:13]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 301:47]
  wire [63:0] mstatus_mstatusNew = {mstatus_mstatusOld_fs == 2'h3,_mstatus_T_3[62:0]}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 302:25]
  wire [63:0] _GEN_53 = _T_693 & addr == 12'h100 ? mstatus_mstatusNew : mstatus; // @[src/main/scala/nutcore/backend/fu/CSR.scala 278:24 src/main/scala/utils/RegMap.scala 50:{72,76}]
  wire [63:0] _pmpaddr3_T_2 = pmpaddr3 & 64'hffffffffc0000000; // @[src/main/scala/utils/BitUtils.scala 34:37]
  wire [63:0] _pmpaddr3_T_3 = _pmpaddr1_T | _pmpaddr3_T_2; // @[src/main/scala/utils/BitUtils.scala 34:26]
  wire [63:0] _GEN_88 = _T_693 & addr == 12'h143 ? wdata : stval; // @[src/main/scala/nutcore/backend/fu/CSR.scala 340:18 src/main/scala/utils/RegMap.scala 50:{72,76}]
  wire [1:0] mstatus_mstatusOld_1_fs = wdata[14:13]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 301:47]
  wire [63:0] mstatus_mstatusNew_1 = {mstatus_mstatusOld_1_fs == 2'h3,wdata[62:0]}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 302:25]
  wire [63:0] _GEN_97 = _T_693 & addr == 12'h300 ? mstatus_mstatusNew_1 : _GEN_53; // @[src/main/scala/utils/RegMap.scala 50:{72,76}]
  wire [63:0] _pmpaddr0_T_2 = pmpaddr0 & 64'hffffffffc0000000; // @[src/main/scala/utils/BitUtils.scala 34:37]
  wire [63:0] _pmpaddr0_T_3 = _pmpaddr1_T | _pmpaddr0_T_2; // @[src/main/scala/utils/BitUtils.scala 34:26]
  wire [63:0] _mideleg_T = wdata & 64'h222; // @[src/main/scala/utils/BitUtils.scala 34:14]
  wire [63:0] _mideleg_T_2 = mideleg & 64'hfffffffffffffddd; // @[src/main/scala/utils/BitUtils.scala 34:37]
  wire [63:0] _mideleg_T_3 = _mideleg_T | _mideleg_T_2; // @[src/main/scala/utils/BitUtils.scala 34:26]
  wire [63:0] _pmpaddr2_T_2 = pmpaddr2 & 64'hffffffffc0000000; // @[src/main/scala/utils/BitUtils.scala 34:37]
  wire [63:0] _pmpaddr2_T_3 = _pmpaddr1_T | _pmpaddr2_T_2; // @[src/main/scala/utils/BitUtils.scala 34:26]
  wire [63:0] _GEN_143 = _T_693 & addr == 12'h341 ? wdata : mepc; // @[src/main/scala/nutcore/backend/fu/CSR.scala 256:21 src/main/scala/utils/RegMap.scala 50:{72,76}]
  wire [63:0] _GEN_144 = _T_693 & addr == 12'h343 ? wdata : mtval; // @[src/main/scala/nutcore/backend/fu/CSR.scala 255:22 src/main/scala/utils/RegMap.scala 50:{72,76}]
  wire [63:0] _GEN_151 = _T_693 & addr == 12'h142 ? wdata : scause; // @[src/main/scala/nutcore/backend/fu/CSR.scala 339:23 src/main/scala/utils/RegMap.scala 50:{72,76}]
  wire  _isIllegalAddr_illegalAddr_T_1 = _rdata_T_162 ? 1'h0 : 1'h1; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_3 = _rdata_T_163 ? 1'h0 : _isIllegalAddr_illegalAddr_T_1; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_5 = _rdata_T_164 ? 1'h0 : _isIllegalAddr_illegalAddr_T_3; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_7 = _rdata_T_165 ? 1'h0 : _isIllegalAddr_illegalAddr_T_5; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_9 = _rdata_T_166 ? 1'h0 : _isIllegalAddr_illegalAddr_T_7; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_11 = _rdata_T_167 ? 1'h0 : _isIllegalAddr_illegalAddr_T_9; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_13 = _rdata_T_168 ? 1'h0 : _isIllegalAddr_illegalAddr_T_11; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_15 = _rdata_T_169 ? 1'h0 : _isIllegalAddr_illegalAddr_T_13; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_17 = _rdata_T_170 ? 1'h0 : _isIllegalAddr_illegalAddr_T_15; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_19 = _rdata_T_171 ? 1'h0 : _isIllegalAddr_illegalAddr_T_17; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_21 = _rdata_T_172 ? 1'h0 : _isIllegalAddr_illegalAddr_T_19; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_23 = _rdata_T_173 ? 1'h0 : _isIllegalAddr_illegalAddr_T_21; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_25 = _rdata_T_174 ? 1'h0 : _isIllegalAddr_illegalAddr_T_23; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_27 = _rdata_T_175 ? 1'h0 : _isIllegalAddr_illegalAddr_T_25; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_29 = _rdata_T_176 ? 1'h0 : _isIllegalAddr_illegalAddr_T_27; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_31 = _rdata_T_177 ? 1'h0 : _isIllegalAddr_illegalAddr_T_29; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_33 = _rdata_T_178 ? 1'h0 : _isIllegalAddr_illegalAddr_T_31; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_35 = _rdata_T_179 ? 1'h0 : _isIllegalAddr_illegalAddr_T_33; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_37 = _rdata_T_180 ? 1'h0 : _isIllegalAddr_illegalAddr_T_35; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_39 = _rdata_T_181 ? 1'h0 : _isIllegalAddr_illegalAddr_T_37; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_41 = _rdata_T_182 ? 1'h0 : _isIllegalAddr_illegalAddr_T_39; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_43 = _rdata_T_183 ? 1'h0 : _isIllegalAddr_illegalAddr_T_41; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_45 = _rdata_T_184 ? 1'h0 : _isIllegalAddr_illegalAddr_T_43; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_47 = _rdata_T_185 ? 1'h0 : _isIllegalAddr_illegalAddr_T_45; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_49 = _rdata_T_186 ? 1'h0 : _isIllegalAddr_illegalAddr_T_47; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_51 = _rdata_T_187 ? 1'h0 : _isIllegalAddr_illegalAddr_T_49; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_53 = _rdata_T_188 ? 1'h0 : _isIllegalAddr_illegalAddr_T_51; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_55 = _rdata_T_189 ? 1'h0 : _isIllegalAddr_illegalAddr_T_53; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_57 = _rdata_T_190 ? 1'h0 : _isIllegalAddr_illegalAddr_T_55; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_59 = _rdata_T_191 ? 1'h0 : _isIllegalAddr_illegalAddr_T_57; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_61 = _rdata_T_192 ? 1'h0 : _isIllegalAddr_illegalAddr_T_59; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_63 = _rdata_T_193 ? 1'h0 : _isIllegalAddr_illegalAddr_T_61; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_65 = _rdata_T_194 ? 1'h0 : _isIllegalAddr_illegalAddr_T_63; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_67 = _rdata_T_195 ? 1'h0 : _isIllegalAddr_illegalAddr_T_65; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_69 = _rdata_T_196 ? 1'h0 : _isIllegalAddr_illegalAddr_T_67; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_71 = _rdata_T_197 ? 1'h0 : _isIllegalAddr_illegalAddr_T_69; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_73 = _rdata_T_198 ? 1'h0 : _isIllegalAddr_illegalAddr_T_71; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_75 = _rdata_T_199 ? 1'h0 : _isIllegalAddr_illegalAddr_T_73; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_77 = _rdata_T_200 ? 1'h0 : _isIllegalAddr_illegalAddr_T_75; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_79 = _rdata_T_201 ? 1'h0 : _isIllegalAddr_illegalAddr_T_77; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_81 = _rdata_T_202 ? 1'h0 : _isIllegalAddr_illegalAddr_T_79; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_83 = _rdata_T_203 ? 1'h0 : _isIllegalAddr_illegalAddr_T_81; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_85 = _rdata_T_204 ? 1'h0 : _isIllegalAddr_illegalAddr_T_83; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_87 = _rdata_T_205 ? 1'h0 : _isIllegalAddr_illegalAddr_T_85; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_89 = _rdata_T_206 ? 1'h0 : _isIllegalAddr_illegalAddr_T_87; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_91 = _rdata_T_207 ? 1'h0 : _isIllegalAddr_illegalAddr_T_89; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_93 = _rdata_T_208 ? 1'h0 : _isIllegalAddr_illegalAddr_T_91; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_95 = _rdata_T_209 ? 1'h0 : _isIllegalAddr_illegalAddr_T_93; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_97 = _rdata_T_210 ? 1'h0 : _isIllegalAddr_illegalAddr_T_95; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_99 = _rdata_T_211 ? 1'h0 : _isIllegalAddr_illegalAddr_T_97; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_101 = _rdata_T_212 ? 1'h0 : _isIllegalAddr_illegalAddr_T_99; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_103 = _rdata_T_213 ? 1'h0 : _isIllegalAddr_illegalAddr_T_101; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_105 = _rdata_T_214 ? 1'h0 : _isIllegalAddr_illegalAddr_T_103; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_107 = _rdata_T_215 ? 1'h0 : _isIllegalAddr_illegalAddr_T_105; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_109 = _rdata_T_216 ? 1'h0 : _isIllegalAddr_illegalAddr_T_107; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_111 = _rdata_T_217 ? 1'h0 : _isIllegalAddr_illegalAddr_T_109; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_113 = _rdata_T_218 ? 1'h0 : _isIllegalAddr_illegalAddr_T_111; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_115 = _rdata_T_219 ? 1'h0 : _isIllegalAddr_illegalAddr_T_113; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_117 = _rdata_T_220 ? 1'h0 : _isIllegalAddr_illegalAddr_T_115; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_119 = _rdata_T_221 ? 1'h0 : _isIllegalAddr_illegalAddr_T_117; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_121 = _rdata_T_222 ? 1'h0 : _isIllegalAddr_illegalAddr_T_119; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_123 = _rdata_T_223 ? 1'h0 : _isIllegalAddr_illegalAddr_T_121; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_125 = _rdata_T_224 ? 1'h0 : _isIllegalAddr_illegalAddr_T_123; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_127 = _rdata_T_225 ? 1'h0 : _isIllegalAddr_illegalAddr_T_125; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_129 = _rdata_T_226 ? 1'h0 : _isIllegalAddr_illegalAddr_T_127; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_131 = _rdata_T_227 ? 1'h0 : _isIllegalAddr_illegalAddr_T_129; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_133 = _rdata_T_228 ? 1'h0 : _isIllegalAddr_illegalAddr_T_131; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_135 = _rdata_T_229 ? 1'h0 : _isIllegalAddr_illegalAddr_T_133; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_137 = _rdata_T_230 ? 1'h0 : _isIllegalAddr_illegalAddr_T_135; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_139 = _rdata_T_231 ? 1'h0 : _isIllegalAddr_illegalAddr_T_137; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_141 = _rdata_T_232 ? 1'h0 : _isIllegalAddr_illegalAddr_T_139; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_143 = _rdata_T_233 ? 1'h0 : _isIllegalAddr_illegalAddr_T_141; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_145 = _rdata_T_234 ? 1'h0 : _isIllegalAddr_illegalAddr_T_143; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_147 = _rdata_T_235 ? 1'h0 : _isIllegalAddr_illegalAddr_T_145; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_149 = _rdata_T_236 ? 1'h0 : _isIllegalAddr_illegalAddr_T_147; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_151 = _rdata_T_237 ? 1'h0 : _isIllegalAddr_illegalAddr_T_149; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_153 = _rdata_T_238 ? 1'h0 : _isIllegalAddr_illegalAddr_T_151; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_155 = _rdata_T_239 ? 1'h0 : _isIllegalAddr_illegalAddr_T_153; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_157 = _rdata_T_240 ? 1'h0 : _isIllegalAddr_illegalAddr_T_155; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_159 = _rdata_T_241 ? 1'h0 : _isIllegalAddr_illegalAddr_T_157; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_161 = _rdata_T_242 ? 1'h0 : _isIllegalAddr_illegalAddr_T_159; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_163 = _rdata_T_243 ? 1'h0 : _isIllegalAddr_illegalAddr_T_161; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_165 = _rdata_T_244 ? 1'h0 : _isIllegalAddr_illegalAddr_T_163; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_167 = _rdata_T_245 ? 1'h0 : _isIllegalAddr_illegalAddr_T_165; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_169 = _rdata_T_246 ? 1'h0 : _isIllegalAddr_illegalAddr_T_167; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_171 = _rdata_T_247 ? 1'h0 : _isIllegalAddr_illegalAddr_T_169; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_173 = _rdata_T_248 ? 1'h0 : _isIllegalAddr_illegalAddr_T_171; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_175 = _rdata_T_249 ? 1'h0 : _isIllegalAddr_illegalAddr_T_173; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_177 = _rdata_T_250 ? 1'h0 : _isIllegalAddr_illegalAddr_T_175; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_179 = _rdata_T_251 ? 1'h0 : _isIllegalAddr_illegalAddr_T_177; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_181 = _rdata_T_252 ? 1'h0 : _isIllegalAddr_illegalAddr_T_179; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_183 = _rdata_T_253 ? 1'h0 : _isIllegalAddr_illegalAddr_T_181; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_185 = _rdata_T_254 ? 1'h0 : _isIllegalAddr_illegalAddr_T_183; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_187 = _rdata_T_255 ? 1'h0 : _isIllegalAddr_illegalAddr_T_185; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_189 = _rdata_T_256 ? 1'h0 : _isIllegalAddr_illegalAddr_T_187; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_191 = _rdata_T_257 ? 1'h0 : _isIllegalAddr_illegalAddr_T_189; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_193 = _rdata_T_258 ? 1'h0 : _isIllegalAddr_illegalAddr_T_191; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_195 = _rdata_T_259 ? 1'h0 : _isIllegalAddr_illegalAddr_T_193; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_197 = _rdata_T_260 ? 1'h0 : _isIllegalAddr_illegalAddr_T_195; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_199 = _rdata_T_261 ? 1'h0 : _isIllegalAddr_illegalAddr_T_197; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_201 = _rdata_T_262 ? 1'h0 : _isIllegalAddr_illegalAddr_T_199; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_203 = _rdata_T_263 ? 1'h0 : _isIllegalAddr_illegalAddr_T_201; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_205 = _rdata_T_264 ? 1'h0 : _isIllegalAddr_illegalAddr_T_203; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_207 = _rdata_T_265 ? 1'h0 : _isIllegalAddr_illegalAddr_T_205; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_209 = _rdata_T_266 ? 1'h0 : _isIllegalAddr_illegalAddr_T_207; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_211 = _rdata_T_267 ? 1'h0 : _isIllegalAddr_illegalAddr_T_209; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_213 = _rdata_T_268 ? 1'h0 : _isIllegalAddr_illegalAddr_T_211; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_215 = _rdata_T_269 ? 1'h0 : _isIllegalAddr_illegalAddr_T_213; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_217 = _rdata_T_270 ? 1'h0 : _isIllegalAddr_illegalAddr_T_215; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_219 = _rdata_T_271 ? 1'h0 : _isIllegalAddr_illegalAddr_T_217; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_221 = _rdata_T_272 ? 1'h0 : _isIllegalAddr_illegalAddr_T_219; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_223 = _rdata_T_273 ? 1'h0 : _isIllegalAddr_illegalAddr_T_221; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_225 = _rdata_T_274 ? 1'h0 : _isIllegalAddr_illegalAddr_T_223; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_227 = _rdata_T_275 ? 1'h0 : _isIllegalAddr_illegalAddr_T_225; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_229 = _rdata_T_276 ? 1'h0 : _isIllegalAddr_illegalAddr_T_227; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_231 = _rdata_T_277 ? 1'h0 : _isIllegalAddr_illegalAddr_T_229; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_233 = _rdata_T_278 ? 1'h0 : _isIllegalAddr_illegalAddr_T_231; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_235 = _rdata_T_279 ? 1'h0 : _isIllegalAddr_illegalAddr_T_233; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_237 = _rdata_T_280 ? 1'h0 : _isIllegalAddr_illegalAddr_T_235; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_239 = _rdata_T_281 ? 1'h0 : _isIllegalAddr_illegalAddr_T_237; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_241 = _rdata_T_282 ? 1'h0 : _isIllegalAddr_illegalAddr_T_239; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_243 = _rdata_T_283 ? 1'h0 : _isIllegalAddr_illegalAddr_T_241; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_245 = _rdata_T_284 ? 1'h0 : _isIllegalAddr_illegalAddr_T_243; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_247 = _rdata_T_285 ? 1'h0 : _isIllegalAddr_illegalAddr_T_245; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_249 = _rdata_T_286 ? 1'h0 : _isIllegalAddr_illegalAddr_T_247; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_251 = _rdata_T_287 ? 1'h0 : _isIllegalAddr_illegalAddr_T_249; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_253 = _rdata_T_288 ? 1'h0 : _isIllegalAddr_illegalAddr_T_251; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_255 = _rdata_T_289 ? 1'h0 : _isIllegalAddr_illegalAddr_T_253; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_257 = _rdata_T_290 ? 1'h0 : _isIllegalAddr_illegalAddr_T_255; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_259 = _rdata_T_291 ? 1'h0 : _isIllegalAddr_illegalAddr_T_257; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_261 = _rdata_T_292 ? 1'h0 : _isIllegalAddr_illegalAddr_T_259; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_263 = _rdata_T_293 ? 1'h0 : _isIllegalAddr_illegalAddr_T_261; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_265 = _rdata_T_294 ? 1'h0 : _isIllegalAddr_illegalAddr_T_263; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_267 = _rdata_T_295 ? 1'h0 : _isIllegalAddr_illegalAddr_T_265; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_269 = _rdata_T_296 ? 1'h0 : _isIllegalAddr_illegalAddr_T_267; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_271 = _rdata_T_297 ? 1'h0 : _isIllegalAddr_illegalAddr_T_269; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_273 = _rdata_T_298 ? 1'h0 : _isIllegalAddr_illegalAddr_T_271; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_275 = _rdata_T_299 ? 1'h0 : _isIllegalAddr_illegalAddr_T_273; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_277 = _rdata_T_300 ? 1'h0 : _isIllegalAddr_illegalAddr_T_275; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_279 = _rdata_T_301 ? 1'h0 : _isIllegalAddr_illegalAddr_T_277; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_281 = _rdata_T_302 ? 1'h0 : _isIllegalAddr_illegalAddr_T_279; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_283 = _rdata_T_303 ? 1'h0 : _isIllegalAddr_illegalAddr_T_281; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_285 = _rdata_T_304 ? 1'h0 : _isIllegalAddr_illegalAddr_T_283; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_287 = _rdata_T_305 ? 1'h0 : _isIllegalAddr_illegalAddr_T_285; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_289 = _rdata_T_306 ? 1'h0 : _isIllegalAddr_illegalAddr_T_287; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_291 = _rdata_T_307 ? 1'h0 : _isIllegalAddr_illegalAddr_T_289; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_293 = _rdata_T_308 ? 1'h0 : _isIllegalAddr_illegalAddr_T_291; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_295 = _rdata_T_309 ? 1'h0 : _isIllegalAddr_illegalAddr_T_293; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_297 = _rdata_T_310 ? 1'h0 : _isIllegalAddr_illegalAddr_T_295; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_299 = _rdata_T_311 ? 1'h0 : _isIllegalAddr_illegalAddr_T_297; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_301 = _rdata_T_312 ? 1'h0 : _isIllegalAddr_illegalAddr_T_299; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_303 = _rdata_T_313 ? 1'h0 : _isIllegalAddr_illegalAddr_T_301; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_305 = _rdata_T_314 ? 1'h0 : _isIllegalAddr_illegalAddr_T_303; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_307 = _rdata_T_315 ? 1'h0 : _isIllegalAddr_illegalAddr_T_305; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_309 = _rdata_T_316 ? 1'h0 : _isIllegalAddr_illegalAddr_T_307; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_311 = _rdata_T_317 ? 1'h0 : _isIllegalAddr_illegalAddr_T_309; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_313 = _rdata_T_318 ? 1'h0 : _isIllegalAddr_illegalAddr_T_311; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_315 = _rdata_T_319 ? 1'h0 : _isIllegalAddr_illegalAddr_T_313; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_317 = _rdata_T_320 ? 1'h0 : _isIllegalAddr_illegalAddr_T_315; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_319 = _rdata_T_321 ? 1'h0 : _isIllegalAddr_illegalAddr_T_317; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_321 = _rdata_T_322 ? 1'h0 : _isIllegalAddr_illegalAddr_T_319; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  isIllegalAddr = _rdata_T_323 ? 1'h0 : _isIllegalAddr_illegalAddr_T_321; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  resetSatp = _T_710 & wen; // @[src/main/scala/nutcore/backend/fu/CSR.scala 481:35]
  wire [63:0] _mipReg_T = wdata & 64'h77f; // @[src/main/scala/utils/BitUtils.scala 34:14]
  wire [63:0] _mipReg_T_2 = mipReg & 64'hfffffffffffff880; // @[src/main/scala/utils/BitUtils.scala 34:37]
  wire [63:0] _mipReg_T_3 = _mipReg_T | _mipReg_T_2; // @[src/main/scala/utils/BitUtils.scala 34:26]
  wire [63:0] _mipReg_T_6 = mipReg & _mie_T_1; // @[src/main/scala/utils/BitUtils.scala 34:37]
  wire [63:0] _mipReg_T_7 = _mie_T | _mipReg_T_6; // @[src/main/scala/utils/BitUtils.scala 34:26]
  wire  _isEbreak_T_1 = io_in_bits_func == 7'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 494:46]
  wire  isEbreak = addr == 12'h1 & io_in_bits_func == 7'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 494:38]
  wire  isEcall = addr == 12'h0 & _isEbreak_T_1; // @[src/main/scala/nutcore/backend/fu/CSR.scala 495:36]
  wire  isMret = _T_740 & _isEbreak_T_1; // @[src/main/scala/nutcore/backend/fu/CSR.scala 496:36]
  wire  isSret = addr == 12'h102 & _isEbreak_T_1; // @[src/main/scala/nutcore/backend/fu/CSR.scala 497:36]
  wire  isUret = addr == 12'h2 & _isEbreak_T_1; // @[src/main/scala/nutcore/backend/fu/CSR.scala 498:36]
  reg [63:0] c; // @[src/main/scala/utils/GTimer.scala 24:20]
  wire [63:0] _c_T_1 = c + 64'h1; // @[src/main/scala/utils/GTimer.scala 25:12]
  wire  _T_1013 = wen & DISPLAY_ENABLE; // @[src/main/scala/utils/Debug.scala 55:16]
  wire  _T_1015 = ~reset; // @[src/main/scala/utils/Debug.scala 56:24]
  reg [63:0] c_1; // @[src/main/scala/utils/GTimer.scala 24:20]
  wire [63:0] _c_T_3 = c_1 + 64'h1; // @[src/main/scala/utils/GTimer.scala 25:12]
  reg [63:0] c_2; // @[src/main/scala/utils/GTimer.scala 24:20]
  wire [63:0] _c_T_5 = c_2 + 64'h1; // @[src/main/scala/utils/GTimer.scala 25:12]
  wire  hasInstrPageFault = io_cfIn_exceptionVec_12 & io_in_valid; // @[src/main/scala/nutcore/backend/fu/CSR.scala 555:63]
  wire  _T_1024 = hasInstrPageFault | io_dmemMMU_loadPF | io_dmemMMU_storePF; // @[src/main/scala/nutcore/backend/fu/CSR.scala 564:46]
  wire [38:0] _tval_T_1 = io_cfIn_pc + 39'h2; // @[src/main/scala/nutcore/backend/fu/CSR.scala 565:88]
  wire  tval_signBit = _tval_T_1[38]; // @[src/main/scala/utils/BitUtils.scala 41:20]
  wire [24:0] _tval_T_4 = tval_signBit ? 25'h1ffffff : 25'h0; // @[src/main/scala/utils/BitUtils.scala 42:46]
  wire [63:0] _tval_T_5 = {_tval_T_4,_tval_T_1}; // @[src/main/scala/utils/BitUtils.scala 42:41]
  wire  tval_signBit_1 = io_cfIn_pc[38]; // @[src/main/scala/utils/BitUtils.scala 41:20]
  wire [24:0] _tval_T_8 = tval_signBit_1 ? 25'h1ffffff : 25'h0; // @[src/main/scala/utils/BitUtils.scala 42:46]
  wire [63:0] _tval_T_9 = {_tval_T_8,io_cfIn_pc}; // @[src/main/scala/utils/BitUtils.scala 42:41]
  wire [63:0] _tval_T_10 = io_cfIn_crossPageIPFFix ? _tval_T_5 : _tval_T_9; // @[src/main/scala/nutcore/backend/fu/CSR.scala 565:42]
  wire  tval_signBit_2 = io_dmemMMU_addr[38]; // @[src/main/scala/utils/BitUtils.scala 41:20]
  wire [24:0] _tval_T_12 = tval_signBit_2 ? 25'h1ffffff : 25'h0; // @[src/main/scala/utils/BitUtils.scala 42:46]
  wire [63:0] _tval_T_13 = {_tval_T_12,io_dmemMMU_addr}; // @[src/main/scala/utils/BitUtils.scala 42:41]
  wire [63:0] tval = hasInstrPageFault ? _tval_T_10 : _tval_T_13; // @[src/main/scala/nutcore/backend/fu/CSR.scala 565:19]
  wire  _T_1025 = priviledgeMode == 2'h3; // @[src/main/scala/nutcore/backend/fu/CSR.scala 566:25]
  wire [63:0] _GEN_160 = priviledgeMode == 2'h3 ? tval : _GEN_144; // @[src/main/scala/nutcore/backend/fu/CSR.scala 566:35 567:13]
  wire [63:0] _GEN_161 = priviledgeMode == 2'h3 ? _GEN_88 : tval; // @[src/main/scala/nutcore/backend/fu/CSR.scala 566:35 569:13]
  reg [63:0] c_3; // @[src/main/scala/utils/GTimer.scala 24:20]
  wire [63:0] _c_T_7 = c_3 + 64'h1; // @[src/main/scala/utils/GTimer.scala 25:12]
  reg [63:0] c_4; // @[src/main/scala/utils/GTimer.scala 24:20]
  wire [63:0] _c_T_9 = c_4 + 64'h1; // @[src/main/scala/utils/GTimer.scala 25:12]
  wire [63:0] _GEN_162 = hasInstrPageFault | io_dmemMMU_loadPF | io_dmemMMU_storePF ? _GEN_160 : _GEN_144; // @[src/main/scala/nutcore/backend/fu/CSR.scala 564:67]
  wire [63:0] _GEN_163 = hasInstrPageFault | io_dmemMMU_loadPF | io_dmemMMU_storePF ? _GEN_161 : _GEN_88; // @[src/main/scala/nutcore/backend/fu/CSR.scala 564:67]
  wire  _T_1034 = io_cfIn_exceptionVec_4 | io_cfIn_exceptionVec_6; // @[src/main/scala/nutcore/backend/fu/CSR.scala 574:30]
  wire [38:0] dmemAddrMisalignedAddr = LSUADDR[38:0]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 543:36 561:28]
  wire  mtval_signBit = dmemAddrMisalignedAddr[38]; // @[src/main/scala/utils/BitUtils.scala 41:20]
  wire [24:0] _mtval_T_5 = mtval_signBit ? 25'h1ffffff : 25'h0; // @[src/main/scala/utils/BitUtils.scala 42:46]
  wire [63:0] _mtval_T_6 = {_mtval_T_5,dmemAddrMisalignedAddr}; // @[src/main/scala/utils/BitUtils.scala 42:41]
  reg [63:0] c_5; // @[src/main/scala/utils/GTimer.scala 24:20]
  wire [63:0] _c_T_11 = c_5 + 64'h1; // @[src/main/scala/utils/GTimer.scala 25:12]
  reg [63:0] c_6; // @[src/main/scala/utils/GTimer.scala 24:20]
  wire [63:0] _c_T_13 = c_6 + 64'h1; // @[src/main/scala/utils/GTimer.scala 25:12]
  wire [63:0] _GEN_164 = _T_1034 ? _mtval_T_6 : _GEN_162; // @[src/main/scala/nutcore/backend/fu/CSR.scala 575:3 576:11]
  wire  mipRaiseIntr_e_s = mip_e_s | meip_0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 598:31]
  wire [11:0] _ideleg_T = {mip_e_m,mip_e_h,mipRaiseIntr_e_s,mip_e_u,mip_t_m,mip_t_h,lo}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 600:41]
  wire [63:0] _GEN_333 = {{52'd0}, _ideleg_T}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 600:26]
  wire [63:0] ideleg = mideleg & _GEN_333; // @[src/main/scala/nutcore/backend/fu/CSR.scala 600:26]
  wire  _intrVecEnable_0_T = priviledgeMode == 2'h1; // @[src/main/scala/nutcore/backend/fu/CSR.scala 601:72]
  wire  _intrVecEnable_0_T_6 = priviledgeMode < 2'h3; // @[src/main/scala/nutcore/backend/fu/CSR.scala 602:106]
  wire  _intrVecEnable_0_T_7 = _T_1025 & mstatusStruct_ie_m | priviledgeMode < 2'h3; // @[src/main/scala/nutcore/backend/fu/CSR.scala 602:87]
  wire  intrVecEnable_0 = ideleg[0] ? priviledgeMode == 2'h1 & mstatusStruct_ie_s | priviledgeMode < 2'h1 :
    _intrVecEnable_0_T_7; // @[src/main/scala/nutcore/backend/fu/CSR.scala 601:51]
  wire  intrVecEnable_1 = ideleg[1] ? priviledgeMode == 2'h1 & mstatusStruct_ie_s | priviledgeMode < 2'h1 :
    _intrVecEnable_0_T_7; // @[src/main/scala/nutcore/backend/fu/CSR.scala 601:51]
  wire  intrVecEnable_2 = ideleg[2] ? priviledgeMode == 2'h1 & mstatusStruct_ie_s | priviledgeMode < 2'h1 :
    _intrVecEnable_0_T_7; // @[src/main/scala/nutcore/backend/fu/CSR.scala 601:51]
  wire  intrVecEnable_3 = ideleg[3] ? priviledgeMode == 2'h1 & mstatusStruct_ie_s | priviledgeMode < 2'h1 :
    _intrVecEnable_0_T_7; // @[src/main/scala/nutcore/backend/fu/CSR.scala 601:51]
  wire  intrVecEnable_4 = ideleg[4] ? priviledgeMode == 2'h1 & mstatusStruct_ie_s | priviledgeMode < 2'h1 :
    _intrVecEnable_0_T_7; // @[src/main/scala/nutcore/backend/fu/CSR.scala 601:51]
  wire  intrVecEnable_5 = ideleg[5] ? priviledgeMode == 2'h1 & mstatusStruct_ie_s | priviledgeMode < 2'h1 :
    _intrVecEnable_0_T_7; // @[src/main/scala/nutcore/backend/fu/CSR.scala 601:51]
  wire  intrVecEnable_6 = ideleg[6] ? priviledgeMode == 2'h1 & mstatusStruct_ie_s | priviledgeMode < 2'h1 :
    _intrVecEnable_0_T_7; // @[src/main/scala/nutcore/backend/fu/CSR.scala 601:51]
  wire  intrVecEnable_7 = ideleg[7] ? priviledgeMode == 2'h1 & mstatusStruct_ie_s | priviledgeMode < 2'h1 :
    _intrVecEnable_0_T_7; // @[src/main/scala/nutcore/backend/fu/CSR.scala 601:51]
  wire  intrVecEnable_8 = ideleg[8] ? priviledgeMode == 2'h1 & mstatusStruct_ie_s | priviledgeMode < 2'h1 :
    _intrVecEnable_0_T_7; // @[src/main/scala/nutcore/backend/fu/CSR.scala 601:51]
  wire  intrVecEnable_9 = ideleg[9] ? priviledgeMode == 2'h1 & mstatusStruct_ie_s | priviledgeMode < 2'h1 :
    _intrVecEnable_0_T_7; // @[src/main/scala/nutcore/backend/fu/CSR.scala 601:51]
  wire  intrVecEnable_10 = ideleg[10] ? priviledgeMode == 2'h1 & mstatusStruct_ie_s | priviledgeMode < 2'h1 :
    _intrVecEnable_0_T_7; // @[src/main/scala/nutcore/backend/fu/CSR.scala 601:51]
  wire  intrVecEnable_11 = ideleg[11] ? priviledgeMode == 2'h1 & mstatusStruct_ie_s | priviledgeMode < 2'h1 :
    _intrVecEnable_0_T_7; // @[src/main/scala/nutcore/backend/fu/CSR.scala 601:51]
  wire [11:0] _intrVec_T_2 = mie[11:0] & _ideleg_T; // @[src/main/scala/nutcore/backend/fu/CSR.scala 606:27]
  wire [5:0] intrVec_lo_1 = {intrVecEnable_5,intrVecEnable_4,intrVecEnable_3,intrVecEnable_2,intrVecEnable_1,
    intrVecEnable_0}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 606:65]
  wire [11:0] _intrVec_T_3 = {intrVecEnable_11,intrVecEnable_10,intrVecEnable_9,intrVecEnable_8,intrVecEnable_7,
    intrVecEnable_6,intrVec_lo_1}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 606:65]
  wire [11:0] intrVec = _intrVec_T_2 & _intrVec_T_3; // @[src/main/scala/nutcore/backend/fu/CSR.scala 606:49]
  wire [2:0] _intrNO_T = io_cfIn_intrVec_4 ? 3'h4 : 3'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 610:69]
  wire [3:0] _intrNO_T_1 = io_cfIn_intrVec_8 ? 4'h8 : {{1'd0}, _intrNO_T}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 610:69]
  wire [3:0] _intrNO_T_2 = io_cfIn_intrVec_0 ? 4'h0 : _intrNO_T_1; // @[src/main/scala/nutcore/backend/fu/CSR.scala 610:69]
  wire [3:0] _intrNO_T_3 = io_cfIn_intrVec_5 ? 4'h5 : _intrNO_T_2; // @[src/main/scala/nutcore/backend/fu/CSR.scala 610:69]
  wire [3:0] _intrNO_T_4 = io_cfIn_intrVec_9 ? 4'h9 : _intrNO_T_3; // @[src/main/scala/nutcore/backend/fu/CSR.scala 610:69]
  wire [3:0] _intrNO_T_5 = io_cfIn_intrVec_1 ? 4'h1 : _intrNO_T_4; // @[src/main/scala/nutcore/backend/fu/CSR.scala 610:69]
  wire [3:0] _intrNO_T_6 = io_cfIn_intrVec_7 ? 4'h7 : _intrNO_T_5; // @[src/main/scala/nutcore/backend/fu/CSR.scala 610:69]
  wire [3:0] _intrNO_T_7 = io_cfIn_intrVec_11 ? 4'hb : _intrNO_T_6; // @[src/main/scala/nutcore/backend/fu/CSR.scala 610:69]
  wire [3:0] intrNO = io_cfIn_intrVec_3 ? 4'h3 : _intrNO_T_7; // @[src/main/scala/nutcore/backend/fu/CSR.scala 610:69]
  wire [5:0] raiseIntr_lo = {io_cfIn_intrVec_5,io_cfIn_intrVec_4,io_cfIn_intrVec_3,io_cfIn_intrVec_2,io_cfIn_intrVec_1,
    io_cfIn_intrVec_0}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 612:35]
  wire [11:0] _raiseIntr_T = {io_cfIn_intrVec_11,io_cfIn_intrVec_10,io_cfIn_intrVec_9,io_cfIn_intrVec_8,
    io_cfIn_intrVec_7,io_cfIn_intrVec_6,raiseIntr_lo}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 612:35]
  wire  raiseIntr = |_raiseIntr_T; // @[src/main/scala/nutcore/backend/fu/CSR.scala 612:42]
  wire  csrExceptionVec_3 = io_in_valid & isEbreak; // @[src/main/scala/nutcore/backend/fu/CSR.scala 619:46]
  wire  csrExceptionVec_11 = _T_1025 & io_in_valid & isEcall; // @[src/main/scala/nutcore/backend/fu/CSR.scala 620:70]
  wire  csrExceptionVec_9 = _intrVecEnable_0_T & io_in_valid & isEcall; // @[src/main/scala/nutcore/backend/fu/CSR.scala 621:70]
  wire  csrExceptionVec_8 = priviledgeMode == 2'h0 & io_in_valid & isEcall; // @[src/main/scala/nutcore/backend/fu/CSR.scala 622:70]
  wire  csrExceptionVec_2 = (isIllegalAddr | isIllegalAccess) & wen; // @[src/main/scala/nutcore/backend/fu/CSR.scala 623:71]
  wire [7:0] raiseExceptionVec_lo = {4'h0,csrExceptionVec_3,csrExceptionVec_2,2'h0}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 627:43]
  wire [15:0] _raiseExceptionVec_T = {io_dmemMMU_storePF,1'h0,io_dmemMMU_loadPF,1'h0,csrExceptionVec_11,1'h0,
    csrExceptionVec_9,csrExceptionVec_8,raiseExceptionVec_lo}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 627:43]
  wire [7:0] raiseExceptionVec_lo_1 = {1'h0,io_cfIn_exceptionVec_6,1'h0,io_cfIn_exceptionVec_4,1'h0,
    io_cfIn_exceptionVec_2,io_cfIn_exceptionVec_1,1'h0}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 627:68]
  wire [15:0] _raiseExceptionVec_T_1 = {2'h0,1'h0,io_cfIn_exceptionVec_12,4'h0,raiseExceptionVec_lo_1}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 627:68]
  wire [15:0] raiseExceptionVec = _raiseExceptionVec_T | _raiseExceptionVec_T_1; // @[src/main/scala/nutcore/backend/fu/CSR.scala 627:50]
  wire  raiseException = |raiseExceptionVec; // @[src/main/scala/nutcore/backend/fu/CSR.scala 628:42]
  wire [2:0] _exceptionNO_T_1 = raiseExceptionVec[5] ? 3'h5 : 3'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 629:74]
  wire [2:0] _exceptionNO_T_3 = raiseExceptionVec[7] ? 3'h7 : _exceptionNO_T_1; // @[src/main/scala/nutcore/backend/fu/CSR.scala 629:74]
  wire [3:0] _exceptionNO_T_5 = raiseExceptionVec[13] ? 4'hd : {{1'd0}, _exceptionNO_T_3}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 629:74]
  wire [3:0] _exceptionNO_T_7 = raiseExceptionVec[15] ? 4'hf : _exceptionNO_T_5; // @[src/main/scala/nutcore/backend/fu/CSR.scala 629:74]
  wire [3:0] _exceptionNO_T_9 = raiseExceptionVec[4] ? 4'h4 : _exceptionNO_T_7; // @[src/main/scala/nutcore/backend/fu/CSR.scala 629:74]
  wire [3:0] _exceptionNO_T_11 = raiseExceptionVec[6] ? 4'h6 : _exceptionNO_T_9; // @[src/main/scala/nutcore/backend/fu/CSR.scala 629:74]
  wire [3:0] _exceptionNO_T_13 = raiseExceptionVec[8] ? 4'h8 : _exceptionNO_T_11; // @[src/main/scala/nutcore/backend/fu/CSR.scala 629:74]
  wire [3:0] _exceptionNO_T_15 = raiseExceptionVec[9] ? 4'h9 : _exceptionNO_T_13; // @[src/main/scala/nutcore/backend/fu/CSR.scala 629:74]
  wire [3:0] _exceptionNO_T_17 = raiseExceptionVec[11] ? 4'hb : _exceptionNO_T_15; // @[src/main/scala/nutcore/backend/fu/CSR.scala 629:74]
  wire [3:0] _exceptionNO_T_19 = raiseExceptionVec[0] ? 4'h0 : _exceptionNO_T_17; // @[src/main/scala/nutcore/backend/fu/CSR.scala 629:74]
  wire [3:0] _exceptionNO_T_21 = raiseExceptionVec[2] ? 4'h2 : _exceptionNO_T_19; // @[src/main/scala/nutcore/backend/fu/CSR.scala 629:74]
  wire [3:0] _exceptionNO_T_23 = raiseExceptionVec[1] ? 4'h1 : _exceptionNO_T_21; // @[src/main/scala/nutcore/backend/fu/CSR.scala 629:74]
  wire [3:0] _exceptionNO_T_25 = raiseExceptionVec[12] ? 4'hc : _exceptionNO_T_23; // @[src/main/scala/nutcore/backend/fu/CSR.scala 629:74]
  wire [3:0] exceptionNO = raiseExceptionVec[3] ? 4'h3 : _exceptionNO_T_25; // @[src/main/scala/nutcore/backend/fu/CSR.scala 629:74]
  wire [63:0] _causeNO_T = {raiseIntr, 63'h0}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 632:28]
  wire [3:0] _causeNO_T_1 = raiseIntr ? intrNO : exceptionNO; // @[src/main/scala/nutcore/backend/fu/CSR.scala 632:46]
  wire [63:0] _GEN_334 = {{60'd0}, _causeNO_T_1}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 632:41]
  wire [63:0] causeNO = _causeNO_T | _GEN_334; // @[src/main/scala/nutcore/backend/fu/CSR.scala 632:41]
  wire  raiseExceptionIntr = (raiseException | raiseIntr) & io_instrValid; // @[src/main/scala/nutcore/backend/fu/CSR.scala 635:58]
  wire [38:0] _io_redirect_target_T_1 = io_cfIn_pc + 39'h4; // @[src/main/scala/nutcore/backend/fu/CSR.scala 640:51]
  wire [63:0] deleg = raiseIntr ? mideleg : medeleg; // @[src/main/scala/nutcore/backend/fu/CSR.scala 650:18]
  wire [63:0] _delegS_T_1 = deleg >> causeNO[3:0]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 652:22]
  wire  delegS = _delegS_T_1[0] & _intrVecEnable_0_T_6; // @[src/main/scala/nutcore/backend/fu/CSR.scala 652:38]
  wire [63:0] _trapTarget_T = delegS ? stvec : mtvec; // @[src/main/scala/nutcore/backend/fu/CSR.scala 656:20]
  wire [38:0] trapTarget = _trapTarget_T[38:0]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 656:42]
  wire [38:0] _GEN_172 = io_in_valid & isSret ? sepc[38:0] : mepc[38:0]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 674:26 684:15]
  wire [38:0] retTarget = io_in_valid & isUret ? 39'h0 : _GEN_172; // @[src/main/scala/nutcore/backend/fu/CSR.scala 687:26 695:15]
  wire [38:0] _io_redirect_target_T_2 = raiseExceptionIntr ? trapTarget : retTarget; // @[src/main/scala/nutcore/backend/fu/CSR.scala 640:61]
  reg [63:0] c_7; // @[src/main/scala/utils/GTimer.scala 24:20]
  wire [63:0] _c_T_15 = c_7 + 64'h1; // @[src/main/scala/utils/GTimer.scala 25:12]
  wire  _T_1109 = raiseExceptionIntr & DISPLAY_ENABLE; // @[src/main/scala/utils/Debug.scala 55:16]
  reg [63:0] c_8; // @[src/main/scala/utils/GTimer.scala 24:20]
  wire [63:0] _c_T_17 = c_8 + 64'h1; // @[src/main/scala/utils/GTimer.scala 25:12]
  reg [63:0] c_9; // @[src/main/scala/utils/GTimer.scala 24:20]
  wire [63:0] _c_T_19 = c_9 + 64'h1; // @[src/main/scala/utils/GTimer.scala 25:12]
  reg [63:0] c_10; // @[src/main/scala/utils/GTimer.scala 24:20]
  wire [63:0] _c_T_21 = c_10 + 64'h1; // @[src/main/scala/utils/GTimer.scala 25:12]
  reg [63:0] c_11; // @[src/main/scala/utils/GTimer.scala 24:20]
  wire [63:0] _c_T_23 = c_11 + 64'h1; // @[src/main/scala/utils/GTimer.scala 25:12]
  wire  _T_1125 = io_redirect_valid & DISPLAY_ENABLE; // @[src/main/scala/utils/Debug.scala 55:16]
  reg [63:0] c_12; // @[src/main/scala/utils/GTimer.scala 24:20]
  wire [63:0] _c_T_25 = c_12 + 64'h1; // @[src/main/scala/utils/GTimer.scala 25:12]
  wire  _T_1130 = resetSatp & DISPLAY_ENABLE; // @[src/main/scala/utils/Debug.scala 55:16]
  wire  tvalWen = ~(_T_1024 | io_cfIn_exceptionVec_4 | io_cfIn_exceptionVec_6) | raiseIntr; // @[src/main/scala/nutcore/backend/fu/CSR.scala 653:130]
  wire [5:0] mstatus_lo_lo = {mstatusStruct_pie_s,mstatusStruct_pie_u,mstatusStruct_pie_m,mstatusStruct_ie_h,
    mstatusStruct_ie_s,mstatusStruct_ie_u}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 669:27]
  wire [14:0] mstatus_lo = {mstatusStruct_fs,2'h0,mstatusStruct_hpp,mstatusStruct_spp,1'h1,mstatusStruct_pie_h,
    mstatus_lo_lo}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 669:27]
  wire [6:0] mstatus_hi_lo = {mstatusStruct_tw,mstatusStruct_tvm,mstatusStruct_mxr,mstatusStruct_sum,mstatusStruct_mprv,
    mstatusStruct_xs}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 669:27]
  wire [63:0] _mstatus_T_8 = {mstatusStruct_sd,mstatusStruct_pad1,mstatusStruct_sxl,mstatusStruct_uxl,mstatusStruct_pad0
    ,mstatusStruct_tsr,mstatus_hi_lo,mstatus_lo}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 669:27]
  wire [1:0] _GEN_165 = io_in_valid & isMret ? mstatusStruct_mpp : priviledgeMode; // @[src/main/scala/nutcore/backend/fu/CSR.scala 661:26 666:20 369:31]
  wire [63:0] _GEN_166 = io_in_valid & isMret ? _mstatus_T_8 : _GEN_97; // @[src/main/scala/nutcore/backend/fu/CSR.scala 661:26 669:13]
  wire [1:0] _priviledgeMode_T = {1'h0,mstatusStruct_spp}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 679:26]
  wire [5:0] mstatus_lo_lo_1 = {1'h1,mstatusStruct_pie_u,mstatusStruct_ie_m,mstatusStruct_ie_h,mstatusStruct_pie_s,
    mstatusStruct_ie_u}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 682:27]
  wire [14:0] mstatus_lo_1 = {mstatusStruct_fs,mstatusStruct_mpp,mstatusStruct_hpp,1'h0,mstatusStruct_pie_m,
    mstatusStruct_pie_h,mstatus_lo_lo_1}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 682:27]
  wire [63:0] _mstatus_T_9 = {mstatusStruct_sd,mstatusStruct_pad1,mstatusStruct_sxl,mstatusStruct_uxl,mstatusStruct_pad0
    ,mstatusStruct_tsr,mstatus_hi_lo,mstatus_lo_1}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 682:27]
  wire [5:0] mstatus_lo_lo_2 = {mstatusStruct_pie_s,1'h1,mstatusStruct_ie_m,mstatusStruct_ie_h,mstatusStruct_ie_s,
    mstatusStruct_pie_u}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 694:27]
  wire [14:0] mstatus_lo_2 = {mstatusStruct_fs,mstatusStruct_mpp,mstatusStruct_hpp,mstatusStruct_spp,mstatusStruct_pie_m
    ,mstatusStruct_pie_h,mstatus_lo_lo_2}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 694:27]
  wire [63:0] _mstatus_T_10 = {mstatusStruct_sd,mstatusStruct_pad1,mstatusStruct_sxl,mstatusStruct_uxl,
    mstatusStruct_pad0,mstatusStruct_tsr,mstatus_hi_lo,mstatus_lo_2}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 694:27]
  wire [1:0] _GEN_180 = delegS ? priviledgeMode : {{1'd0}, mstatusStruct_spp}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 702:19 705:22 700:30]
  wire  mstatusNew_3_pie_s = delegS ? mstatusStruct_ie_s : mstatusStruct_pie_s; // @[src/main/scala/nutcore/backend/fu/CSR.scala 702:19 706:24 700:30]
  wire  mstatusNew_3_ie_s = delegS ? 1'h0 : mstatusStruct_ie_s; // @[src/main/scala/nutcore/backend/fu/CSR.scala 702:19 707:23 700:30]
  wire [1:0] mstatusNew_3_mpp = delegS ? mstatusStruct_mpp : priviledgeMode; // @[src/main/scala/nutcore/backend/fu/CSR.scala 702:19 700:30 715:22]
  wire  mstatusNew_3_pie_m = delegS ? mstatusStruct_pie_m : mstatusStruct_ie_m; // @[src/main/scala/nutcore/backend/fu/CSR.scala 702:19 700:30 716:24]
  wire  mstatusNew_3_ie_m = delegS & mstatusStruct_ie_m; // @[src/main/scala/nutcore/backend/fu/CSR.scala 702:19 700:30 717:23]
  wire [5:0] mstatus_lo_lo_3 = {mstatusNew_3_pie_s,mstatusStruct_pie_u,mstatusNew_3_ie_m,mstatusStruct_ie_h,
    mstatusNew_3_ie_s,mstatusStruct_ie_u}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 729:27]
  wire  mstatusNew_3_spp = _GEN_180[0]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 700:30]
  wire [14:0] mstatus_lo_3 = {mstatusStruct_fs,mstatusNew_3_mpp,mstatusStruct_hpp,mstatusNew_3_spp,mstatusNew_3_pie_m,
    mstatusStruct_pie_h,mstatus_lo_lo_3}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 729:27]
  wire [63:0] _mstatus_T_11 = {mstatusStruct_sd,mstatusStruct_pad1,mstatusStruct_sxl,mstatusStruct_uxl,
    mstatusStruct_pad0,mstatusStruct_tsr,mstatus_hi_lo,mstatus_lo_3}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 729:27]
  wire [63:0] _perfCnts_0_T_5 = perfCnts_0 + 64'h1; // @[src/main/scala/nutcore/backend/fu/CSR.scala 838:71]
  wire  _WIRE_1 = 1'h1; // @[src/main/scala/nutcore/backend/fu/CSR.scala 855:{33,33}]
  wire [63:0] _perfCnts_2_T_5 = perfCnts_2 + 64'h1; // @[src/main/scala/nutcore/backend/fu/CSR.scala 838:71]
  wire [63:0] _perfCnts_3_T_5 = perfCnts_3 + 64'h1; // @[src/main/scala/nutcore/backend/fu/CSR.scala 838:71]
  wire [63:0] _perfCnts_4_T_5 = perfCnts_4 + 64'h1; // @[src/main/scala/nutcore/backend/fu/CSR.scala 838:71]
  wire [63:0] _perfCnts_5_T_5 = perfCnts_5 + 64'h1; // @[src/main/scala/nutcore/backend/fu/CSR.scala 838:71]
  wire [63:0] _perfCnts_6_T_5 = perfCnts_6 + 64'h1; // @[src/main/scala/nutcore/backend/fu/CSR.scala 838:71]
  wire [63:0] _perfCnts_7_T_5 = perfCnts_7 + 64'h1; // @[src/main/scala/nutcore/backend/fu/CSR.scala 838:71]
  wire [63:0] _perfCnts_8_T_5 = perfCnts_8 + 64'h1; // @[src/main/scala/nutcore/backend/fu/CSR.scala 838:71]
  wire [63:0] _perfCnts_9_T_5 = perfCnts_9 + 64'h1; // @[src/main/scala/nutcore/backend/fu/CSR.scala 838:71]
  wire [63:0] _perfCnts_10_T_5 = perfCnts_10 + 64'h1; // @[src/main/scala/nutcore/backend/fu/CSR.scala 838:71]
  wire [63:0] _perfCnts_11_T_5 = perfCnts_11 + 64'h1; // @[src/main/scala/nutcore/backend/fu/CSR.scala 838:71]
  wire [63:0] _perfCnts_14_T_5 = perfCnts_14 + 64'h1; // @[src/main/scala/nutcore/backend/fu/CSR.scala 838:71]
  wire [63:0] _perfCnts_15_T_5 = perfCnts_15 + 64'h1; // @[src/main/scala/nutcore/backend/fu/CSR.scala 838:71]
  wire [63:0] _perfCnts_16_T_5 = perfCnts_16 + 64'h1; // @[src/main/scala/nutcore/backend/fu/CSR.scala 838:71]
  wire [63:0] _perfCnts_17_T_5 = perfCnts_17 + 64'h1; // @[src/main/scala/nutcore/backend/fu/CSR.scala 838:71]
  wire [63:0] _perfCnts_18_T_5 = perfCnts_18 + 64'h1; // @[src/main/scala/nutcore/backend/fu/CSR.scala 838:71]
  wire [63:0] _perfCnts_19_T_5 = perfCnts_19 + 64'h1; // @[src/main/scala/nutcore/backend/fu/CSR.scala 838:71]
  wire [63:0] _perfCnts_20_T_5 = perfCnts_20 + 64'h1; // @[src/main/scala/nutcore/backend/fu/CSR.scala 838:71]
  wire [63:0] _perfCnts_21_T_5 = perfCnts_21 + 64'h1; // @[src/main/scala/nutcore/backend/fu/CSR.scala 838:71]
  wire [63:0] _perfCnts_22_T_5 = perfCnts_22 + 64'h1; // @[src/main/scala/nutcore/backend/fu/CSR.scala 838:71]
  wire [63:0] _perfCnts_23_T_5 = perfCnts_23 + 64'h1; // @[src/main/scala/nutcore/backend/fu/CSR.scala 838:71]
  wire [63:0] _perfCnts_25_T_5 = perfCnts_25 + 64'h1; // @[src/main/scala/nutcore/backend/fu/CSR.scala 838:71]
  wire [63:0] _perfCnts_26_T_5 = perfCnts_26 + 64'h1; // @[src/main/scala/nutcore/backend/fu/CSR.scala 838:71]
  wire [63:0] _perfCnts_27_T_5 = perfCnts_27 + 64'h1; // @[src/main/scala/nutcore/backend/fu/CSR.scala 838:71]
  wire [63:0] _perfCnts_28_T_5 = perfCnts_28 + 64'h1; // @[src/main/scala/nutcore/backend/fu/CSR.scala 838:71]
  wire [63:0] _perfCnts_29_T_5 = perfCnts_29 + 64'h1; // @[src/main/scala/nutcore/backend/fu/CSR.scala 838:71]
  wire [63:0] _perfCnts_30_T_5 = perfCnts_30 + 64'h1; // @[src/main/scala/nutcore/backend/fu/CSR.scala 838:71]
  wire [63:0] _perfCnts_31_T_5 = perfCnts_31 + 64'h1; // @[src/main/scala/nutcore/backend/fu/CSR.scala 838:71]
  wire [63:0] _perfCnts_32_T_5 = perfCnts_32 + 64'h1; // @[src/main/scala/nutcore/backend/fu/CSR.scala 838:71]
  wire [63:0] _perfCnts_49_T_5 = perfCnts_49 + 64'h1; // @[src/main/scala/nutcore/backend/fu/CSR.scala 838:71]
  wire [63:0] _perfCnts_50_T_5 = perfCnts_50 + 64'h1; // @[src/main/scala/nutcore/backend/fu/CSR.scala 838:71]
  wire [63:0] _perfCnts_51_T_5 = perfCnts_51 + 64'h1; // @[src/main/scala/nutcore/backend/fu/CSR.scala 838:71]
  wire [63:0] _perfCnts_52_T_5 = perfCnts_52 + 64'h1; // @[src/main/scala/nutcore/backend/fu/CSR.scala 838:71]
  wire [63:0] _perfCnts_53_T_5 = perfCnts_53 + 64'h1; // @[src/main/scala/nutcore/backend/fu/CSR.scala 838:71]
  wire [63:0] _perfCnts_2_T_7 = perfCnts_2 + 64'h2; // @[src/main/scala/nutcore/backend/fu/CSR.scala 848:86]
  wire [64:0] _perfCnts_99_T_6 = {{1'd0}, perfCnts_99}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 850:69]
  wire [64:0] _perfCnts_100_T_6 = {{1'd0}, perfCnts_100}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 851:69]
  wire [64:0] _perfCnts_101_T_6 = {{1'd0}, perfCnts_102}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 852:69]
  wire [11:0] _WIRE = intrVec; // @[src/main/scala/nutcore/backend/fu/CSR.scala 606:49]
  wire  _GEN_335 = _T_1024 & DISPLAY_ENABLE; // @[src/main/scala/utils/Debug.scala 56:24]
  wire  _GEN_337 = _T_1034 & DISPLAY_ENABLE; // @[src/main/scala/utils/Debug.scala 56:24]
  assign io_out_valid = io_in_valid; // @[src/main/scala/nutcore/backend/fu/CSR.scala 733:16]
  assign io_out_bits = _rdata_T_645 | _rdata_T_485; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign io_redirect_target = resetSatp ? _io_redirect_target_T_1 : _io_redirect_target_T_2; // @[src/main/scala/nutcore/backend/fu/CSR.scala 640:28]
  assign io_redirect_valid = io_in_valid & _isEbreak_T_1 | raiseExceptionIntr | resetSatp; // @[src/main/scala/nutcore/backend/fu/CSR.scala 638:80]
  assign io_intrNO = raiseIntr ? causeNO : 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 633:19]
  assign io_imemMMU_priviledgeMode = priviledgeMode; // @[src/main/scala/nutcore/backend/fu/CSR.scala 529:29]
  assign io_dmemMMU_priviledgeMode = mstatusStruct_mprv ? mstatusStruct_mpp : priviledgeMode; // @[src/main/scala/nutcore/backend/fu/CSR.scala 530:35]
  assign io_dmemMMU_status_sum = mstatus[18]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 299:39]
  assign io_dmemMMU_status_mxr = mstatus[19]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 299:39]
  assign io_wenFix = |raiseExceptionVec; // @[src/main/scala/nutcore/backend/fu/CSR.scala 628:42]
  assign lr_0 = lr;
  assign lrAddr_0 = lrAddr;
  assign satp_0 = satp;
  assign _WIRE_4 = _WIRE;
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 252:22]
      mtvec <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 252:22]
    end else if (_T_693 & addr == 12'h305) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      mtvec <= wdata; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 253:27]
      mcounteren <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 253:27]
    end else if (_T_693 & addr == 12'h306) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      mcounteren <= wdata; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 254:23]
      mcause <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 254:23]
    end else if (raiseExceptionIntr) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 698:29]
      if (delegS) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 702:19]
        mcause <= _GEN_34;
      end else begin
        mcause <= causeNO; // @[src/main/scala/nutcore/backend/fu/CSR.scala 713:14]
      end
    end else begin
      mcause <= _GEN_34;
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 255:22]
      mtval <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 255:22]
    end else if (raiseExceptionIntr) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 698:29]
      if (delegS) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 702:19]
        mtval <= _GEN_164;
      end else if (tvalWen) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 719:20]
        mtval <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 719:27]
      end else begin
        mtval <= _GEN_164;
      end
    end else begin
      mtval <= _GEN_164;
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 256:21]
      mepc <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 256:21]
    end else if (raiseExceptionIntr) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 698:29]
      if (delegS) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 702:19]
        mepc <= _GEN_143;
      end else begin
        mepc <= _tval_T_9; // @[src/main/scala/nutcore/backend/fu/CSR.scala 714:12]
      end
    end else begin
      mepc <= _GEN_143;
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 258:20]
      mie <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 258:20]
    end else if (_T_693 & addr == 12'h304) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      mie <= wdata; // @[src/main/scala/utils/RegMap.scala 50:76]
    end else if (_T_693 & addr == 12'h104) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      mie <= _mie_T_3; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 260:24]
      mipReg <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 260:24]
    end else if (_T_693 & addr == 12'h144) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      mipReg <= _mipReg_T_7; // @[src/main/scala/utils/RegMap.scala 50:76]
    end else if (_T_693 & addr == 12'h344) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      mipReg <= _mipReg_T_3; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 270:21]
      misa <= 64'h8000000000141105; // @[src/main/scala/nutcore/backend/fu/CSR.scala 270:21]
    end else if (_T_693 & addr == 12'h301) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      misa <= wdata; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 278:24]
      mstatus <= 64'ha00001800; // @[src/main/scala/nutcore/backend/fu/CSR.scala 278:24]
    end else if (raiseExceptionIntr) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 698:29]
      mstatus <= _mstatus_T_11; // @[src/main/scala/nutcore/backend/fu/CSR.scala 729:13]
    end else if (io_in_valid & isUret) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 687:26]
      mstatus <= _mstatus_T_10; // @[src/main/scala/nutcore/backend/fu/CSR.scala 694:13]
    end else if (io_in_valid & isSret) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 674:26]
      mstatus <= _mstatus_T_9; // @[src/main/scala/nutcore/backend/fu/CSR.scala 682:13]
    end else begin
      mstatus <= _GEN_166;
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 306:24]
      medeleg <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 306:24]
    end else if (_T_693 & addr == 12'h302) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      medeleg <= _medeleg_T_3; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 307:24]
      mideleg <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 307:24]
    end else if (_T_693 & addr == 12'h303) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      mideleg <= _mideleg_T_3; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 308:25]
      mscratch <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 308:25]
    end else if (_T_693 & addr == 12'h340) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      mscratch <= wdata; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 310:24]
      pmpcfg0 <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 310:24]
    end else if (_T_693 & addr == 12'h3a0) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      pmpcfg0 <= wdata; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 311:24]
      pmpcfg1 <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 311:24]
    end else if (_T_693 & addr == 12'h3a1) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      pmpcfg1 <= wdata; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 312:24]
      pmpcfg2 <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 312:24]
    end else if (_T_693 & addr == 12'h3a2) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      pmpcfg2 <= wdata; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 313:24]
      pmpcfg3 <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 313:24]
    end else if (_T_693 & addr == 12'h3a3) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      pmpcfg3 <= wdata; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 314:25]
      pmpaddr0 <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 314:25]
    end else if (_T_693 & addr == 12'h3b0) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      pmpaddr0 <= _pmpaddr0_T_3; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 315:25]
      pmpaddr1 <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 315:25]
    end else if (_T_693 & addr == 12'h3b1) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      pmpaddr1 <= _pmpaddr1_T_3; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 316:25]
      pmpaddr2 <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 316:25]
    end else if (_T_693 & addr == 12'h3b2) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      pmpaddr2 <= _pmpaddr2_T_3; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 317:25]
      pmpaddr3 <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 317:25]
    end else if (_T_693 & addr == 12'h3b3) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      pmpaddr3 <= _pmpaddr3_T_3; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 332:22]
      stvec <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 332:22]
    end else if (_T_693 & addr == 12'h105) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      stvec <= wdata; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 337:21]
      satp <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 337:21]
    end else if (_T_693 & addr == 12'h180) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      satp <= wdata; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 338:21]
      sepc <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 338:21]
    end else if (raiseExceptionIntr) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 698:29]
      if (delegS) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 702:19]
        sepc <= _tval_T_9; // @[src/main/scala/nutcore/backend/fu/CSR.scala 704:12]
      end else begin
        sepc <= _GEN_32;
      end
    end else begin
      sepc <= _GEN_32;
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 339:23]
      scause <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 339:23]
    end else if (raiseExceptionIntr) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 698:29]
      if (delegS) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 702:19]
        scause <= causeNO; // @[src/main/scala/nutcore/backend/fu/CSR.scala 703:14]
      end else begin
        scause <= _GEN_151;
      end
    end else begin
      scause <= _GEN_151;
    end
    if (raiseExceptionIntr) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 698:29]
      if (delegS) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 702:19]
        if (tvalWen) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 709:20]
          stval <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 709:27]
        end else begin
          stval <= _GEN_163;
        end
      end else begin
        stval <= _GEN_163;
      end
    end else begin
      stval <= _GEN_163;
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 341:25]
      sscratch <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 341:25]
    end else if (_T_693 & addr == 12'h140) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      sscratch <= wdata; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 342:27]
      scounteren <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 342:27]
    end else if (_T_693 & addr == 12'h106) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      scounteren <= wdata; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 355:19]
      lr <= 1'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 355:19]
    end else if (io_in_valid & isSret) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 674:26]
      lr <= 1'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 683:8]
    end else if (io_in_valid & isMret) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 661:26]
      lr <= 1'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 670:8]
    end else if (set_lr) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 363:14]
      lr <= set_lr_val; // @[src/main/scala/nutcore/backend/fu/CSR.scala 364:8]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 356:23]
      lrAddr <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 356:23]
    end else if (set_lr) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 363:14]
      lrAddr <= set_lr_addr; // @[src/main/scala/nutcore/backend/fu/CSR.scala 365:12]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 369:31]
      priviledgeMode <= 2'h3; // @[src/main/scala/nutcore/backend/fu/CSR.scala 369:31]
    end else if (raiseExceptionIntr) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 698:29]
      if (delegS) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 702:19]
        priviledgeMode <= 2'h1; // @[src/main/scala/nutcore/backend/fu/CSR.scala 708:22]
      end else begin
        priviledgeMode <= 2'h3; // @[src/main/scala/nutcore/backend/fu/CSR.scala 718:22]
      end
    end else if (io_in_valid & isUret) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 687:26]
      priviledgeMode <= 2'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 692:20]
    end else if (io_in_valid & isSret) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 674:26]
      priviledgeMode <= _priviledgeMode_T; // @[src/main/scala/nutcore/backend/fu/CSR.scala 679:20]
    end else begin
      priviledgeMode <= _GEN_165;
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
      perfCnts_0 <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
    end else begin
      perfCnts_0 <= _perfCnts_0_T_5;
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
      perfCnts_1 <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
    end else if (_T_693 & addr == 12'hb01) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      perfCnts_1 <= wdata; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
      perfCnts_2 <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
    end else if (perfCntCondMultiCommit) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 848:35]
      perfCnts_2 <= _perfCnts_2_T_7; // @[src/main/scala/nutcore/backend/fu/CSR.scala 848:60]
    end else if (perfCntCondMinstret) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 838:62]
      perfCnts_2 <= _perfCnts_2_T_5; // @[src/main/scala/nutcore/backend/fu/CSR.scala 838:66]
    end else if (_T_693 & addr == 12'hb02) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      perfCnts_2 <= wdata; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
      perfCnts_3 <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
    end else if (perfCntCondMultiCommit) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 838:62]
      perfCnts_3 <= _perfCnts_3_T_5; // @[src/main/scala/nutcore/backend/fu/CSR.scala 838:66]
    end else if (_T_693 & addr == 12'hb03) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      perfCnts_3 <= wdata; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
      perfCnts_4 <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
    end else if (perfCntCondMimemStall) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 838:62]
      perfCnts_4 <= _perfCnts_4_T_5; // @[src/main/scala/nutcore/backend/fu/CSR.scala 838:66]
    end else if (_T_693 & addr == 12'hb04) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      perfCnts_4 <= wdata; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
      perfCnts_5 <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
    end else if (perfCntCondMaluInstr) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 838:62]
      perfCnts_5 <= _perfCnts_5_T_5; // @[src/main/scala/nutcore/backend/fu/CSR.scala 838:66]
    end else if (_T_693 & addr == 12'hb05) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      perfCnts_5 <= wdata; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
      perfCnts_6 <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
    end else if (perfCntCondMbruInstr) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 838:62]
      perfCnts_6 <= _perfCnts_6_T_5; // @[src/main/scala/nutcore/backend/fu/CSR.scala 838:66]
    end else if (_T_693 & addr == 12'hb06) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      perfCnts_6 <= wdata; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
      perfCnts_7 <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
    end else if (perfCntCondMlsuInstr) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 838:62]
      perfCnts_7 <= _perfCnts_7_T_5; // @[src/main/scala/nutcore/backend/fu/CSR.scala 838:66]
    end else if (_T_693 & addr == 12'hb07) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      perfCnts_7 <= wdata; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
      perfCnts_8 <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
    end else if (perfCntCondMmduInstr) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 838:62]
      perfCnts_8 <= _perfCnts_8_T_5; // @[src/main/scala/nutcore/backend/fu/CSR.scala 838:66]
    end else if (_T_693 & addr == 12'hb08) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      perfCnts_8 <= wdata; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
      perfCnts_9 <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
    end else if (perfCntCondMcsrInstr) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 838:62]
      perfCnts_9 <= _perfCnts_9_T_5; // @[src/main/scala/nutcore/backend/fu/CSR.scala 838:66]
    end else if (_T_693 & addr == 12'hb09) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      perfCnts_9 <= wdata; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
      perfCnts_10 <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
    end else if (perfCntCondMloadInstr) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 838:62]
      perfCnts_10 <= _perfCnts_10_T_5; // @[src/main/scala/nutcore/backend/fu/CSR.scala 838:66]
    end else if (_T_693 & addr == 12'hb0a) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      perfCnts_10 <= wdata; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
      perfCnts_11 <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
    end else if (perfCntCondMmmioInstr) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 838:62]
      perfCnts_11 <= _perfCnts_11_T_5; // @[src/main/scala/nutcore/backend/fu/CSR.scala 838:66]
    end else if (_T_693 & addr == 12'hb0b) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      perfCnts_11 <= wdata; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
      perfCnts_12 <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
    end else if (_T_693 & addr == 12'hb0c) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      perfCnts_12 <= wdata; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
      perfCnts_13 <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
    end else if (_T_693 & addr == 12'hb0d) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      perfCnts_13 <= wdata; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
      perfCnts_14 <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
    end else if (perfCntCondMmulInstr) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 838:62]
      perfCnts_14 <= _perfCnts_14_T_5; // @[src/main/scala/nutcore/backend/fu/CSR.scala 838:66]
    end else if (_T_693 & addr == 12'hb0e) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      perfCnts_14 <= wdata; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
      perfCnts_15 <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
    end else if (perfCntCondMifuFlush) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 838:62]
      perfCnts_15 <= _perfCnts_15_T_5; // @[src/main/scala/nutcore/backend/fu/CSR.scala 838:66]
    end else if (_T_693 & addr == 12'hb0f) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      perfCnts_15 <= wdata; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
      perfCnts_16 <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
    end else if (MbpBRight) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 838:62]
      perfCnts_16 <= _perfCnts_16_T_5; // @[src/main/scala/nutcore/backend/fu/CSR.scala 838:66]
    end else if (_T_693 & addr == 12'hb10) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      perfCnts_16 <= wdata; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
      perfCnts_17 <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
    end else if (MbpBWrong) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 838:62]
      perfCnts_17 <= _perfCnts_17_T_5; // @[src/main/scala/nutcore/backend/fu/CSR.scala 838:66]
    end else if (_T_693 & addr == 12'hb11) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      perfCnts_17 <= wdata; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
      perfCnts_18 <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
    end else if (MbpJRight) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 838:62]
      perfCnts_18 <= _perfCnts_18_T_5; // @[src/main/scala/nutcore/backend/fu/CSR.scala 838:66]
    end else if (_T_693 & addr == 12'hb12) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      perfCnts_18 <= wdata; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
      perfCnts_19 <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
    end else if (MbpJWrong) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 838:62]
      perfCnts_19 <= _perfCnts_19_T_5; // @[src/main/scala/nutcore/backend/fu/CSR.scala 838:66]
    end else if (_T_693 & addr == 12'hb13) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      perfCnts_19 <= wdata; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
      perfCnts_20 <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
    end else if (MbpIRight) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 838:62]
      perfCnts_20 <= _perfCnts_20_T_5; // @[src/main/scala/nutcore/backend/fu/CSR.scala 838:66]
    end else if (_T_693 & addr == 12'hb14) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      perfCnts_20 <= wdata; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
      perfCnts_21 <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
    end else if (MbpIWrong) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 838:62]
      perfCnts_21 <= _perfCnts_21_T_5; // @[src/main/scala/nutcore/backend/fu/CSR.scala 838:66]
    end else if (_T_693 & addr == 12'hb15) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      perfCnts_21 <= wdata; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
      perfCnts_22 <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
    end else if (MbpRRight) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 838:62]
      perfCnts_22 <= _perfCnts_22_T_5; // @[src/main/scala/nutcore/backend/fu/CSR.scala 838:66]
    end else if (_T_693 & addr == 12'hb16) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      perfCnts_22 <= wdata; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
      perfCnts_23 <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
    end else if (MbpRWrong) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 838:62]
      perfCnts_23 <= _perfCnts_23_T_5; // @[src/main/scala/nutcore/backend/fu/CSR.scala 838:66]
    end else if (_T_693 & addr == 12'hb17) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      perfCnts_23 <= wdata; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
      perfCnts_24 <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
    end else if (_T_693 & addr == 12'hb18) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      perfCnts_24 <= wdata; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
      perfCnts_25 <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
    end else if (Custom1) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 838:62]
      perfCnts_25 <= _perfCnts_25_T_5; // @[src/main/scala/nutcore/backend/fu/CSR.scala 838:66]
    end else if (_T_693 & addr == 12'hb19) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      perfCnts_25 <= wdata; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
      perfCnts_26 <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
    end else if (Custom2) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 838:62]
      perfCnts_26 <= _perfCnts_26_T_5; // @[src/main/scala/nutcore/backend/fu/CSR.scala 838:66]
    end else if (_T_693 & addr == 12'hb1a) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      perfCnts_26 <= wdata; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
      perfCnts_27 <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
    end else if (Custom3) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 838:62]
      perfCnts_27 <= _perfCnts_27_T_5; // @[src/main/scala/nutcore/backend/fu/CSR.scala 838:66]
    end else if (_T_693 & addr == 12'hb1b) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      perfCnts_27 <= wdata; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
      perfCnts_28 <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
    end else if (Custom4) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 838:62]
      perfCnts_28 <= _perfCnts_28_T_5; // @[src/main/scala/nutcore/backend/fu/CSR.scala 838:66]
    end else if (_T_693 & addr == 12'hb1c) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      perfCnts_28 <= wdata; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
      perfCnts_29 <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
    end else if (Custom5) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 838:62]
      perfCnts_29 <= _perfCnts_29_T_5; // @[src/main/scala/nutcore/backend/fu/CSR.scala 838:66]
    end else if (_T_693 & addr == 12'hb1d) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      perfCnts_29 <= wdata; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
      perfCnts_30 <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
    end else if (Custom6) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 838:62]
      perfCnts_30 <= _perfCnts_30_T_5; // @[src/main/scala/nutcore/backend/fu/CSR.scala 838:66]
    end else if (_T_693 & addr == 12'hb1e) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      perfCnts_30 <= wdata; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
      perfCnts_31 <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
    end else if (Custom7) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 838:62]
      perfCnts_31 <= _perfCnts_31_T_5; // @[src/main/scala/nutcore/backend/fu/CSR.scala 838:66]
    end else if (_T_693 & addr == 12'hb1f) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      perfCnts_31 <= wdata; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
      perfCnts_32 <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
    end else if (Custom8) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 838:62]
      perfCnts_32 <= _perfCnts_32_T_5; // @[src/main/scala/nutcore/backend/fu/CSR.scala 838:66]
    end else if (_T_693 & addr == 12'hb20) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      perfCnts_32 <= wdata; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
      perfCnts_33 <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
    end else if (_T_693 & addr == 12'hb21) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      perfCnts_33 <= wdata; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
      perfCnts_34 <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
    end else if (_T_693 & addr == 12'hb22) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      perfCnts_34 <= wdata; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
      perfCnts_35 <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
    end else if (_T_693 & addr == 12'hb23) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      perfCnts_35 <= wdata; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
      perfCnts_36 <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
    end else if (_T_693 & addr == 12'hb24) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      perfCnts_36 <= wdata; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
      perfCnts_37 <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
    end else if (_T_693 & addr == 12'hb25) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      perfCnts_37 <= wdata; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
      perfCnts_38 <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
    end else if (_T_693 & addr == 12'hb26) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      perfCnts_38 <= wdata; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
      perfCnts_39 <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
    end else if (_T_693 & addr == 12'hb27) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      perfCnts_39 <= wdata; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
      perfCnts_40 <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
    end else if (_T_693 & addr == 12'hb28) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      perfCnts_40 <= wdata; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
      perfCnts_41 <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
    end else if (_T_693 & addr == 12'hb29) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      perfCnts_41 <= wdata; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
      perfCnts_42 <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
    end else if (_T_693 & addr == 12'hb2a) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      perfCnts_42 <= wdata; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
      perfCnts_43 <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
    end else if (_T_693 & addr == 12'hb2b) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      perfCnts_43 <= wdata; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
      perfCnts_44 <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
    end else if (_T_693 & addr == 12'hb2c) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      perfCnts_44 <= wdata; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
      perfCnts_45 <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
    end else if (_T_693 & addr == 12'hb2d) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      perfCnts_45 <= wdata; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
      perfCnts_46 <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
    end else if (_T_693 & addr == 12'hb2e) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      perfCnts_46 <= wdata; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
      perfCnts_47 <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
    end else if (_T_693 & addr == 12'hb2f) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      perfCnts_47 <= wdata; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
      perfCnts_48 <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
    end else if (_T_693 & addr == 12'hb30) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      perfCnts_48 <= wdata; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
      perfCnts_49 <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
    end else if (perfCntCondMrawStall) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 838:62]
      perfCnts_49 <= _perfCnts_49_T_5; // @[src/main/scala/nutcore/backend/fu/CSR.scala 838:66]
    end else if (_T_693 & addr == 12'hb31) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      perfCnts_49 <= wdata; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
      perfCnts_50 <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
    end else if (perfCntCondMexuBusy) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 838:62]
      perfCnts_50 <= _perfCnts_50_T_5; // @[src/main/scala/nutcore/backend/fu/CSR.scala 838:66]
    end else if (_T_693 & addr == 12'hb32) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      perfCnts_50 <= wdata; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
      perfCnts_51 <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
    end else if (perfCntCondMloadStall) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 838:62]
      perfCnts_51 <= _perfCnts_51_T_5; // @[src/main/scala/nutcore/backend/fu/CSR.scala 838:66]
    end else if (_T_693 & addr == 12'hb33) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      perfCnts_51 <= wdata; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
      perfCnts_52 <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
    end else if (perfCntCondMstoreStall) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 838:62]
      perfCnts_52 <= _perfCnts_52_T_5; // @[src/main/scala/nutcore/backend/fu/CSR.scala 838:66]
    end else if (_T_693 & addr == 12'hb34) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      perfCnts_52 <= wdata; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
      perfCnts_53 <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
    end else if (perfCntCondISUIssue) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 838:62]
      perfCnts_53 <= _perfCnts_53_T_5; // @[src/main/scala/nutcore/backend/fu/CSR.scala 838:66]
    end else if (_T_693 & addr == 12'hb35) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      perfCnts_53 <= wdata; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
      perfCnts_54 <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
    end else if (_T_693 & addr == 12'hb36) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      perfCnts_54 <= wdata; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
      perfCnts_55 <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
    end else if (_T_693 & addr == 12'hb37) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      perfCnts_55 <= wdata; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
      perfCnts_56 <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
    end else if (_T_693 & addr == 12'hb38) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      perfCnts_56 <= wdata; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
      perfCnts_57 <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
    end else if (_T_693 & addr == 12'hb39) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      perfCnts_57 <= wdata; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
      perfCnts_58 <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
    end else if (_T_693 & addr == 12'hb3a) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      perfCnts_58 <= wdata; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
      perfCnts_59 <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
    end else if (_T_693 & addr == 12'hb3b) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      perfCnts_59 <= wdata; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
      perfCnts_60 <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
    end else if (_T_693 & addr == 12'hb3c) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      perfCnts_60 <= wdata; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
      perfCnts_61 <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
    end else if (_T_693 & addr == 12'hb3d) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      perfCnts_61 <= wdata; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
      perfCnts_62 <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
    end else if (_T_693 & addr == 12'hb3e) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      perfCnts_62 <= wdata; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
      perfCnts_63 <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
    end else if (_T_693 & addr == 12'hb3f) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      perfCnts_63 <= wdata; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
      perfCnts_64 <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
    end else if (_T_693 & addr == 12'hb40) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      perfCnts_64 <= wdata; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
      perfCnts_65 <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
    end else if (_T_693 & addr == 12'hb41) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      perfCnts_65 <= wdata; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
      perfCnts_66 <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
    end else if (_T_693 & addr == 12'hb42) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      perfCnts_66 <= wdata; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
      perfCnts_67 <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
    end else if (_T_693 & addr == 12'hb43) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      perfCnts_67 <= wdata; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
      perfCnts_68 <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
    end else if (_T_693 & addr == 12'hb44) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      perfCnts_68 <= wdata; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
      perfCnts_69 <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
    end else if (_T_693 & addr == 12'hb45) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      perfCnts_69 <= wdata; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
      perfCnts_70 <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
    end else if (_T_693 & addr == 12'hb46) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      perfCnts_70 <= wdata; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
      perfCnts_71 <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
    end else if (_T_693 & addr == 12'hb47) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      perfCnts_71 <= wdata; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
      perfCnts_72 <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
    end else if (_T_693 & addr == 12'hb48) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      perfCnts_72 <= wdata; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
      perfCnts_73 <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
    end else if (_T_693 & addr == 12'hb49) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      perfCnts_73 <= wdata; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
      perfCnts_74 <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
    end else if (_T_693 & addr == 12'hb4a) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      perfCnts_74 <= wdata; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
      perfCnts_75 <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
    end else if (_T_693 & addr == 12'hb4b) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      perfCnts_75 <= wdata; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
      perfCnts_76 <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
    end else if (_T_693 & addr == 12'hb4c) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      perfCnts_76 <= wdata; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
      perfCnts_77 <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
    end else if (_T_693 & addr == 12'hb4d) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      perfCnts_77 <= wdata; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
      perfCnts_78 <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
    end else if (_T_693 & addr == 12'hb4e) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      perfCnts_78 <= wdata; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
      perfCnts_79 <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
    end else if (_T_693 & addr == 12'hb4f) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      perfCnts_79 <= wdata; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
      perfCnts_80 <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
    end else if (_T_693 & addr == 12'hb50) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      perfCnts_80 <= wdata; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
      perfCnts_81 <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
    end else if (_T_693 & addr == 12'hb51) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      perfCnts_81 <= wdata; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
      perfCnts_82 <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
    end else if (_T_693 & addr == 12'hb52) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      perfCnts_82 <= wdata; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
      perfCnts_83 <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
    end else if (_T_693 & addr == 12'hb53) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      perfCnts_83 <= wdata; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
      perfCnts_84 <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
    end else if (_T_693 & addr == 12'hb54) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      perfCnts_84 <= wdata; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
      perfCnts_85 <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
    end else if (_T_693 & addr == 12'hb55) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      perfCnts_85 <= wdata; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
      perfCnts_86 <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
    end else if (_T_693 & addr == 12'hb56) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      perfCnts_86 <= wdata; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
      perfCnts_87 <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
    end else if (_T_693 & addr == 12'hb57) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      perfCnts_87 <= wdata; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
      perfCnts_88 <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
    end else if (_T_693 & addr == 12'hb58) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      perfCnts_88 <= wdata; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
      perfCnts_89 <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
    end else if (_T_693 & addr == 12'hb59) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      perfCnts_89 <= wdata; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
      perfCnts_90 <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
    end else if (_T_693 & addr == 12'hb5a) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      perfCnts_90 <= wdata; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
      perfCnts_91 <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
    end else if (_T_693 & addr == 12'hb5b) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      perfCnts_91 <= wdata; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
      perfCnts_92 <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
    end else if (_T_693 & addr == 12'hb5c) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      perfCnts_92 <= wdata; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
      perfCnts_93 <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
    end else if (_T_693 & addr == 12'hb5d) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      perfCnts_93 <= wdata; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
      perfCnts_94 <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
    end else if (_T_693 & addr == 12'hb5e) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      perfCnts_94 <= wdata; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
      perfCnts_95 <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
    end else if (_T_693 & addr == 12'hb5f) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      perfCnts_95 <= wdata; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
      perfCnts_96 <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
    end else if (_T_693 & addr == 12'hb60) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      perfCnts_96 <= wdata; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
      perfCnts_97 <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
    end else if (_T_693 & addr == 12'hb61) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      perfCnts_97 <= wdata; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
      perfCnts_98 <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
    end else if (_T_693 & addr == 12'hb62) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      perfCnts_98 <= wdata; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
      perfCnts_99 <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
    end else begin
      perfCnts_99 <= _perfCnts_99_T_6[63:0];
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
      perfCnts_100 <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
    end else begin
      perfCnts_100 <= _perfCnts_100_T_6[63:0];
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
      perfCnts_101 <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
    end else begin
      perfCnts_101 <= _perfCnts_101_T_6[63:0];
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
      perfCnts_102 <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
    end else if (_T_693 & addr == 12'hb66) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      perfCnts_102 <= wdata; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
      perfCnts_103 <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
    end else if (_T_693 & addr == 12'hb67) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      perfCnts_103 <= wdata; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
      perfCnts_104 <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
    end else if (_T_693 & addr == 12'hb68) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      perfCnts_104 <= wdata; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
      perfCnts_105 <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
    end else if (_T_693 & addr == 12'hb69) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      perfCnts_105 <= wdata; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
      perfCnts_106 <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
    end else if (_T_693 & addr == 12'hb6a) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      perfCnts_106 <= wdata; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
      perfCnts_107 <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
    end else if (_T_693 & addr == 12'hb6b) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      perfCnts_107 <= wdata; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
      perfCnts_108 <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
    end else if (_T_693 & addr == 12'hb6c) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      perfCnts_108 <= wdata; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
      perfCnts_109 <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
    end else if (_T_693 & addr == 12'hb6d) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      perfCnts_109 <= wdata; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
      perfCnts_110 <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
    end else if (_T_693 & addr == 12'hb6e) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      perfCnts_110 <= wdata; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
      perfCnts_111 <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
    end else if (_T_693 & addr == 12'hb6f) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      perfCnts_111 <= wdata; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
      perfCnts_112 <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
    end else if (_T_693 & addr == 12'hb70) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      perfCnts_112 <= wdata; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
      perfCnts_113 <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
    end else if (_T_693 & addr == 12'hb71) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      perfCnts_113 <= wdata; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
      perfCnts_114 <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
    end else if (_T_693 & addr == 12'hb72) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      perfCnts_114 <= wdata; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
      perfCnts_115 <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
    end else if (_T_693 & addr == 12'hb73) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      perfCnts_115 <= wdata; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
      perfCnts_116 <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
    end else if (_T_693 & addr == 12'hb74) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      perfCnts_116 <= wdata; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
      perfCnts_117 <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
    end else if (_T_693 & addr == 12'hb75) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      perfCnts_117 <= wdata; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
      perfCnts_118 <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
    end else if (_T_693 & addr == 12'hb76) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      perfCnts_118 <= wdata; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
      perfCnts_119 <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
    end else if (_T_693 & addr == 12'hb77) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      perfCnts_119 <= wdata; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
      perfCnts_120 <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
    end else if (_T_693 & addr == 12'hb78) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      perfCnts_120 <= wdata; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
      perfCnts_121 <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
    end else if (_T_693 & addr == 12'hb79) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      perfCnts_121 <= wdata; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
      perfCnts_122 <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
    end else if (_T_693 & addr == 12'hb7a) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      perfCnts_122 <= wdata; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
      perfCnts_123 <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
    end else if (_T_693 & addr == 12'hb7b) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      perfCnts_123 <= wdata; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
      perfCnts_124 <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
    end else if (_T_693 & addr == 12'hb7c) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      perfCnts_124 <= wdata; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
      perfCnts_125 <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
    end else if (_T_693 & addr == 12'hb7d) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      perfCnts_125 <= wdata; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
      perfCnts_126 <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
    end else if (_T_693 & addr == 12'hb7e) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      perfCnts_126 <= wdata; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
      perfCnts_127 <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 374:47]
    end else if (_T_693 & addr == 12'hb7f) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      perfCnts_127 <= wdata; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/utils/GTimer.scala 24:20]
      c <= 64'h0; // @[src/main/scala/utils/GTimer.scala 24:20]
    end else begin
      c <= _c_T_1; // @[src/main/scala/utils/GTimer.scala 25:7]
    end
    if (reset) begin // @[src/main/scala/utils/GTimer.scala 24:20]
      c_1 <= 64'h0; // @[src/main/scala/utils/GTimer.scala 24:20]
    end else begin
      c_1 <= _c_T_3; // @[src/main/scala/utils/GTimer.scala 25:7]
    end
    if (reset) begin // @[src/main/scala/utils/GTimer.scala 24:20]
      c_2 <= 64'h0; // @[src/main/scala/utils/GTimer.scala 24:20]
    end else begin
      c_2 <= _c_T_5; // @[src/main/scala/utils/GTimer.scala 25:7]
    end
    if (reset) begin // @[src/main/scala/utils/GTimer.scala 24:20]
      c_3 <= 64'h0; // @[src/main/scala/utils/GTimer.scala 24:20]
    end else begin
      c_3 <= _c_T_7; // @[src/main/scala/utils/GTimer.scala 25:7]
    end
    if (reset) begin // @[src/main/scala/utils/GTimer.scala 24:20]
      c_4 <= 64'h0; // @[src/main/scala/utils/GTimer.scala 24:20]
    end else begin
      c_4 <= _c_T_9; // @[src/main/scala/utils/GTimer.scala 25:7]
    end
    if (reset) begin // @[src/main/scala/utils/GTimer.scala 24:20]
      c_5 <= 64'h0; // @[src/main/scala/utils/GTimer.scala 24:20]
    end else begin
      c_5 <= _c_T_11; // @[src/main/scala/utils/GTimer.scala 25:7]
    end
    if (reset) begin // @[src/main/scala/utils/GTimer.scala 24:20]
      c_6 <= 64'h0; // @[src/main/scala/utils/GTimer.scala 24:20]
    end else begin
      c_6 <= _c_T_13; // @[src/main/scala/utils/GTimer.scala 25:7]
    end
    if (reset) begin // @[src/main/scala/utils/GTimer.scala 24:20]
      c_7 <= 64'h0; // @[src/main/scala/utils/GTimer.scala 24:20]
    end else begin
      c_7 <= _c_T_15; // @[src/main/scala/utils/GTimer.scala 25:7]
    end
    if (reset) begin // @[src/main/scala/utils/GTimer.scala 24:20]
      c_8 <= 64'h0; // @[src/main/scala/utils/GTimer.scala 24:20]
    end else begin
      c_8 <= _c_T_17; // @[src/main/scala/utils/GTimer.scala 25:7]
    end
    if (reset) begin // @[src/main/scala/utils/GTimer.scala 24:20]
      c_9 <= 64'h0; // @[src/main/scala/utils/GTimer.scala 24:20]
    end else begin
      c_9 <= _c_T_19; // @[src/main/scala/utils/GTimer.scala 25:7]
    end
    if (reset) begin // @[src/main/scala/utils/GTimer.scala 24:20]
      c_10 <= 64'h0; // @[src/main/scala/utils/GTimer.scala 24:20]
    end else begin
      c_10 <= _c_T_21; // @[src/main/scala/utils/GTimer.scala 25:7]
    end
    if (reset) begin // @[src/main/scala/utils/GTimer.scala 24:20]
      c_11 <= 64'h0; // @[src/main/scala/utils/GTimer.scala 24:20]
    end else begin
      c_11 <= _c_T_23; // @[src/main/scala/utils/GTimer.scala 25:7]
    end
    if (reset) begin // @[src/main/scala/utils/GTimer.scala 24:20]
      c_12 <= 64'h0; // @[src/main/scala/utils/GTimer.scala 24:20]
    end else begin
      c_12 <= _c_T_25; // @[src/main/scala/utils/GTimer.scala 25:7]
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1013 & ~reset) begin
          $fwrite(32'h80000002,"[%d] CSR: ",c); // @[src/main/scala/utils/Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1013 & _T_1015) begin
          $fwrite(32'h80000002,"csr write: pc %x addr %x rdata %x wdata %x func %x\n",io_cfIn_pc,addr,rdata,wdata,
            io_in_bits_func); // @[src/main/scala/utils/Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1013 & ~reset) begin
          $fwrite(32'h80000002,"[%d] CSR: ",c_2); // @[src/main/scala/utils/Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1013 & _T_1015) begin
          $fwrite(32'h80000002,"[MST] time %d pc %x mstatus %x mideleg %x medeleg %x mode %x\n",c_1,io_cfIn_pc,mstatus,
            mideleg,medeleg,priviledgeMode); // @[src/main/scala/utils/Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1024 & DISPLAY_ENABLE & ~reset) begin
          $fwrite(32'h80000002,"[%d] CSR: ",c_4); // @[src/main/scala/utils/Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_335 & _T_1015) begin
          $fwrite(32'h80000002,"[PF] %d: ipf %b tval %x := addr %x pc %x priviledgeMode %x\n",c_3,hasInstrPageFault,tval
            ,_tval_T_13,io_cfIn_pc,priviledgeMode); // @[src/main/scala/utils/Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1034 & DISPLAY_ENABLE & ~reset) begin
          $fwrite(32'h80000002,"[%d] CSR: ",c_6); // @[src/main/scala/utils/Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_337 & _T_1015) begin
          $fwrite(32'h80000002,"[ML] %d: addr %x pc %x priviledgeMode %x\n",c_5,_mtval_T_6,io_cfIn_pc,priviledgeMode); // @[src/main/scala/utils/Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1109 & ~reset) begin
          $fwrite(32'h80000002,"[%d] CSR: ",c_7); // @[src/main/scala/utils/Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1109 & _T_1015) begin
          $fwrite(32'h80000002,"excin %b excgen %b",_raiseExceptionVec_T,_raiseExceptionVec_T_1); // @[src/main/scala/utils/Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1109 & ~reset) begin
          $fwrite(32'h80000002,"[%d] CSR: ",c_8); // @[src/main/scala/utils/Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1109 & _T_1015) begin
          $fwrite(32'h80000002,"int/exc: pc %x int (%d):%x exc: (%d):%x\n",io_cfIn_pc,intrNO,_raiseIntr_T,exceptionNO,
            raiseExceptionVec); // @[src/main/scala/utils/Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1109 & ~reset) begin
          $fwrite(32'h80000002,"[%d] CSR: ",c_10); // @[src/main/scala/utils/Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1109 & _T_1015) begin
          $fwrite(32'h80000002,"[MST] time %d pc %x mstatus %x mideleg %x medeleg %x mode %x\n",c_9,io_cfIn_pc,mstatus,
            mideleg,medeleg,priviledgeMode); // @[src/main/scala/utils/Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1125 & ~reset) begin
          $fwrite(32'h80000002,"[%d] CSR: ",c_11); // @[src/main/scala/utils/Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1125 & _T_1015) begin
          $fwrite(32'h80000002,"redirect to %x\n",io_redirect_target); // @[src/main/scala/utils/Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1130 & ~reset) begin
          $fwrite(32'h80000002,"[%d] CSR: ",c_12); // @[src/main/scala/utils/Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1130 & _T_1015) begin
          $fwrite(32'h80000002,"satp reset\n"); // @[src/main/scala/utils/Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_1015) begin
          $fwrite(32'h80000002,"======== PerfCnt =========\n"); // @[src/main/scala/nutcore/backend/fu/CSR.scala 879:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_1015) begin
          $fwrite(32'h80000002,"%d <- Mcycle\n",perfCnts_0); // @[src/main/scala/nutcore/backend/fu/CSR.scala 881:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_1015) begin
          $fwrite(32'h80000002,"%d <- Minstret\n",perfCnts_2); // @[src/main/scala/nutcore/backend/fu/CSR.scala 881:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_1015) begin
          $fwrite(32'h80000002,"%d <- MultiCommit\n",perfCnts_3); // @[src/main/scala/nutcore/backend/fu/CSR.scala 881:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_1015) begin
          $fwrite(32'h80000002,"%d <- MimemStall\n",perfCnts_4); // @[src/main/scala/nutcore/backend/fu/CSR.scala 881:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_1015) begin
          $fwrite(32'h80000002,"%d <- MaluInstr\n",perfCnts_5); // @[src/main/scala/nutcore/backend/fu/CSR.scala 881:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_1015) begin
          $fwrite(32'h80000002,"%d <- MbruInstr\n",perfCnts_6); // @[src/main/scala/nutcore/backend/fu/CSR.scala 881:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_1015) begin
          $fwrite(32'h80000002,"%d <- MlsuInstr\n",perfCnts_7); // @[src/main/scala/nutcore/backend/fu/CSR.scala 881:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_1015) begin
          $fwrite(32'h80000002,"%d <- MmduInstr\n",perfCnts_8); // @[src/main/scala/nutcore/backend/fu/CSR.scala 881:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_1015) begin
          $fwrite(32'h80000002,"%d <- McsrInstr\n",perfCnts_9); // @[src/main/scala/nutcore/backend/fu/CSR.scala 881:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_1015) begin
          $fwrite(32'h80000002,"%d <- MloadInstr\n",perfCnts_10); // @[src/main/scala/nutcore/backend/fu/CSR.scala 881:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_1015) begin
          $fwrite(32'h80000002,"%d <- MmmioInstr\n",perfCnts_11); // @[src/main/scala/nutcore/backend/fu/CSR.scala 881:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_1015) begin
          $fwrite(32'h80000002,"%d <- MmulInstr\n",perfCnts_14); // @[src/main/scala/nutcore/backend/fu/CSR.scala 881:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_1015) begin
          $fwrite(32'h80000002,"%d <- MifuFlush\n",perfCnts_15); // @[src/main/scala/nutcore/backend/fu/CSR.scala 881:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_1015) begin
          $fwrite(32'h80000002,"%d <- MbpBRight\n",perfCnts_16); // @[src/main/scala/nutcore/backend/fu/CSR.scala 881:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_1015) begin
          $fwrite(32'h80000002,"%d <- MbpBWrong\n",perfCnts_17); // @[src/main/scala/nutcore/backend/fu/CSR.scala 881:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_1015) begin
          $fwrite(32'h80000002,"%d <- MbpJRight\n",perfCnts_18); // @[src/main/scala/nutcore/backend/fu/CSR.scala 881:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_1015) begin
          $fwrite(32'h80000002,"%d <- MbpJWrong\n",perfCnts_19); // @[src/main/scala/nutcore/backend/fu/CSR.scala 881:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_1015) begin
          $fwrite(32'h80000002,"%d <- MbpIRight\n",perfCnts_20); // @[src/main/scala/nutcore/backend/fu/CSR.scala 881:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_1015) begin
          $fwrite(32'h80000002,"%d <- MbpIWrong\n",perfCnts_21); // @[src/main/scala/nutcore/backend/fu/CSR.scala 881:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_1015) begin
          $fwrite(32'h80000002,"%d <- MbpRRight\n",perfCnts_22); // @[src/main/scala/nutcore/backend/fu/CSR.scala 881:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_1015) begin
          $fwrite(32'h80000002,"%d <- MbpRWrong\n",perfCnts_23); // @[src/main/scala/nutcore/backend/fu/CSR.scala 881:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_1015) begin
          $fwrite(32'h80000002,"%d <- Custom1\n",perfCnts_25); // @[src/main/scala/nutcore/backend/fu/CSR.scala 881:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_1015) begin
          $fwrite(32'h80000002,"%d <- Custom2\n",perfCnts_26); // @[src/main/scala/nutcore/backend/fu/CSR.scala 881:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_1015) begin
          $fwrite(32'h80000002,"%d <- Custom3\n",perfCnts_27); // @[src/main/scala/nutcore/backend/fu/CSR.scala 881:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_1015) begin
          $fwrite(32'h80000002,"%d <- Custom4\n",perfCnts_28); // @[src/main/scala/nutcore/backend/fu/CSR.scala 881:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_1015) begin
          $fwrite(32'h80000002,"%d <- Custom5\n",perfCnts_29); // @[src/main/scala/nutcore/backend/fu/CSR.scala 881:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_1015) begin
          $fwrite(32'h80000002,"%d <- Custom6\n",perfCnts_30); // @[src/main/scala/nutcore/backend/fu/CSR.scala 881:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_1015) begin
          $fwrite(32'h80000002,"%d <- Custom7\n",perfCnts_31); // @[src/main/scala/nutcore/backend/fu/CSR.scala 881:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_1015) begin
          $fwrite(32'h80000002,"%d <- Custom8\n",perfCnts_32); // @[src/main/scala/nutcore/backend/fu/CSR.scala 881:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_1015) begin
          $fwrite(32'h80000002,"%d <- MrawStall\n",perfCnts_49); // @[src/main/scala/nutcore/backend/fu/CSR.scala 881:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_1015) begin
          $fwrite(32'h80000002,"%d <- MexuBusy\n",perfCnts_50); // @[src/main/scala/nutcore/backend/fu/CSR.scala 881:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_1015) begin
          $fwrite(32'h80000002,"%d <- MloadStall\n",perfCnts_51); // @[src/main/scala/nutcore/backend/fu/CSR.scala 881:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_1015) begin
          $fwrite(32'h80000002,"%d <- MstoreStall\n",perfCnts_52); // @[src/main/scala/nutcore/backend/fu/CSR.scala 881:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_1015) begin
          $fwrite(32'h80000002,"%d <- ISUIssue\n",perfCnts_53); // @[src/main/scala/nutcore/backend/fu/CSR.scala 881:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_1015) begin
          $fwrite(32'h80000002,"======== PerfCntCSV =========\n\n"); // @[src/main/scala/nutcore/backend/fu/CSR.scala 883:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_1015) begin
          $fwrite(32'h80000002,"Mcycle, "); // @[src/main/scala/nutcore/backend/fu/CSR.scala 885:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_1015) begin
          $fwrite(32'h80000002,"Minstret, "); // @[src/main/scala/nutcore/backend/fu/CSR.scala 885:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_1015) begin
          $fwrite(32'h80000002,"MultiCommit, "); // @[src/main/scala/nutcore/backend/fu/CSR.scala 885:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_1015) begin
          $fwrite(32'h80000002,"MimemStall, "); // @[src/main/scala/nutcore/backend/fu/CSR.scala 885:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_1015) begin
          $fwrite(32'h80000002,"MaluInstr, "); // @[src/main/scala/nutcore/backend/fu/CSR.scala 885:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_1015) begin
          $fwrite(32'h80000002,"MbruInstr, "); // @[src/main/scala/nutcore/backend/fu/CSR.scala 885:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_1015) begin
          $fwrite(32'h80000002,"MlsuInstr, "); // @[src/main/scala/nutcore/backend/fu/CSR.scala 885:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_1015) begin
          $fwrite(32'h80000002,"MmduInstr, "); // @[src/main/scala/nutcore/backend/fu/CSR.scala 885:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_1015) begin
          $fwrite(32'h80000002,"McsrInstr, "); // @[src/main/scala/nutcore/backend/fu/CSR.scala 885:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_1015) begin
          $fwrite(32'h80000002,"MloadInstr, "); // @[src/main/scala/nutcore/backend/fu/CSR.scala 885:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_1015) begin
          $fwrite(32'h80000002,"MmmioInstr, "); // @[src/main/scala/nutcore/backend/fu/CSR.scala 885:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_1015) begin
          $fwrite(32'h80000002,"MmulInstr, "); // @[src/main/scala/nutcore/backend/fu/CSR.scala 885:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_1015) begin
          $fwrite(32'h80000002,"MifuFlush, "); // @[src/main/scala/nutcore/backend/fu/CSR.scala 885:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_1015) begin
          $fwrite(32'h80000002,"MbpBRight, "); // @[src/main/scala/nutcore/backend/fu/CSR.scala 885:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_1015) begin
          $fwrite(32'h80000002,"MbpBWrong, "); // @[src/main/scala/nutcore/backend/fu/CSR.scala 885:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_1015) begin
          $fwrite(32'h80000002,"MbpJRight, "); // @[src/main/scala/nutcore/backend/fu/CSR.scala 885:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_1015) begin
          $fwrite(32'h80000002,"MbpJWrong, "); // @[src/main/scala/nutcore/backend/fu/CSR.scala 885:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_1015) begin
          $fwrite(32'h80000002,"MbpIRight, "); // @[src/main/scala/nutcore/backend/fu/CSR.scala 885:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_1015) begin
          $fwrite(32'h80000002,"MbpIWrong, "); // @[src/main/scala/nutcore/backend/fu/CSR.scala 885:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_1015) begin
          $fwrite(32'h80000002,"MbpRRight, "); // @[src/main/scala/nutcore/backend/fu/CSR.scala 885:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_1015) begin
          $fwrite(32'h80000002,"MbpRWrong, "); // @[src/main/scala/nutcore/backend/fu/CSR.scala 885:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_1015) begin
          $fwrite(32'h80000002,"Custom1, "); // @[src/main/scala/nutcore/backend/fu/CSR.scala 885:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_1015) begin
          $fwrite(32'h80000002,"Custom2, "); // @[src/main/scala/nutcore/backend/fu/CSR.scala 885:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_1015) begin
          $fwrite(32'h80000002,"Custom3, "); // @[src/main/scala/nutcore/backend/fu/CSR.scala 885:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_1015) begin
          $fwrite(32'h80000002,"Custom4, "); // @[src/main/scala/nutcore/backend/fu/CSR.scala 885:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_1015) begin
          $fwrite(32'h80000002,"Custom5, "); // @[src/main/scala/nutcore/backend/fu/CSR.scala 885:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_1015) begin
          $fwrite(32'h80000002,"Custom6, "); // @[src/main/scala/nutcore/backend/fu/CSR.scala 885:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_1015) begin
          $fwrite(32'h80000002,"Custom7, "); // @[src/main/scala/nutcore/backend/fu/CSR.scala 885:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_1015) begin
          $fwrite(32'h80000002,"Custom8, "); // @[src/main/scala/nutcore/backend/fu/CSR.scala 885:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_1015) begin
          $fwrite(32'h80000002,"MrawStall, "); // @[src/main/scala/nutcore/backend/fu/CSR.scala 885:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_1015) begin
          $fwrite(32'h80000002,"MexuBusy, "); // @[src/main/scala/nutcore/backend/fu/CSR.scala 885:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_1015) begin
          $fwrite(32'h80000002,"MloadStall, "); // @[src/main/scala/nutcore/backend/fu/CSR.scala 885:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_1015) begin
          $fwrite(32'h80000002,"MstoreStall, "); // @[src/main/scala/nutcore/backend/fu/CSR.scala 885:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_1015) begin
          $fwrite(32'h80000002,"ISUIssue, "); // @[src/main/scala/nutcore/backend/fu/CSR.scala 885:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_1015) begin
          $fwrite(32'h80000002,"\n\n\n"); // @[src/main/scala/nutcore/backend/fu/CSR.scala 886:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_1015) begin
          $fwrite(32'h80000002,"%d, ",perfCnts_0); // @[src/main/scala/nutcore/backend/fu/CSR.scala 888:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_1015) begin
          $fwrite(32'h80000002,"%d, ",perfCnts_2); // @[src/main/scala/nutcore/backend/fu/CSR.scala 888:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_1015) begin
          $fwrite(32'h80000002,"%d, ",perfCnts_3); // @[src/main/scala/nutcore/backend/fu/CSR.scala 888:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_1015) begin
          $fwrite(32'h80000002,"%d, ",perfCnts_4); // @[src/main/scala/nutcore/backend/fu/CSR.scala 888:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_1015) begin
          $fwrite(32'h80000002,"%d, ",perfCnts_5); // @[src/main/scala/nutcore/backend/fu/CSR.scala 888:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_1015) begin
          $fwrite(32'h80000002,"%d, ",perfCnts_6); // @[src/main/scala/nutcore/backend/fu/CSR.scala 888:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_1015) begin
          $fwrite(32'h80000002,"%d, ",perfCnts_7); // @[src/main/scala/nutcore/backend/fu/CSR.scala 888:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_1015) begin
          $fwrite(32'h80000002,"%d, ",perfCnts_8); // @[src/main/scala/nutcore/backend/fu/CSR.scala 888:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_1015) begin
          $fwrite(32'h80000002,"%d, ",perfCnts_9); // @[src/main/scala/nutcore/backend/fu/CSR.scala 888:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_1015) begin
          $fwrite(32'h80000002,"%d, ",perfCnts_10); // @[src/main/scala/nutcore/backend/fu/CSR.scala 888:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_1015) begin
          $fwrite(32'h80000002,"%d, ",perfCnts_11); // @[src/main/scala/nutcore/backend/fu/CSR.scala 888:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_1015) begin
          $fwrite(32'h80000002,"%d, ",perfCnts_14); // @[src/main/scala/nutcore/backend/fu/CSR.scala 888:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_1015) begin
          $fwrite(32'h80000002,"%d, ",perfCnts_15); // @[src/main/scala/nutcore/backend/fu/CSR.scala 888:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_1015) begin
          $fwrite(32'h80000002,"%d, ",perfCnts_16); // @[src/main/scala/nutcore/backend/fu/CSR.scala 888:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_1015) begin
          $fwrite(32'h80000002,"%d, ",perfCnts_17); // @[src/main/scala/nutcore/backend/fu/CSR.scala 888:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_1015) begin
          $fwrite(32'h80000002,"%d, ",perfCnts_18); // @[src/main/scala/nutcore/backend/fu/CSR.scala 888:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_1015) begin
          $fwrite(32'h80000002,"%d, ",perfCnts_19); // @[src/main/scala/nutcore/backend/fu/CSR.scala 888:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_1015) begin
          $fwrite(32'h80000002,"%d, ",perfCnts_20); // @[src/main/scala/nutcore/backend/fu/CSR.scala 888:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_1015) begin
          $fwrite(32'h80000002,"%d, ",perfCnts_21); // @[src/main/scala/nutcore/backend/fu/CSR.scala 888:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_1015) begin
          $fwrite(32'h80000002,"%d, ",perfCnts_22); // @[src/main/scala/nutcore/backend/fu/CSR.scala 888:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_1015) begin
          $fwrite(32'h80000002,"%d, ",perfCnts_23); // @[src/main/scala/nutcore/backend/fu/CSR.scala 888:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_1015) begin
          $fwrite(32'h80000002,"%d, ",perfCnts_25); // @[src/main/scala/nutcore/backend/fu/CSR.scala 888:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_1015) begin
          $fwrite(32'h80000002,"%d, ",perfCnts_26); // @[src/main/scala/nutcore/backend/fu/CSR.scala 888:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_1015) begin
          $fwrite(32'h80000002,"%d, ",perfCnts_27); // @[src/main/scala/nutcore/backend/fu/CSR.scala 888:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_1015) begin
          $fwrite(32'h80000002,"%d, ",perfCnts_28); // @[src/main/scala/nutcore/backend/fu/CSR.scala 888:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_1015) begin
          $fwrite(32'h80000002,"%d, ",perfCnts_29); // @[src/main/scala/nutcore/backend/fu/CSR.scala 888:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_1015) begin
          $fwrite(32'h80000002,"%d, ",perfCnts_30); // @[src/main/scala/nutcore/backend/fu/CSR.scala 888:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_1015) begin
          $fwrite(32'h80000002,"%d, ",perfCnts_31); // @[src/main/scala/nutcore/backend/fu/CSR.scala 888:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_1015) begin
          $fwrite(32'h80000002,"%d, ",perfCnts_32); // @[src/main/scala/nutcore/backend/fu/CSR.scala 888:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_1015) begin
          $fwrite(32'h80000002,"%d, ",perfCnts_49); // @[src/main/scala/nutcore/backend/fu/CSR.scala 888:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_1015) begin
          $fwrite(32'h80000002,"%d, ",perfCnts_50); // @[src/main/scala/nutcore/backend/fu/CSR.scala 888:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_1015) begin
          $fwrite(32'h80000002,"%d, ",perfCnts_51); // @[src/main/scala/nutcore/backend/fu/CSR.scala 888:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_1015) begin
          $fwrite(32'h80000002,"%d, ",perfCnts_52); // @[src/main/scala/nutcore/backend/fu/CSR.scala 888:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_1015) begin
          $fwrite(32'h80000002,"%d, ",perfCnts_53); // @[src/main/scala/nutcore/backend/fu/CSR.scala 888:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_1015) begin
          $fwrite(32'h80000002,"\n\n\n"); // @[src/main/scala/nutcore/backend/fu/CSR.scala 889:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  mtvec = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  mcounteren = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  mcause = _RAND_2[63:0];
  _RAND_3 = {2{`RANDOM}};
  mtval = _RAND_3[63:0];
  _RAND_4 = {2{`RANDOM}};
  mepc = _RAND_4[63:0];
  _RAND_5 = {2{`RANDOM}};
  mie = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  mipReg = _RAND_6[63:0];
  _RAND_7 = {2{`RANDOM}};
  misa = _RAND_7[63:0];
  _RAND_8 = {2{`RANDOM}};
  mstatus = _RAND_8[63:0];
  _RAND_9 = {2{`RANDOM}};
  medeleg = _RAND_9[63:0];
  _RAND_10 = {2{`RANDOM}};
  mideleg = _RAND_10[63:0];
  _RAND_11 = {2{`RANDOM}};
  mscratch = _RAND_11[63:0];
  _RAND_12 = {2{`RANDOM}};
  pmpcfg0 = _RAND_12[63:0];
  _RAND_13 = {2{`RANDOM}};
  pmpcfg1 = _RAND_13[63:0];
  _RAND_14 = {2{`RANDOM}};
  pmpcfg2 = _RAND_14[63:0];
  _RAND_15 = {2{`RANDOM}};
  pmpcfg3 = _RAND_15[63:0];
  _RAND_16 = {2{`RANDOM}};
  pmpaddr0 = _RAND_16[63:0];
  _RAND_17 = {2{`RANDOM}};
  pmpaddr1 = _RAND_17[63:0];
  _RAND_18 = {2{`RANDOM}};
  pmpaddr2 = _RAND_18[63:0];
  _RAND_19 = {2{`RANDOM}};
  pmpaddr3 = _RAND_19[63:0];
  _RAND_20 = {2{`RANDOM}};
  stvec = _RAND_20[63:0];
  _RAND_21 = {2{`RANDOM}};
  satp = _RAND_21[63:0];
  _RAND_22 = {2{`RANDOM}};
  sepc = _RAND_22[63:0];
  _RAND_23 = {2{`RANDOM}};
  scause = _RAND_23[63:0];
  _RAND_24 = {2{`RANDOM}};
  stval = _RAND_24[63:0];
  _RAND_25 = {2{`RANDOM}};
  sscratch = _RAND_25[63:0];
  _RAND_26 = {2{`RANDOM}};
  scounteren = _RAND_26[63:0];
  _RAND_27 = {1{`RANDOM}};
  lr = _RAND_27[0:0];
  _RAND_28 = {2{`RANDOM}};
  lrAddr = _RAND_28[63:0];
  _RAND_29 = {1{`RANDOM}};
  priviledgeMode = _RAND_29[1:0];
  _RAND_30 = {2{`RANDOM}};
  perfCnts_0 = _RAND_30[63:0];
  _RAND_31 = {2{`RANDOM}};
  perfCnts_1 = _RAND_31[63:0];
  _RAND_32 = {2{`RANDOM}};
  perfCnts_2 = _RAND_32[63:0];
  _RAND_33 = {2{`RANDOM}};
  perfCnts_3 = _RAND_33[63:0];
  _RAND_34 = {2{`RANDOM}};
  perfCnts_4 = _RAND_34[63:0];
  _RAND_35 = {2{`RANDOM}};
  perfCnts_5 = _RAND_35[63:0];
  _RAND_36 = {2{`RANDOM}};
  perfCnts_6 = _RAND_36[63:0];
  _RAND_37 = {2{`RANDOM}};
  perfCnts_7 = _RAND_37[63:0];
  _RAND_38 = {2{`RANDOM}};
  perfCnts_8 = _RAND_38[63:0];
  _RAND_39 = {2{`RANDOM}};
  perfCnts_9 = _RAND_39[63:0];
  _RAND_40 = {2{`RANDOM}};
  perfCnts_10 = _RAND_40[63:0];
  _RAND_41 = {2{`RANDOM}};
  perfCnts_11 = _RAND_41[63:0];
  _RAND_42 = {2{`RANDOM}};
  perfCnts_12 = _RAND_42[63:0];
  _RAND_43 = {2{`RANDOM}};
  perfCnts_13 = _RAND_43[63:0];
  _RAND_44 = {2{`RANDOM}};
  perfCnts_14 = _RAND_44[63:0];
  _RAND_45 = {2{`RANDOM}};
  perfCnts_15 = _RAND_45[63:0];
  _RAND_46 = {2{`RANDOM}};
  perfCnts_16 = _RAND_46[63:0];
  _RAND_47 = {2{`RANDOM}};
  perfCnts_17 = _RAND_47[63:0];
  _RAND_48 = {2{`RANDOM}};
  perfCnts_18 = _RAND_48[63:0];
  _RAND_49 = {2{`RANDOM}};
  perfCnts_19 = _RAND_49[63:0];
  _RAND_50 = {2{`RANDOM}};
  perfCnts_20 = _RAND_50[63:0];
  _RAND_51 = {2{`RANDOM}};
  perfCnts_21 = _RAND_51[63:0];
  _RAND_52 = {2{`RANDOM}};
  perfCnts_22 = _RAND_52[63:0];
  _RAND_53 = {2{`RANDOM}};
  perfCnts_23 = _RAND_53[63:0];
  _RAND_54 = {2{`RANDOM}};
  perfCnts_24 = _RAND_54[63:0];
  _RAND_55 = {2{`RANDOM}};
  perfCnts_25 = _RAND_55[63:0];
  _RAND_56 = {2{`RANDOM}};
  perfCnts_26 = _RAND_56[63:0];
  _RAND_57 = {2{`RANDOM}};
  perfCnts_27 = _RAND_57[63:0];
  _RAND_58 = {2{`RANDOM}};
  perfCnts_28 = _RAND_58[63:0];
  _RAND_59 = {2{`RANDOM}};
  perfCnts_29 = _RAND_59[63:0];
  _RAND_60 = {2{`RANDOM}};
  perfCnts_30 = _RAND_60[63:0];
  _RAND_61 = {2{`RANDOM}};
  perfCnts_31 = _RAND_61[63:0];
  _RAND_62 = {2{`RANDOM}};
  perfCnts_32 = _RAND_62[63:0];
  _RAND_63 = {2{`RANDOM}};
  perfCnts_33 = _RAND_63[63:0];
  _RAND_64 = {2{`RANDOM}};
  perfCnts_34 = _RAND_64[63:0];
  _RAND_65 = {2{`RANDOM}};
  perfCnts_35 = _RAND_65[63:0];
  _RAND_66 = {2{`RANDOM}};
  perfCnts_36 = _RAND_66[63:0];
  _RAND_67 = {2{`RANDOM}};
  perfCnts_37 = _RAND_67[63:0];
  _RAND_68 = {2{`RANDOM}};
  perfCnts_38 = _RAND_68[63:0];
  _RAND_69 = {2{`RANDOM}};
  perfCnts_39 = _RAND_69[63:0];
  _RAND_70 = {2{`RANDOM}};
  perfCnts_40 = _RAND_70[63:0];
  _RAND_71 = {2{`RANDOM}};
  perfCnts_41 = _RAND_71[63:0];
  _RAND_72 = {2{`RANDOM}};
  perfCnts_42 = _RAND_72[63:0];
  _RAND_73 = {2{`RANDOM}};
  perfCnts_43 = _RAND_73[63:0];
  _RAND_74 = {2{`RANDOM}};
  perfCnts_44 = _RAND_74[63:0];
  _RAND_75 = {2{`RANDOM}};
  perfCnts_45 = _RAND_75[63:0];
  _RAND_76 = {2{`RANDOM}};
  perfCnts_46 = _RAND_76[63:0];
  _RAND_77 = {2{`RANDOM}};
  perfCnts_47 = _RAND_77[63:0];
  _RAND_78 = {2{`RANDOM}};
  perfCnts_48 = _RAND_78[63:0];
  _RAND_79 = {2{`RANDOM}};
  perfCnts_49 = _RAND_79[63:0];
  _RAND_80 = {2{`RANDOM}};
  perfCnts_50 = _RAND_80[63:0];
  _RAND_81 = {2{`RANDOM}};
  perfCnts_51 = _RAND_81[63:0];
  _RAND_82 = {2{`RANDOM}};
  perfCnts_52 = _RAND_82[63:0];
  _RAND_83 = {2{`RANDOM}};
  perfCnts_53 = _RAND_83[63:0];
  _RAND_84 = {2{`RANDOM}};
  perfCnts_54 = _RAND_84[63:0];
  _RAND_85 = {2{`RANDOM}};
  perfCnts_55 = _RAND_85[63:0];
  _RAND_86 = {2{`RANDOM}};
  perfCnts_56 = _RAND_86[63:0];
  _RAND_87 = {2{`RANDOM}};
  perfCnts_57 = _RAND_87[63:0];
  _RAND_88 = {2{`RANDOM}};
  perfCnts_58 = _RAND_88[63:0];
  _RAND_89 = {2{`RANDOM}};
  perfCnts_59 = _RAND_89[63:0];
  _RAND_90 = {2{`RANDOM}};
  perfCnts_60 = _RAND_90[63:0];
  _RAND_91 = {2{`RANDOM}};
  perfCnts_61 = _RAND_91[63:0];
  _RAND_92 = {2{`RANDOM}};
  perfCnts_62 = _RAND_92[63:0];
  _RAND_93 = {2{`RANDOM}};
  perfCnts_63 = _RAND_93[63:0];
  _RAND_94 = {2{`RANDOM}};
  perfCnts_64 = _RAND_94[63:0];
  _RAND_95 = {2{`RANDOM}};
  perfCnts_65 = _RAND_95[63:0];
  _RAND_96 = {2{`RANDOM}};
  perfCnts_66 = _RAND_96[63:0];
  _RAND_97 = {2{`RANDOM}};
  perfCnts_67 = _RAND_97[63:0];
  _RAND_98 = {2{`RANDOM}};
  perfCnts_68 = _RAND_98[63:0];
  _RAND_99 = {2{`RANDOM}};
  perfCnts_69 = _RAND_99[63:0];
  _RAND_100 = {2{`RANDOM}};
  perfCnts_70 = _RAND_100[63:0];
  _RAND_101 = {2{`RANDOM}};
  perfCnts_71 = _RAND_101[63:0];
  _RAND_102 = {2{`RANDOM}};
  perfCnts_72 = _RAND_102[63:0];
  _RAND_103 = {2{`RANDOM}};
  perfCnts_73 = _RAND_103[63:0];
  _RAND_104 = {2{`RANDOM}};
  perfCnts_74 = _RAND_104[63:0];
  _RAND_105 = {2{`RANDOM}};
  perfCnts_75 = _RAND_105[63:0];
  _RAND_106 = {2{`RANDOM}};
  perfCnts_76 = _RAND_106[63:0];
  _RAND_107 = {2{`RANDOM}};
  perfCnts_77 = _RAND_107[63:0];
  _RAND_108 = {2{`RANDOM}};
  perfCnts_78 = _RAND_108[63:0];
  _RAND_109 = {2{`RANDOM}};
  perfCnts_79 = _RAND_109[63:0];
  _RAND_110 = {2{`RANDOM}};
  perfCnts_80 = _RAND_110[63:0];
  _RAND_111 = {2{`RANDOM}};
  perfCnts_81 = _RAND_111[63:0];
  _RAND_112 = {2{`RANDOM}};
  perfCnts_82 = _RAND_112[63:0];
  _RAND_113 = {2{`RANDOM}};
  perfCnts_83 = _RAND_113[63:0];
  _RAND_114 = {2{`RANDOM}};
  perfCnts_84 = _RAND_114[63:0];
  _RAND_115 = {2{`RANDOM}};
  perfCnts_85 = _RAND_115[63:0];
  _RAND_116 = {2{`RANDOM}};
  perfCnts_86 = _RAND_116[63:0];
  _RAND_117 = {2{`RANDOM}};
  perfCnts_87 = _RAND_117[63:0];
  _RAND_118 = {2{`RANDOM}};
  perfCnts_88 = _RAND_118[63:0];
  _RAND_119 = {2{`RANDOM}};
  perfCnts_89 = _RAND_119[63:0];
  _RAND_120 = {2{`RANDOM}};
  perfCnts_90 = _RAND_120[63:0];
  _RAND_121 = {2{`RANDOM}};
  perfCnts_91 = _RAND_121[63:0];
  _RAND_122 = {2{`RANDOM}};
  perfCnts_92 = _RAND_122[63:0];
  _RAND_123 = {2{`RANDOM}};
  perfCnts_93 = _RAND_123[63:0];
  _RAND_124 = {2{`RANDOM}};
  perfCnts_94 = _RAND_124[63:0];
  _RAND_125 = {2{`RANDOM}};
  perfCnts_95 = _RAND_125[63:0];
  _RAND_126 = {2{`RANDOM}};
  perfCnts_96 = _RAND_126[63:0];
  _RAND_127 = {2{`RANDOM}};
  perfCnts_97 = _RAND_127[63:0];
  _RAND_128 = {2{`RANDOM}};
  perfCnts_98 = _RAND_128[63:0];
  _RAND_129 = {2{`RANDOM}};
  perfCnts_99 = _RAND_129[63:0];
  _RAND_130 = {2{`RANDOM}};
  perfCnts_100 = _RAND_130[63:0];
  _RAND_131 = {2{`RANDOM}};
  perfCnts_101 = _RAND_131[63:0];
  _RAND_132 = {2{`RANDOM}};
  perfCnts_102 = _RAND_132[63:0];
  _RAND_133 = {2{`RANDOM}};
  perfCnts_103 = _RAND_133[63:0];
  _RAND_134 = {2{`RANDOM}};
  perfCnts_104 = _RAND_134[63:0];
  _RAND_135 = {2{`RANDOM}};
  perfCnts_105 = _RAND_135[63:0];
  _RAND_136 = {2{`RANDOM}};
  perfCnts_106 = _RAND_136[63:0];
  _RAND_137 = {2{`RANDOM}};
  perfCnts_107 = _RAND_137[63:0];
  _RAND_138 = {2{`RANDOM}};
  perfCnts_108 = _RAND_138[63:0];
  _RAND_139 = {2{`RANDOM}};
  perfCnts_109 = _RAND_139[63:0];
  _RAND_140 = {2{`RANDOM}};
  perfCnts_110 = _RAND_140[63:0];
  _RAND_141 = {2{`RANDOM}};
  perfCnts_111 = _RAND_141[63:0];
  _RAND_142 = {2{`RANDOM}};
  perfCnts_112 = _RAND_142[63:0];
  _RAND_143 = {2{`RANDOM}};
  perfCnts_113 = _RAND_143[63:0];
  _RAND_144 = {2{`RANDOM}};
  perfCnts_114 = _RAND_144[63:0];
  _RAND_145 = {2{`RANDOM}};
  perfCnts_115 = _RAND_145[63:0];
  _RAND_146 = {2{`RANDOM}};
  perfCnts_116 = _RAND_146[63:0];
  _RAND_147 = {2{`RANDOM}};
  perfCnts_117 = _RAND_147[63:0];
  _RAND_148 = {2{`RANDOM}};
  perfCnts_118 = _RAND_148[63:0];
  _RAND_149 = {2{`RANDOM}};
  perfCnts_119 = _RAND_149[63:0];
  _RAND_150 = {2{`RANDOM}};
  perfCnts_120 = _RAND_150[63:0];
  _RAND_151 = {2{`RANDOM}};
  perfCnts_121 = _RAND_151[63:0];
  _RAND_152 = {2{`RANDOM}};
  perfCnts_122 = _RAND_152[63:0];
  _RAND_153 = {2{`RANDOM}};
  perfCnts_123 = _RAND_153[63:0];
  _RAND_154 = {2{`RANDOM}};
  perfCnts_124 = _RAND_154[63:0];
  _RAND_155 = {2{`RANDOM}};
  perfCnts_125 = _RAND_155[63:0];
  _RAND_156 = {2{`RANDOM}};
  perfCnts_126 = _RAND_156[63:0];
  _RAND_157 = {2{`RANDOM}};
  perfCnts_127 = _RAND_157[63:0];
  _RAND_158 = {2{`RANDOM}};
  c = _RAND_158[63:0];
  _RAND_159 = {2{`RANDOM}};
  c_1 = _RAND_159[63:0];
  _RAND_160 = {2{`RANDOM}};
  c_2 = _RAND_160[63:0];
  _RAND_161 = {2{`RANDOM}};
  c_3 = _RAND_161[63:0];
  _RAND_162 = {2{`RANDOM}};
  c_4 = _RAND_162[63:0];
  _RAND_163 = {2{`RANDOM}};
  c_5 = _RAND_163[63:0];
  _RAND_164 = {2{`RANDOM}};
  c_6 = _RAND_164[63:0];
  _RAND_165 = {2{`RANDOM}};
  c_7 = _RAND_165[63:0];
  _RAND_166 = {2{`RANDOM}};
  c_8 = _RAND_166[63:0];
  _RAND_167 = {2{`RANDOM}};
  c_9 = _RAND_167[63:0];
  _RAND_168 = {2{`RANDOM}};
  c_10 = _RAND_168[63:0];
  _RAND_169 = {2{`RANDOM}};
  c_11 = _RAND_169[63:0];
  _RAND_170 = {2{`RANDOM}};
  c_12 = _RAND_170[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module MOU(
  input         clock,
  input         reset,
  input         io_in_valid, // @[src/main/scala/nutcore/backend/fu/MOU.scala 38:14]
  input  [6:0]  io_in_bits_func, // @[src/main/scala/nutcore/backend/fu/MOU.scala 38:14]
  input  [38:0] io_cfIn_pc, // @[src/main/scala/nutcore/backend/fu/MOU.scala 38:14]
  output [38:0] io_redirect_target, // @[src/main/scala/nutcore/backend/fu/MOU.scala 38:14]
  output        io_redirect_valid, // @[src/main/scala/nutcore/backend/fu/MOU.scala 38:14]
  input         DISPLAY_ENABLE,
  output        _WIRE_11,
  output        _WIRE_1_4
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  wire  flushICache = io_in_valid & io_in_bits_func == 7'h1; // @[src/main/scala/nutcore/backend/fu/MOU.scala 52:27]
  reg [63:0] c; // @[src/main/scala/utils/GTimer.scala 24:20]
  wire [63:0] _c_T_1 = c + 64'h1; // @[src/main/scala/utils/GTimer.scala 25:12]
  wire  _T = flushICache & DISPLAY_ENABLE; // @[src/main/scala/utils/Debug.scala 55:16]
  wire  _T_2 = ~reset; // @[src/main/scala/utils/Debug.scala 56:24]
  wire  flushTLB = io_in_valid & io_in_bits_func == 7'h2; // @[src/main/scala/nutcore/backend/fu/MOU.scala 56:24]
  reg [63:0] c_1; // @[src/main/scala/utils/GTimer.scala 24:20]
  wire [63:0] _c_T_3 = c_1 + 64'h1; // @[src/main/scala/utils/GTimer.scala 25:12]
  wire  _T_5 = flushTLB & DISPLAY_ENABLE; // @[src/main/scala/utils/Debug.scala 55:16]
  wire  _WIRE = flushICache; // @[src/main/scala/nutcore/backend/fu/MOU.scala 52:27]
  wire  _WIRE_1 = flushTLB; // @[src/main/scala/nutcore/backend/fu/MOU.scala 56:24]
  assign io_redirect_target = io_cfIn_pc + 39'h4; // @[src/main/scala/nutcore/backend/fu/MOU.scala 49:36]
  assign io_redirect_valid = io_in_valid; // @[src/main/scala/nutcore/backend/fu/MOU.scala 50:21]
  assign _WIRE_11 = _WIRE;
  assign _WIRE_1_4 = _WIRE_1;
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/utils/GTimer.scala 24:20]
      c <= 64'h0; // @[src/main/scala/utils/GTimer.scala 24:20]
    end else begin
      c <= _c_T_1; // @[src/main/scala/utils/GTimer.scala 25:7]
    end
    if (reset) begin // @[src/main/scala/utils/GTimer.scala 24:20]
      c_1 <= 64'h0; // @[src/main/scala/utils/GTimer.scala 24:20]
    end else begin
      c_1 <= _c_T_3; // @[src/main/scala/utils/GTimer.scala 25:7]
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T & ~reset) begin
          $fwrite(32'h80000002,"[%d] MOU: ",c); // @[src/main/scala/utils/Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T & _T_2) begin
          $fwrite(32'h80000002,"Flush I$ at %x\n",io_cfIn_pc); // @[src/main/scala/utils/Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_5 & ~reset) begin
          $fwrite(32'h80000002,"[%d] MOU: ",c_1); // @[src/main/scala/utils/Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_5 & _T_2) begin
          $fwrite(32'h80000002,"Sfence.vma at %x\n",io_cfIn_pc); // @[src/main/scala/utils/Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  c = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  c_1 = _RAND_1[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module EXU(
  input         clock,
  input         reset,
  output        io__in_ready, // @[src/main/scala/nutcore/backend/seq/EXU.scala 29:14]
  input         io__in_valid, // @[src/main/scala/nutcore/backend/seq/EXU.scala 29:14]
  input  [63:0] io__in_bits_cf_instr, // @[src/main/scala/nutcore/backend/seq/EXU.scala 29:14]
  input  [38:0] io__in_bits_cf_pc, // @[src/main/scala/nutcore/backend/seq/EXU.scala 29:14]
  input  [38:0] io__in_bits_cf_pnpc, // @[src/main/scala/nutcore/backend/seq/EXU.scala 29:14]
  input         io__in_bits_cf_exceptionVec_1, // @[src/main/scala/nutcore/backend/seq/EXU.scala 29:14]
  input         io__in_bits_cf_exceptionVec_2, // @[src/main/scala/nutcore/backend/seq/EXU.scala 29:14]
  input         io__in_bits_cf_exceptionVec_12, // @[src/main/scala/nutcore/backend/seq/EXU.scala 29:14]
  input         io__in_bits_cf_intrVec_0, // @[src/main/scala/nutcore/backend/seq/EXU.scala 29:14]
  input         io__in_bits_cf_intrVec_1, // @[src/main/scala/nutcore/backend/seq/EXU.scala 29:14]
  input         io__in_bits_cf_intrVec_2, // @[src/main/scala/nutcore/backend/seq/EXU.scala 29:14]
  input         io__in_bits_cf_intrVec_3, // @[src/main/scala/nutcore/backend/seq/EXU.scala 29:14]
  input         io__in_bits_cf_intrVec_4, // @[src/main/scala/nutcore/backend/seq/EXU.scala 29:14]
  input         io__in_bits_cf_intrVec_5, // @[src/main/scala/nutcore/backend/seq/EXU.scala 29:14]
  input         io__in_bits_cf_intrVec_6, // @[src/main/scala/nutcore/backend/seq/EXU.scala 29:14]
  input         io__in_bits_cf_intrVec_7, // @[src/main/scala/nutcore/backend/seq/EXU.scala 29:14]
  input         io__in_bits_cf_intrVec_8, // @[src/main/scala/nutcore/backend/seq/EXU.scala 29:14]
  input         io__in_bits_cf_intrVec_9, // @[src/main/scala/nutcore/backend/seq/EXU.scala 29:14]
  input         io__in_bits_cf_intrVec_10, // @[src/main/scala/nutcore/backend/seq/EXU.scala 29:14]
  input         io__in_bits_cf_intrVec_11, // @[src/main/scala/nutcore/backend/seq/EXU.scala 29:14]
  input  [3:0]  io__in_bits_cf_brIdx, // @[src/main/scala/nutcore/backend/seq/EXU.scala 29:14]
  input         io__in_bits_cf_crossPageIPFFix, // @[src/main/scala/nutcore/backend/seq/EXU.scala 29:14]
  input  [2:0]  io__in_bits_ctrl_fuType, // @[src/main/scala/nutcore/backend/seq/EXU.scala 29:14]
  input  [6:0]  io__in_bits_ctrl_fuOpType, // @[src/main/scala/nutcore/backend/seq/EXU.scala 29:14]
  input         io__in_bits_ctrl_rfWen, // @[src/main/scala/nutcore/backend/seq/EXU.scala 29:14]
  input  [4:0]  io__in_bits_ctrl_rfDest, // @[src/main/scala/nutcore/backend/seq/EXU.scala 29:14]
  input         io__in_bits_ctrl_isNutCoreTrap, // @[src/main/scala/nutcore/backend/seq/EXU.scala 29:14]
  input  [63:0] io__in_bits_data_src1, // @[src/main/scala/nutcore/backend/seq/EXU.scala 29:14]
  input  [63:0] io__in_bits_data_src2, // @[src/main/scala/nutcore/backend/seq/EXU.scala 29:14]
  input  [63:0] io__in_bits_data_imm, // @[src/main/scala/nutcore/backend/seq/EXU.scala 29:14]
  input         io__out_ready, // @[src/main/scala/nutcore/backend/seq/EXU.scala 29:14]
  output        io__out_valid, // @[src/main/scala/nutcore/backend/seq/EXU.scala 29:14]
  output [63:0] io__out_bits_decode_cf_instr, // @[src/main/scala/nutcore/backend/seq/EXU.scala 29:14]
  output [38:0] io__out_bits_decode_cf_pc, // @[src/main/scala/nutcore/backend/seq/EXU.scala 29:14]
  output [38:0] io__out_bits_decode_cf_redirect_target, // @[src/main/scala/nutcore/backend/seq/EXU.scala 29:14]
  output        io__out_bits_decode_cf_redirect_valid, // @[src/main/scala/nutcore/backend/seq/EXU.scala 29:14]
  output [2:0]  io__out_bits_decode_ctrl_fuType, // @[src/main/scala/nutcore/backend/seq/EXU.scala 29:14]
  output        io__out_bits_decode_ctrl_rfWen, // @[src/main/scala/nutcore/backend/seq/EXU.scala 29:14]
  output [4:0]  io__out_bits_decode_ctrl_rfDest, // @[src/main/scala/nutcore/backend/seq/EXU.scala 29:14]
  output        io__out_bits_isMMIO, // @[src/main/scala/nutcore/backend/seq/EXU.scala 29:14]
  output [63:0] io__out_bits_intrNO, // @[src/main/scala/nutcore/backend/seq/EXU.scala 29:14]
  output [63:0] io__out_bits_commits_0, // @[src/main/scala/nutcore/backend/seq/EXU.scala 29:14]
  output [63:0] io__out_bits_commits_1, // @[src/main/scala/nutcore/backend/seq/EXU.scala 29:14]
  output [63:0] io__out_bits_commits_2, // @[src/main/scala/nutcore/backend/seq/EXU.scala 29:14]
  output [63:0] io__out_bits_commits_3, // @[src/main/scala/nutcore/backend/seq/EXU.scala 29:14]
  input         io__flush, // @[src/main/scala/nutcore/backend/seq/EXU.scala 29:14]
  input         io__dmem_req_ready, // @[src/main/scala/nutcore/backend/seq/EXU.scala 29:14]
  output        io__dmem_req_valid, // @[src/main/scala/nutcore/backend/seq/EXU.scala 29:14]
  output [38:0] io__dmem_req_bits_addr, // @[src/main/scala/nutcore/backend/seq/EXU.scala 29:14]
  output [2:0]  io__dmem_req_bits_size, // @[src/main/scala/nutcore/backend/seq/EXU.scala 29:14]
  output [3:0]  io__dmem_req_bits_cmd, // @[src/main/scala/nutcore/backend/seq/EXU.scala 29:14]
  output [7:0]  io__dmem_req_bits_wmask, // @[src/main/scala/nutcore/backend/seq/EXU.scala 29:14]
  output [63:0] io__dmem_req_bits_wdata, // @[src/main/scala/nutcore/backend/seq/EXU.scala 29:14]
  input         io__dmem_resp_valid, // @[src/main/scala/nutcore/backend/seq/EXU.scala 29:14]
  input  [63:0] io__dmem_resp_bits_rdata, // @[src/main/scala/nutcore/backend/seq/EXU.scala 29:14]
  output        io__forward_valid, // @[src/main/scala/nutcore/backend/seq/EXU.scala 29:14]
  output        io__forward_wb_rfWen, // @[src/main/scala/nutcore/backend/seq/EXU.scala 29:14]
  output [4:0]  io__forward_wb_rfDest, // @[src/main/scala/nutcore/backend/seq/EXU.scala 29:14]
  output [63:0] io__forward_wb_rfData, // @[src/main/scala/nutcore/backend/seq/EXU.scala 29:14]
  output [2:0]  io__forward_fuType, // @[src/main/scala/nutcore/backend/seq/EXU.scala 29:14]
  output [1:0]  io__memMMU_imem_priviledgeMode, // @[src/main/scala/nutcore/backend/seq/EXU.scala 29:14]
  output [1:0]  io__memMMU_dmem_priviledgeMode, // @[src/main/scala/nutcore/backend/seq/EXU.scala 29:14]
  output        io__memMMU_dmem_status_sum, // @[src/main/scala/nutcore/backend/seq/EXU.scala 29:14]
  output        io__memMMU_dmem_status_mxr, // @[src/main/scala/nutcore/backend/seq/EXU.scala 29:14]
  input         io__memMMU_dmem_loadPF, // @[src/main/scala/nutcore/backend/seq/EXU.scala 29:14]
  input         io__memMMU_dmem_storePF, // @[src/main/scala/nutcore/backend/seq/EXU.scala 29:14]
  input  [38:0] io__memMMU_dmem_addr, // @[src/main/scala/nutcore/backend/seq/EXU.scala 29:14]
  input         io_extra_meip_0,
  output        REG_valid,
  output [38:0] REG_pc,
  output        REG_isMissPredict,
  output [38:0] REG_actualTarget,
  output        REG_actualTaken,
  output [6:0]  REG_fuOpType,
  output [1:0]  REG_btbType,
  output        REG_isRVC,
  output        _WIRE_6,
  input         _WIRE_1_0,
  output [63:0] satp,
  input         DISPLAY_ENABLE,
  input         _WIRE_1_1,
  input         _WIRE_8,
  input         _WIRE_11,
  input         _WIRE_2_2,
  input         io_extra_mtip,
  output        _WIRE_12,
  input         falseWire,
  output        _WIRE_1_4,
  output [11:0] _WIRE_14,
  input         _WIRE_2_3,
  input         _WIRE_16,
  input         _WIRE_17,
  input         r_0,
  input         io_extra_msip,
  input         io_in_valid
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  wire  alu_clock; // @[src/main/scala/nutcore/backend/seq/EXU.scala 46:19]
  wire  alu_reset; // @[src/main/scala/nutcore/backend/seq/EXU.scala 46:19]
  wire  alu_io_in_valid; // @[src/main/scala/nutcore/backend/seq/EXU.scala 46:19]
  wire [63:0] alu_io_in_bits_src1; // @[src/main/scala/nutcore/backend/seq/EXU.scala 46:19]
  wire [63:0] alu_io_in_bits_src2; // @[src/main/scala/nutcore/backend/seq/EXU.scala 46:19]
  wire [6:0] alu_io_in_bits_func; // @[src/main/scala/nutcore/backend/seq/EXU.scala 46:19]
  wire  alu_io_out_ready; // @[src/main/scala/nutcore/backend/seq/EXU.scala 46:19]
  wire  alu_io_out_valid; // @[src/main/scala/nutcore/backend/seq/EXU.scala 46:19]
  wire [63:0] alu_io_out_bits; // @[src/main/scala/nutcore/backend/seq/EXU.scala 46:19]
  wire [63:0] alu_io_cfIn_instr; // @[src/main/scala/nutcore/backend/seq/EXU.scala 46:19]
  wire [38:0] alu_io_cfIn_pc; // @[src/main/scala/nutcore/backend/seq/EXU.scala 46:19]
  wire [38:0] alu_io_cfIn_pnpc; // @[src/main/scala/nutcore/backend/seq/EXU.scala 46:19]
  wire [3:0] alu_io_cfIn_brIdx; // @[src/main/scala/nutcore/backend/seq/EXU.scala 46:19]
  wire [38:0] alu_io_redirect_target; // @[src/main/scala/nutcore/backend/seq/EXU.scala 46:19]
  wire  alu_io_redirect_valid; // @[src/main/scala/nutcore/backend/seq/EXU.scala 46:19]
  wire [63:0] alu_io_offset; // @[src/main/scala/nutcore/backend/seq/EXU.scala 46:19]
  wire  alu__WIRE_2_0; // @[src/main/scala/nutcore/backend/seq/EXU.scala 46:19]
  wire  alu_REG_0_valid; // @[src/main/scala/nutcore/backend/seq/EXU.scala 46:19]
  wire [38:0] alu_REG_0_pc; // @[src/main/scala/nutcore/backend/seq/EXU.scala 46:19]
  wire  alu_REG_0_isMissPredict; // @[src/main/scala/nutcore/backend/seq/EXU.scala 46:19]
  wire [38:0] alu_REG_0_actualTarget; // @[src/main/scala/nutcore/backend/seq/EXU.scala 46:19]
  wire  alu_REG_0_actualTaken; // @[src/main/scala/nutcore/backend/seq/EXU.scala 46:19]
  wire [6:0] alu_REG_0_fuOpType; // @[src/main/scala/nutcore/backend/seq/EXU.scala 46:19]
  wire [1:0] alu_REG_0_btbType; // @[src/main/scala/nutcore/backend/seq/EXU.scala 46:19]
  wire  alu_REG_0_isRVC; // @[src/main/scala/nutcore/backend/seq/EXU.scala 46:19]
  wire  alu__WIRE_15_0; // @[src/main/scala/nutcore/backend/seq/EXU.scala 46:19]
  wire  alu_DISPLAY_ENABLE; // @[src/main/scala/nutcore/backend/seq/EXU.scala 46:19]
  wire  alu__WIRE_13_0; // @[src/main/scala/nutcore/backend/seq/EXU.scala 46:19]
  wire  alu__WIRE_6_0; // @[src/main/scala/nutcore/backend/seq/EXU.scala 46:19]
  wire  alu__WIRE_5_0; // @[src/main/scala/nutcore/backend/seq/EXU.scala 46:19]
  wire  alu__WIRE_4_1; // @[src/main/scala/nutcore/backend/seq/EXU.scala 46:19]
  wire  alu__WIRE_3_0; // @[src/main/scala/nutcore/backend/seq/EXU.scala 46:19]
  wire  alu__WIRE_10_0; // @[src/main/scala/nutcore/backend/seq/EXU.scala 46:19]
  wire  alu__WIRE_9_0; // @[src/main/scala/nutcore/backend/seq/EXU.scala 46:19]
  wire  alu__WIRE_8_0; // @[src/main/scala/nutcore/backend/seq/EXU.scala 46:19]
  wire  alu__WIRE_7_0; // @[src/main/scala/nutcore/backend/seq/EXU.scala 46:19]
  wire  alu__WIRE_1_2; // @[src/main/scala/nutcore/backend/seq/EXU.scala 46:19]
  wire  alu__WIRE_12_0; // @[src/main/scala/nutcore/backend/seq/EXU.scala 46:19]
  wire  alu__WIRE_14_0; // @[src/main/scala/nutcore/backend/seq/EXU.scala 46:19]
  wire  alu__WIRE_11_0; // @[src/main/scala/nutcore/backend/seq/EXU.scala 46:19]
  wire  alu__WIRE_16_0; // @[src/main/scala/nutcore/backend/seq/EXU.scala 46:19]
  wire  lsu_clock; // @[src/main/scala/nutcore/backend/seq/EXU.scala 54:19]
  wire  lsu_reset; // @[src/main/scala/nutcore/backend/seq/EXU.scala 54:19]
  wire  lsu_io__in_ready; // @[src/main/scala/nutcore/backend/seq/EXU.scala 54:19]
  wire  lsu_io__in_valid; // @[src/main/scala/nutcore/backend/seq/EXU.scala 54:19]
  wire [63:0] lsu_io__in_bits_src1; // @[src/main/scala/nutcore/backend/seq/EXU.scala 54:19]
  wire [63:0] lsu_io__in_bits_src2; // @[src/main/scala/nutcore/backend/seq/EXU.scala 54:19]
  wire [6:0] lsu_io__in_bits_func; // @[src/main/scala/nutcore/backend/seq/EXU.scala 54:19]
  wire  lsu_io__out_ready; // @[src/main/scala/nutcore/backend/seq/EXU.scala 54:19]
  wire  lsu_io__out_valid; // @[src/main/scala/nutcore/backend/seq/EXU.scala 54:19]
  wire [63:0] lsu_io__out_bits; // @[src/main/scala/nutcore/backend/seq/EXU.scala 54:19]
  wire [63:0] lsu_io__wdata; // @[src/main/scala/nutcore/backend/seq/EXU.scala 54:19]
  wire [31:0] lsu_io__instr; // @[src/main/scala/nutcore/backend/seq/EXU.scala 54:19]
  wire  lsu_io__dmem_req_ready; // @[src/main/scala/nutcore/backend/seq/EXU.scala 54:19]
  wire  lsu_io__dmem_req_valid; // @[src/main/scala/nutcore/backend/seq/EXU.scala 54:19]
  wire [38:0] lsu_io__dmem_req_bits_addr; // @[src/main/scala/nutcore/backend/seq/EXU.scala 54:19]
  wire [2:0] lsu_io__dmem_req_bits_size; // @[src/main/scala/nutcore/backend/seq/EXU.scala 54:19]
  wire [3:0] lsu_io__dmem_req_bits_cmd; // @[src/main/scala/nutcore/backend/seq/EXU.scala 54:19]
  wire [7:0] lsu_io__dmem_req_bits_wmask; // @[src/main/scala/nutcore/backend/seq/EXU.scala 54:19]
  wire [63:0] lsu_io__dmem_req_bits_wdata; // @[src/main/scala/nutcore/backend/seq/EXU.scala 54:19]
  wire  lsu_io__dmem_resp_valid; // @[src/main/scala/nutcore/backend/seq/EXU.scala 54:19]
  wire [63:0] lsu_io__dmem_resp_bits_rdata; // @[src/main/scala/nutcore/backend/seq/EXU.scala 54:19]
  wire  lsu_io__isMMIO; // @[src/main/scala/nutcore/backend/seq/EXU.scala 54:19]
  wire  lsu_io__dtlbPF; // @[src/main/scala/nutcore/backend/seq/EXU.scala 54:19]
  wire  lsu_io__loadAddrMisaligned; // @[src/main/scala/nutcore/backend/seq/EXU.scala 54:19]
  wire  lsu_io__storeAddrMisaligned; // @[src/main/scala/nutcore/backend/seq/EXU.scala 54:19]
  wire  lsu_setLr_0; // @[src/main/scala/nutcore/backend/seq/EXU.scala 54:19]
  wire  lsu_lr_0; // @[src/main/scala/nutcore/backend/seq/EXU.scala 54:19]
  wire  lsu__WIRE_4; // @[src/main/scala/nutcore/backend/seq/EXU.scala 54:19]
  wire [63:0] lsu_lr_addr; // @[src/main/scala/nutcore/backend/seq/EXU.scala 54:19]
  wire  lsu_io_isMMIO; // @[src/main/scala/nutcore/backend/seq/EXU.scala 54:19]
  wire  lsu_DISPLAY_ENABLE; // @[src/main/scala/nutcore/backend/seq/EXU.scala 54:19]
  wire  lsu_DTLBPF; // @[src/main/scala/nutcore/backend/seq/EXU.scala 54:19]
  wire  lsu_r; // @[src/main/scala/nutcore/backend/seq/EXU.scala 54:19]
  wire  lsu_setLrVal_0; // @[src/main/scala/nutcore/backend/seq/EXU.scala 54:19]
  wire [63:0] lsu_io_in_bits_src1; // @[src/main/scala/nutcore/backend/seq/EXU.scala 54:19]
  wire  lsu_DTLBENABLE; // @[src/main/scala/nutcore/backend/seq/EXU.scala 54:19]
  wire  lsu_DTLBFINISH; // @[src/main/scala/nutcore/backend/seq/EXU.scala 54:19]
  wire  lsu_r_1; // @[src/main/scala/nutcore/backend/seq/EXU.scala 54:19]
  wire  lsu_lsuMMIO_0; // @[src/main/scala/nutcore/backend/seq/EXU.scala 54:19]
  wire  lsu__WIRE_16; // @[src/main/scala/nutcore/backend/seq/EXU.scala 54:19]
  wire [63:0] lsu_setLrAddr_0; // @[src/main/scala/nutcore/backend/seq/EXU.scala 54:19]
  wire  mdu_clock; // @[src/main/scala/nutcore/backend/seq/EXU.scala 63:19]
  wire  mdu_reset; // @[src/main/scala/nutcore/backend/seq/EXU.scala 63:19]
  wire  mdu_io_in_ready; // @[src/main/scala/nutcore/backend/seq/EXU.scala 63:19]
  wire  mdu_io_in_valid; // @[src/main/scala/nutcore/backend/seq/EXU.scala 63:19]
  wire [63:0] mdu_io_in_bits_src1; // @[src/main/scala/nutcore/backend/seq/EXU.scala 63:19]
  wire [63:0] mdu_io_in_bits_src2; // @[src/main/scala/nutcore/backend/seq/EXU.scala 63:19]
  wire [6:0] mdu_io_in_bits_func; // @[src/main/scala/nutcore/backend/seq/EXU.scala 63:19]
  wire  mdu_io_out_ready; // @[src/main/scala/nutcore/backend/seq/EXU.scala 63:19]
  wire  mdu_io_out_valid; // @[src/main/scala/nutcore/backend/seq/EXU.scala 63:19]
  wire [63:0] mdu_io_out_bits; // @[src/main/scala/nutcore/backend/seq/EXU.scala 63:19]
  wire  mdu__WIRE_0; // @[src/main/scala/nutcore/backend/seq/EXU.scala 63:19]
  wire  mdu_DISPLAY_ENABLE; // @[src/main/scala/nutcore/backend/seq/EXU.scala 63:19]
  wire  csr_clock; // @[src/main/scala/nutcore/backend/seq/EXU.scala 68:19]
  wire  csr_reset; // @[src/main/scala/nutcore/backend/seq/EXU.scala 68:19]
  wire  csr_io_in_valid; // @[src/main/scala/nutcore/backend/seq/EXU.scala 68:19]
  wire [63:0] csr_io_in_bits_src1; // @[src/main/scala/nutcore/backend/seq/EXU.scala 68:19]
  wire [63:0] csr_io_in_bits_src2; // @[src/main/scala/nutcore/backend/seq/EXU.scala 68:19]
  wire [6:0] csr_io_in_bits_func; // @[src/main/scala/nutcore/backend/seq/EXU.scala 68:19]
  wire  csr_io_out_ready; // @[src/main/scala/nutcore/backend/seq/EXU.scala 68:19]
  wire  csr_io_out_valid; // @[src/main/scala/nutcore/backend/seq/EXU.scala 68:19]
  wire [63:0] csr_io_out_bits; // @[src/main/scala/nutcore/backend/seq/EXU.scala 68:19]
  wire [63:0] csr_io_cfIn_instr; // @[src/main/scala/nutcore/backend/seq/EXU.scala 68:19]
  wire [38:0] csr_io_cfIn_pc; // @[src/main/scala/nutcore/backend/seq/EXU.scala 68:19]
  wire  csr_io_cfIn_exceptionVec_1; // @[src/main/scala/nutcore/backend/seq/EXU.scala 68:19]
  wire  csr_io_cfIn_exceptionVec_2; // @[src/main/scala/nutcore/backend/seq/EXU.scala 68:19]
  wire  csr_io_cfIn_exceptionVec_4; // @[src/main/scala/nutcore/backend/seq/EXU.scala 68:19]
  wire  csr_io_cfIn_exceptionVec_6; // @[src/main/scala/nutcore/backend/seq/EXU.scala 68:19]
  wire  csr_io_cfIn_exceptionVec_12; // @[src/main/scala/nutcore/backend/seq/EXU.scala 68:19]
  wire  csr_io_cfIn_intrVec_0; // @[src/main/scala/nutcore/backend/seq/EXU.scala 68:19]
  wire  csr_io_cfIn_intrVec_1; // @[src/main/scala/nutcore/backend/seq/EXU.scala 68:19]
  wire  csr_io_cfIn_intrVec_2; // @[src/main/scala/nutcore/backend/seq/EXU.scala 68:19]
  wire  csr_io_cfIn_intrVec_3; // @[src/main/scala/nutcore/backend/seq/EXU.scala 68:19]
  wire  csr_io_cfIn_intrVec_4; // @[src/main/scala/nutcore/backend/seq/EXU.scala 68:19]
  wire  csr_io_cfIn_intrVec_5; // @[src/main/scala/nutcore/backend/seq/EXU.scala 68:19]
  wire  csr_io_cfIn_intrVec_6; // @[src/main/scala/nutcore/backend/seq/EXU.scala 68:19]
  wire  csr_io_cfIn_intrVec_7; // @[src/main/scala/nutcore/backend/seq/EXU.scala 68:19]
  wire  csr_io_cfIn_intrVec_8; // @[src/main/scala/nutcore/backend/seq/EXU.scala 68:19]
  wire  csr_io_cfIn_intrVec_9; // @[src/main/scala/nutcore/backend/seq/EXU.scala 68:19]
  wire  csr_io_cfIn_intrVec_10; // @[src/main/scala/nutcore/backend/seq/EXU.scala 68:19]
  wire  csr_io_cfIn_intrVec_11; // @[src/main/scala/nutcore/backend/seq/EXU.scala 68:19]
  wire  csr_io_cfIn_crossPageIPFFix; // @[src/main/scala/nutcore/backend/seq/EXU.scala 68:19]
  wire [38:0] csr_io_redirect_target; // @[src/main/scala/nutcore/backend/seq/EXU.scala 68:19]
  wire  csr_io_redirect_valid; // @[src/main/scala/nutcore/backend/seq/EXU.scala 68:19]
  wire  csr_io_instrValid; // @[src/main/scala/nutcore/backend/seq/EXU.scala 68:19]
  wire [63:0] csr_io_intrNO; // @[src/main/scala/nutcore/backend/seq/EXU.scala 68:19]
  wire [1:0] csr_io_imemMMU_priviledgeMode; // @[src/main/scala/nutcore/backend/seq/EXU.scala 68:19]
  wire [1:0] csr_io_dmemMMU_priviledgeMode; // @[src/main/scala/nutcore/backend/seq/EXU.scala 68:19]
  wire  csr_io_dmemMMU_status_sum; // @[src/main/scala/nutcore/backend/seq/EXU.scala 68:19]
  wire  csr_io_dmemMMU_status_mxr; // @[src/main/scala/nutcore/backend/seq/EXU.scala 68:19]
  wire  csr_io_dmemMMU_loadPF; // @[src/main/scala/nutcore/backend/seq/EXU.scala 68:19]
  wire  csr_io_dmemMMU_storePF; // @[src/main/scala/nutcore/backend/seq/EXU.scala 68:19]
  wire [38:0] csr_io_dmemMMU_addr; // @[src/main/scala/nutcore/backend/seq/EXU.scala 68:19]
  wire  csr_io_wenFix; // @[src/main/scala/nutcore/backend/seq/EXU.scala 68:19]
  wire  csr_set_lr; // @[src/main/scala/nutcore/backend/seq/EXU.scala 68:19]
  wire  csr_lr_0; // @[src/main/scala/nutcore/backend/seq/EXU.scala 68:19]
  wire  csr_MbpBWrong; // @[src/main/scala/nutcore/backend/seq/EXU.scala 68:19]
  wire  csr_perfCntCondMmulInstr; // @[src/main/scala/nutcore/backend/seq/EXU.scala 68:19]
  wire  csr_meip_0; // @[src/main/scala/nutcore/backend/seq/EXU.scala 68:19]
  wire  csr_perfCntCondMlsuInstr; // @[src/main/scala/nutcore/backend/seq/EXU.scala 68:19]
  wire [63:0] csr_lrAddr_0; // @[src/main/scala/nutcore/backend/seq/EXU.scala 68:19]
  wire  csr_perfCntCondMexuBusy; // @[src/main/scala/nutcore/backend/seq/EXU.scala 68:19]
  wire  csr_perfCntCondMmmioInstr; // @[src/main/scala/nutcore/backend/seq/EXU.scala 68:19]
  wire  csr_perfCntCondMaluInstr; // @[src/main/scala/nutcore/backend/seq/EXU.scala 68:19]
  wire  csr_MbpRRight; // @[src/main/scala/nutcore/backend/seq/EXU.scala 68:19]
  wire [63:0] csr_satp_0; // @[src/main/scala/nutcore/backend/seq/EXU.scala 68:19]
  wire  csr_DISPLAY_ENABLE; // @[src/main/scala/nutcore/backend/seq/EXU.scala 68:19]
  wire  csr_MbpIRight; // @[src/main/scala/nutcore/backend/seq/EXU.scala 68:19]
  wire  csr_perfCntCondMcsrInstr; // @[src/main/scala/nutcore/backend/seq/EXU.scala 68:19]
  wire  csr_Custom4; // @[src/main/scala/nutcore/backend/seq/EXU.scala 68:19]
  wire  csr_Custom3; // @[src/main/scala/nutcore/backend/seq/EXU.scala 68:19]
  wire  csr_perfCntCondMifuFlush; // @[src/main/scala/nutcore/backend/seq/EXU.scala 68:19]
  wire  csr_Custom2; // @[src/main/scala/nutcore/backend/seq/EXU.scala 68:19]
  wire  csr_Custom1; // @[src/main/scala/nutcore/backend/seq/EXU.scala 68:19]
  wire  csr_Custom8; // @[src/main/scala/nutcore/backend/seq/EXU.scala 68:19]
  wire  csr_Custom7; // @[src/main/scala/nutcore/backend/seq/EXU.scala 68:19]
  wire  csr_perfCntCondMrawStall; // @[src/main/scala/nutcore/backend/seq/EXU.scala 68:19]
  wire  csr_perfCntCondMloadStall; // @[src/main/scala/nutcore/backend/seq/EXU.scala 68:19]
  wire  csr_Custom6; // @[src/main/scala/nutcore/backend/seq/EXU.scala 68:19]
  wire  csr_Custom5; // @[src/main/scala/nutcore/backend/seq/EXU.scala 68:19]
  wire  csr_perfCntCondISUIssue; // @[src/main/scala/nutcore/backend/seq/EXU.scala 68:19]
  wire  csr_mtip_0; // @[src/main/scala/nutcore/backend/seq/EXU.scala 68:19]
  wire  csr_perfCntCondMultiCommit; // @[src/main/scala/nutcore/backend/seq/EXU.scala 68:19]
  wire  csr_MbpBRight; // @[src/main/scala/nutcore/backend/seq/EXU.scala 68:19]
  wire  csr_perfCntCondMbruInstr; // @[src/main/scala/nutcore/backend/seq/EXU.scala 68:19]
  wire  csr_set_lr_val; // @[src/main/scala/nutcore/backend/seq/EXU.scala 68:19]
  wire  csr_MbpJWrong; // @[src/main/scala/nutcore/backend/seq/EXU.scala 68:19]
  wire  csr_nutcoretrap_0; // @[src/main/scala/nutcore/backend/seq/EXU.scala 68:19]
  wire [63:0] csr_LSUADDR; // @[src/main/scala/nutcore/backend/seq/EXU.scala 68:19]
  wire [11:0] csr__WIRE_4; // @[src/main/scala/nutcore/backend/seq/EXU.scala 68:19]
  wire  csr_perfCntCondMstoreStall; // @[src/main/scala/nutcore/backend/seq/EXU.scala 68:19]
  wire  csr_MbpIWrong; // @[src/main/scala/nutcore/backend/seq/EXU.scala 68:19]
  wire  csr_MbpJRight; // @[src/main/scala/nutcore/backend/seq/EXU.scala 68:19]
  wire  csr_perfCntCondMloadInstr; // @[src/main/scala/nutcore/backend/seq/EXU.scala 68:19]
  wire  csr_perfCntCondMmduInstr; // @[src/main/scala/nutcore/backend/seq/EXU.scala 68:19]
  wire [63:0] csr_set_lr_addr; // @[src/main/scala/nutcore/backend/seq/EXU.scala 68:19]
  wire  csr_perfCntCondMimemStall; // @[src/main/scala/nutcore/backend/seq/EXU.scala 68:19]
  wire  csr_MbpRWrong; // @[src/main/scala/nutcore/backend/seq/EXU.scala 68:19]
  wire  csr_msip_0; // @[src/main/scala/nutcore/backend/seq/EXU.scala 68:19]
  wire  csr_perfCntCondMinstret; // @[src/main/scala/nutcore/backend/seq/EXU.scala 68:19]
  wire  mou_clock; // @[src/main/scala/nutcore/backend/seq/EXU.scala 82:19]
  wire  mou_reset; // @[src/main/scala/nutcore/backend/seq/EXU.scala 82:19]
  wire  mou_io_in_valid; // @[src/main/scala/nutcore/backend/seq/EXU.scala 82:19]
  wire [6:0] mou_io_in_bits_func; // @[src/main/scala/nutcore/backend/seq/EXU.scala 82:19]
  wire [38:0] mou_io_cfIn_pc; // @[src/main/scala/nutcore/backend/seq/EXU.scala 82:19]
  wire [38:0] mou_io_redirect_target; // @[src/main/scala/nutcore/backend/seq/EXU.scala 82:19]
  wire  mou_io_redirect_valid; // @[src/main/scala/nutcore/backend/seq/EXU.scala 82:19]
  wire  mou_DISPLAY_ENABLE; // @[src/main/scala/nutcore/backend/seq/EXU.scala 82:19]
  wire  mou__WIRE_11; // @[src/main/scala/nutcore/backend/seq/EXU.scala 82:19]
  wire  mou__WIRE_1_4; // @[src/main/scala/nutcore/backend/seq/EXU.scala 82:19]
  wire  _fuValids_0_T_2 = ~io__flush; // @[src/main/scala/nutcore/backend/seq/EXU.scala 44:84]
  wire  fuValids_1 = io__in_bits_ctrl_fuType == 3'h1 & io__in_valid & ~io__flush; // @[src/main/scala/nutcore/backend/seq/EXU.scala 44:81]
  wire  fuValids_3 = io__in_bits_ctrl_fuType == 3'h3 & io__in_valid & ~io__flush; // @[src/main/scala/nutcore/backend/seq/EXU.scala 44:81]
  wire [38:0] _io_out_bits_isMMIO_T = io__in_bits_cf_pc ^ 39'h30000000; // @[src/main/scala/nutcore/NutCore.scala 87:11]
  wire  _io_out_bits_isMMIO_T_2 = _io_out_bits_isMMIO_T[31:28] == 4'h0; // @[src/main/scala/nutcore/NutCore.scala 87:44]
  wire [38:0] _io_out_bits_isMMIO_T_3 = io__in_bits_cf_pc ^ 39'h40000000; // @[src/main/scala/nutcore/NutCore.scala 87:11]
  wire  _io_out_bits_isMMIO_T_5 = _io_out_bits_isMMIO_T_3[31:30] == 2'h0; // @[src/main/scala/nutcore/NutCore.scala 87:44]
  wire  _io_out_bits_isMMIO_T_6 = _io_out_bits_isMMIO_T_2 | _io_out_bits_isMMIO_T_5; // @[src/main/scala/nutcore/NutCore.scala 88:15]
  wire  lsuTlbPF = lsu_io__dtlbPF; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 44:12 src/main/scala/nutcore/backend/seq/EXU.scala 55:26]
  wire [38:0] _io_out_bits_decode_cf_redirect_T_target = csr_io_redirect_valid ? csr_io_redirect_target :
    alu_io_redirect_target; // @[src/main/scala/nutcore/backend/seq/EXU.scala 100:10]
  wire  _io_out_bits_decode_cf_redirect_T_valid = csr_io_redirect_valid ? csr_io_redirect_valid : alu_io_redirect_valid; // @[src/main/scala/nutcore/backend/seq/EXU.scala 100:10]
  wire  _T_1 = mou_io_redirect_valid | csr_io_redirect_valid | alu_io_redirect_valid; // @[src/main/scala/nutcore/backend/seq/EXU.scala 102:56]
  reg [63:0] c; // @[src/main/scala/utils/GTimer.scala 24:20]
  wire [63:0] _c_T_1 = c + 64'h1; // @[src/main/scala/utils/GTimer.scala 25:12]
  wire  _T_2 = _T_1 & DISPLAY_ENABLE; // @[src/main/scala/utils/Debug.scala 55:16]
  wire  _T_4 = ~reset; // @[src/main/scala/utils/Debug.scala 56:24]
  reg [63:0] c_1; // @[src/main/scala/utils/GTimer.scala 24:20]
  wire [63:0] _c_T_3 = c_1 + 64'h1; // @[src/main/scala/utils/GTimer.scala 25:12]
  wire  _io_out_valid_T_1 = 3'h1 == io__in_bits_ctrl_fuType ? lsu_io__out_valid : 1'h1; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _io_out_valid_T_3 = 3'h2 == io__in_bits_ctrl_fuType ? mdu_io_out_valid : _io_out_valid_T_1; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _io_forward_wb_rfData_T = alu_io_out_ready & alu_io_out_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  wire  isBru = io__in_bits_ctrl_fuOpType[4]; // @[src/main/scala/nutcore/backend/fu/ALU.scala 62:31]
  wire  _WIRE_3 = mdu_io_out_ready & mdu_io_out_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  wire  nutcoretrap = io__in_bits_ctrl_isNutCoreTrap & io__in_valid; // @[src/main/scala/nutcore/backend/seq/EXU.scala 135:62]
  wire  _WIRE_1 = _io_forward_wb_rfData_T & isBru; // @[src/main/scala/nutcore/backend/seq/EXU.scala 127:50]
  wire  _WIRE_4 = csr_io_out_ready & csr_io_out_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  wire  _WIRE = _io_forward_wb_rfData_T & ~isBru; // @[src/main/scala/nutcore/backend/seq/EXU.scala 126:50]
  wire  _WIRE_2 = lsu_io__out_ready & lsu_io__out_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  ALU alu ( // @[src/main/scala/nutcore/backend/seq/EXU.scala 46:19]
    .clock(alu_clock),
    .reset(alu_reset),
    .io_in_valid(alu_io_in_valid),
    .io_in_bits_src1(alu_io_in_bits_src1),
    .io_in_bits_src2(alu_io_in_bits_src2),
    .io_in_bits_func(alu_io_in_bits_func),
    .io_out_ready(alu_io_out_ready),
    .io_out_valid(alu_io_out_valid),
    .io_out_bits(alu_io_out_bits),
    .io_cfIn_instr(alu_io_cfIn_instr),
    .io_cfIn_pc(alu_io_cfIn_pc),
    .io_cfIn_pnpc(alu_io_cfIn_pnpc),
    .io_cfIn_brIdx(alu_io_cfIn_brIdx),
    .io_redirect_target(alu_io_redirect_target),
    .io_redirect_valid(alu_io_redirect_valid),
    .io_offset(alu_io_offset),
    ._WIRE_2_0(alu__WIRE_2_0),
    .REG_0_valid(alu_REG_0_valid),
    .REG_0_pc(alu_REG_0_pc),
    .REG_0_isMissPredict(alu_REG_0_isMissPredict),
    .REG_0_actualTarget(alu_REG_0_actualTarget),
    .REG_0_actualTaken(alu_REG_0_actualTaken),
    .REG_0_fuOpType(alu_REG_0_fuOpType),
    .REG_0_btbType(alu_REG_0_btbType),
    .REG_0_isRVC(alu_REG_0_isRVC),
    ._WIRE_15_0(alu__WIRE_15_0),
    .DISPLAY_ENABLE(alu_DISPLAY_ENABLE),
    ._WIRE_13_0(alu__WIRE_13_0),
    ._WIRE_6_0(alu__WIRE_6_0),
    ._WIRE_5_0(alu__WIRE_5_0),
    ._WIRE_4_1(alu__WIRE_4_1),
    ._WIRE_3_0(alu__WIRE_3_0),
    ._WIRE_10_0(alu__WIRE_10_0),
    ._WIRE_9_0(alu__WIRE_9_0),
    ._WIRE_8_0(alu__WIRE_8_0),
    ._WIRE_7_0(alu__WIRE_7_0),
    ._WIRE_1_2(alu__WIRE_1_2),
    ._WIRE_12_0(alu__WIRE_12_0),
    ._WIRE_14_0(alu__WIRE_14_0),
    ._WIRE_11_0(alu__WIRE_11_0),
    ._WIRE_16_0(alu__WIRE_16_0)
  );
  UnpipelinedLSU lsu ( // @[src/main/scala/nutcore/backend/seq/EXU.scala 54:19]
    .clock(lsu_clock),
    .reset(lsu_reset),
    .io__in_ready(lsu_io__in_ready),
    .io__in_valid(lsu_io__in_valid),
    .io__in_bits_src1(lsu_io__in_bits_src1),
    .io__in_bits_src2(lsu_io__in_bits_src2),
    .io__in_bits_func(lsu_io__in_bits_func),
    .io__out_ready(lsu_io__out_ready),
    .io__out_valid(lsu_io__out_valid),
    .io__out_bits(lsu_io__out_bits),
    .io__wdata(lsu_io__wdata),
    .io__instr(lsu_io__instr),
    .io__dmem_req_ready(lsu_io__dmem_req_ready),
    .io__dmem_req_valid(lsu_io__dmem_req_valid),
    .io__dmem_req_bits_addr(lsu_io__dmem_req_bits_addr),
    .io__dmem_req_bits_size(lsu_io__dmem_req_bits_size),
    .io__dmem_req_bits_cmd(lsu_io__dmem_req_bits_cmd),
    .io__dmem_req_bits_wmask(lsu_io__dmem_req_bits_wmask),
    .io__dmem_req_bits_wdata(lsu_io__dmem_req_bits_wdata),
    .io__dmem_resp_valid(lsu_io__dmem_resp_valid),
    .io__dmem_resp_bits_rdata(lsu_io__dmem_resp_bits_rdata),
    .io__isMMIO(lsu_io__isMMIO),
    .io__dtlbPF(lsu_io__dtlbPF),
    .io__loadAddrMisaligned(lsu_io__loadAddrMisaligned),
    .io__storeAddrMisaligned(lsu_io__storeAddrMisaligned),
    .setLr_0(lsu_setLr_0),
    .lr_0(lsu_lr_0),
    ._WIRE_4(lsu__WIRE_4),
    .lr_addr(lsu_lr_addr),
    .io_isMMIO(lsu_io_isMMIO),
    .DISPLAY_ENABLE(lsu_DISPLAY_ENABLE),
    .DTLBPF(lsu_DTLBPF),
    .r(lsu_r),
    .setLrVal_0(lsu_setLrVal_0),
    .io_in_bits_src1(lsu_io_in_bits_src1),
    .DTLBENABLE(lsu_DTLBENABLE),
    .DTLBFINISH(lsu_DTLBFINISH),
    .r_1(lsu_r_1),
    .lsuMMIO_0(lsu_lsuMMIO_0),
    ._WIRE_16(lsu__WIRE_16),
    .setLrAddr_0(lsu_setLrAddr_0)
  );
  MDU mdu ( // @[src/main/scala/nutcore/backend/seq/EXU.scala 63:19]
    .clock(mdu_clock),
    .reset(mdu_reset),
    .io_in_ready(mdu_io_in_ready),
    .io_in_valid(mdu_io_in_valid),
    .io_in_bits_src1(mdu_io_in_bits_src1),
    .io_in_bits_src2(mdu_io_in_bits_src2),
    .io_in_bits_func(mdu_io_in_bits_func),
    .io_out_ready(mdu_io_out_ready),
    .io_out_valid(mdu_io_out_valid),
    .io_out_bits(mdu_io_out_bits),
    ._WIRE_0(mdu__WIRE_0),
    .DISPLAY_ENABLE(mdu_DISPLAY_ENABLE)
  );
  CSR csr ( // @[src/main/scala/nutcore/backend/seq/EXU.scala 68:19]
    .clock(csr_clock),
    .reset(csr_reset),
    .io_in_valid(csr_io_in_valid),
    .io_in_bits_src1(csr_io_in_bits_src1),
    .io_in_bits_src2(csr_io_in_bits_src2),
    .io_in_bits_func(csr_io_in_bits_func),
    .io_out_ready(csr_io_out_ready),
    .io_out_valid(csr_io_out_valid),
    .io_out_bits(csr_io_out_bits),
    .io_cfIn_instr(csr_io_cfIn_instr),
    .io_cfIn_pc(csr_io_cfIn_pc),
    .io_cfIn_exceptionVec_1(csr_io_cfIn_exceptionVec_1),
    .io_cfIn_exceptionVec_2(csr_io_cfIn_exceptionVec_2),
    .io_cfIn_exceptionVec_4(csr_io_cfIn_exceptionVec_4),
    .io_cfIn_exceptionVec_6(csr_io_cfIn_exceptionVec_6),
    .io_cfIn_exceptionVec_12(csr_io_cfIn_exceptionVec_12),
    .io_cfIn_intrVec_0(csr_io_cfIn_intrVec_0),
    .io_cfIn_intrVec_1(csr_io_cfIn_intrVec_1),
    .io_cfIn_intrVec_2(csr_io_cfIn_intrVec_2),
    .io_cfIn_intrVec_3(csr_io_cfIn_intrVec_3),
    .io_cfIn_intrVec_4(csr_io_cfIn_intrVec_4),
    .io_cfIn_intrVec_5(csr_io_cfIn_intrVec_5),
    .io_cfIn_intrVec_6(csr_io_cfIn_intrVec_6),
    .io_cfIn_intrVec_7(csr_io_cfIn_intrVec_7),
    .io_cfIn_intrVec_8(csr_io_cfIn_intrVec_8),
    .io_cfIn_intrVec_9(csr_io_cfIn_intrVec_9),
    .io_cfIn_intrVec_10(csr_io_cfIn_intrVec_10),
    .io_cfIn_intrVec_11(csr_io_cfIn_intrVec_11),
    .io_cfIn_crossPageIPFFix(csr_io_cfIn_crossPageIPFFix),
    .io_redirect_target(csr_io_redirect_target),
    .io_redirect_valid(csr_io_redirect_valid),
    .io_instrValid(csr_io_instrValid),
    .io_intrNO(csr_io_intrNO),
    .io_imemMMU_priviledgeMode(csr_io_imemMMU_priviledgeMode),
    .io_dmemMMU_priviledgeMode(csr_io_dmemMMU_priviledgeMode),
    .io_dmemMMU_status_sum(csr_io_dmemMMU_status_sum),
    .io_dmemMMU_status_mxr(csr_io_dmemMMU_status_mxr),
    .io_dmemMMU_loadPF(csr_io_dmemMMU_loadPF),
    .io_dmemMMU_storePF(csr_io_dmemMMU_storePF),
    .io_dmemMMU_addr(csr_io_dmemMMU_addr),
    .io_wenFix(csr_io_wenFix),
    .set_lr(csr_set_lr),
    .lr_0(csr_lr_0),
    .MbpBWrong(csr_MbpBWrong),
    .perfCntCondMmulInstr(csr_perfCntCondMmulInstr),
    .meip_0(csr_meip_0),
    .perfCntCondMlsuInstr(csr_perfCntCondMlsuInstr),
    .lrAddr_0(csr_lrAddr_0),
    .perfCntCondMexuBusy(csr_perfCntCondMexuBusy),
    .perfCntCondMmmioInstr(csr_perfCntCondMmmioInstr),
    .perfCntCondMaluInstr(csr_perfCntCondMaluInstr),
    .MbpRRight(csr_MbpRRight),
    .satp_0(csr_satp_0),
    .DISPLAY_ENABLE(csr_DISPLAY_ENABLE),
    .MbpIRight(csr_MbpIRight),
    .perfCntCondMcsrInstr(csr_perfCntCondMcsrInstr),
    .Custom4(csr_Custom4),
    .Custom3(csr_Custom3),
    .perfCntCondMifuFlush(csr_perfCntCondMifuFlush),
    .Custom2(csr_Custom2),
    .Custom1(csr_Custom1),
    .Custom8(csr_Custom8),
    .Custom7(csr_Custom7),
    .perfCntCondMrawStall(csr_perfCntCondMrawStall),
    .perfCntCondMloadStall(csr_perfCntCondMloadStall),
    .Custom6(csr_Custom6),
    .Custom5(csr_Custom5),
    .perfCntCondISUIssue(csr_perfCntCondISUIssue),
    .mtip_0(csr_mtip_0),
    .perfCntCondMultiCommit(csr_perfCntCondMultiCommit),
    .MbpBRight(csr_MbpBRight),
    .perfCntCondMbruInstr(csr_perfCntCondMbruInstr),
    .set_lr_val(csr_set_lr_val),
    .MbpJWrong(csr_MbpJWrong),
    .nutcoretrap_0(csr_nutcoretrap_0),
    .LSUADDR(csr_LSUADDR),
    ._WIRE_4(csr__WIRE_4),
    .perfCntCondMstoreStall(csr_perfCntCondMstoreStall),
    .MbpIWrong(csr_MbpIWrong),
    .MbpJRight(csr_MbpJRight),
    .perfCntCondMloadInstr(csr_perfCntCondMloadInstr),
    .perfCntCondMmduInstr(csr_perfCntCondMmduInstr),
    .set_lr_addr(csr_set_lr_addr),
    .perfCntCondMimemStall(csr_perfCntCondMimemStall),
    .MbpRWrong(csr_MbpRWrong),
    .msip_0(csr_msip_0),
    .perfCntCondMinstret(csr_perfCntCondMinstret)
  );
  MOU mou ( // @[src/main/scala/nutcore/backend/seq/EXU.scala 82:19]
    .clock(mou_clock),
    .reset(mou_reset),
    .io_in_valid(mou_io_in_valid),
    .io_in_bits_func(mou_io_in_bits_func),
    .io_cfIn_pc(mou_io_cfIn_pc),
    .io_redirect_target(mou_io_redirect_target),
    .io_redirect_valid(mou_io_redirect_valid),
    .DISPLAY_ENABLE(mou_DISPLAY_ENABLE),
    ._WIRE_11(mou__WIRE_11),
    ._WIRE_1_4(mou__WIRE_1_4)
  );
  assign io__in_ready = ~io__in_valid | io__out_valid; // @[src/main/scala/nutcore/backend/seq/EXU.scala 117:31]
  assign io__out_valid = io__in_valid & _io_out_valid_T_3; // @[src/main/scala/nutcore/backend/seq/EXU.scala 106:31]
  assign io__out_bits_decode_cf_instr = io__in_bits_cf_instr; // @[src/main/scala/nutcore/backend/seq/EXU.scala 95:31]
  assign io__out_bits_decode_cf_pc = io__in_bits_cf_pc; // @[src/main/scala/nutcore/backend/seq/EXU.scala 94:28]
  assign io__out_bits_decode_cf_redirect_target = mou_io_redirect_valid ? mou_io_redirect_target :
    _io_out_bits_decode_cf_redirect_T_target; // @[src/main/scala/nutcore/backend/seq/EXU.scala 99:8]
  assign io__out_bits_decode_cf_redirect_valid = mou_io_redirect_valid ? mou_io_redirect_valid :
    _io_out_bits_decode_cf_redirect_T_valid; // @[src/main/scala/nutcore/backend/seq/EXU.scala 99:8]
  assign io__out_bits_decode_ctrl_fuType = io__in_bits_ctrl_fuType; // @[src/main/scala/nutcore/backend/seq/EXU.scala 92:14]
  assign io__out_bits_decode_ctrl_rfWen = io__in_bits_ctrl_rfWen & (~lsuTlbPF & ~lsu_io__loadAddrMisaligned & ~
    lsu_io__storeAddrMisaligned | ~fuValids_1) & ~(csr_io_wenFix & fuValids_3); // @[src/main/scala/nutcore/backend/seq/EXU.scala 90:125]
  assign io__out_bits_decode_ctrl_rfDest = io__in_bits_ctrl_rfDest; // @[src/main/scala/nutcore/backend/seq/EXU.scala 91:14]
  assign io__out_bits_isMMIO = lsu_io__isMMIO | _io_out_bits_isMMIO_T_6 & io__out_valid; // @[src/main/scala/nutcore/backend/seq/EXU.scala 59:39]
  assign io__out_bits_intrNO = csr_io_intrNO; // @[src/main/scala/nutcore/backend/seq/EXU.scala 75:22]
  assign io__out_bits_commits_0 = alu_io_out_bits; // @[src/main/scala/nutcore/backend/seq/EXU.scala 111:35]
  assign io__out_bits_commits_1 = lsu_io__out_bits; // @[src/main/scala/nutcore/backend/seq/EXU.scala 112:35]
  assign io__out_bits_commits_2 = mdu_io_out_bits; // @[src/main/scala/nutcore/backend/seq/EXU.scala 114:35]
  assign io__out_bits_commits_3 = csr_io_out_bits; // @[src/main/scala/nutcore/backend/seq/EXU.scala 113:35]
  assign io__dmem_req_valid = lsu_io__dmem_req_valid; // @[src/main/scala/nutcore/backend/seq/EXU.scala 60:11]
  assign io__dmem_req_bits_addr = lsu_io__dmem_req_bits_addr; // @[src/main/scala/nutcore/backend/seq/EXU.scala 60:11]
  assign io__dmem_req_bits_size = lsu_io__dmem_req_bits_size; // @[src/main/scala/nutcore/backend/seq/EXU.scala 60:11]
  assign io__dmem_req_bits_cmd = lsu_io__dmem_req_bits_cmd; // @[src/main/scala/nutcore/backend/seq/EXU.scala 60:11]
  assign io__dmem_req_bits_wmask = lsu_io__dmem_req_bits_wmask; // @[src/main/scala/nutcore/backend/seq/EXU.scala 60:11]
  assign io__dmem_req_bits_wdata = lsu_io__dmem_req_bits_wdata; // @[src/main/scala/nutcore/backend/seq/EXU.scala 60:11]
  assign io__forward_valid = io__in_valid; // @[src/main/scala/nutcore/backend/seq/EXU.scala 119:20]
  assign io__forward_wb_rfWen = io__in_bits_ctrl_rfWen; // @[src/main/scala/nutcore/backend/seq/EXU.scala 120:23]
  assign io__forward_wb_rfDest = io__in_bits_ctrl_rfDest; // @[src/main/scala/nutcore/backend/seq/EXU.scala 121:24]
  assign io__forward_wb_rfData = _io_forward_wb_rfData_T ? alu_io_out_bits : lsu_io__out_bits; // @[src/main/scala/nutcore/backend/seq/EXU.scala 122:30]
  assign io__forward_fuType = io__in_bits_ctrl_fuType; // @[src/main/scala/nutcore/backend/seq/EXU.scala 123:21]
  assign io__memMMU_imem_priviledgeMode = csr_io_imemMMU_priviledgeMode; // @[src/main/scala/nutcore/backend/seq/EXU.scala 79:18]
  assign io__memMMU_dmem_priviledgeMode = csr_io_dmemMMU_priviledgeMode; // @[src/main/scala/nutcore/backend/seq/EXU.scala 80:18]
  assign io__memMMU_dmem_status_sum = csr_io_dmemMMU_status_sum; // @[src/main/scala/nutcore/backend/seq/EXU.scala 80:18]
  assign io__memMMU_dmem_status_mxr = csr_io_dmemMMU_status_mxr; // @[src/main/scala/nutcore/backend/seq/EXU.scala 80:18]
  assign REG_valid = alu_REG_0_valid;
  assign REG_pc = alu_REG_0_pc;
  assign REG_isMissPredict = alu_REG_0_isMissPredict;
  assign REG_actualTarget = alu_REG_0_actualTarget;
  assign REG_actualTaken = alu_REG_0_actualTaken;
  assign REG_fuOpType = alu_REG_0_fuOpType;
  assign REG_btbType = alu_REG_0_btbType;
  assign REG_isRVC = alu_REG_0_isRVC;
  assign _WIRE_6 = lsu__WIRE_4;
  assign satp = csr_satp_0;
  assign _WIRE_12 = mou__WIRE_11;
  assign _WIRE_1_4 = mou__WIRE_1_4;
  assign _WIRE_14 = csr__WIRE_4;
  assign alu_clock = clock;
  assign alu_reset = reset;
  assign alu_io_in_valid = io__in_bits_ctrl_fuType == 3'h0 & io__in_valid & ~io__flush; // @[src/main/scala/nutcore/backend/seq/EXU.scala 44:81]
  assign alu_io_in_bits_src1 = io__in_bits_data_src1; // @[src/main/scala/nutcore/backend/seq/EXU.scala 38:34]
  assign alu_io_in_bits_src2 = io__in_bits_data_src2; // @[src/main/scala/nutcore/backend/seq/EXU.scala 39:34]
  assign alu_io_in_bits_func = io__in_bits_ctrl_fuOpType; // @[src/main/scala/nutcore/backend/fu/ALU.scala 83:15]
  assign alu_io_out_ready = 1'h1; // @[src/main/scala/nutcore/backend/seq/EXU.scala 50:20]
  assign alu_io_cfIn_instr = io__in_bits_cf_instr; // @[src/main/scala/nutcore/backend/seq/EXU.scala 48:15]
  assign alu_io_cfIn_pc = io__in_bits_cf_pc; // @[src/main/scala/nutcore/backend/seq/EXU.scala 48:15]
  assign alu_io_cfIn_pnpc = io__in_bits_cf_pnpc; // @[src/main/scala/nutcore/backend/seq/EXU.scala 48:15]
  assign alu_io_cfIn_brIdx = io__in_bits_cf_brIdx; // @[src/main/scala/nutcore/backend/seq/EXU.scala 48:15]
  assign alu_io_offset = io__in_bits_data_imm; // @[src/main/scala/nutcore/backend/seq/EXU.scala 49:17]
  assign alu_DISPLAY_ENABLE = DISPLAY_ENABLE;
  assign lsu_clock = clock;
  assign lsu_reset = reset;
  assign lsu_io__in_valid = io__in_bits_ctrl_fuType == 3'h1 & io__in_valid & ~io__flush; // @[src/main/scala/nutcore/backend/seq/EXU.scala 44:81]
  assign lsu_io__in_bits_src1 = io__in_bits_data_src1; // @[src/main/scala/nutcore/backend/seq/EXU.scala 38:34]
  assign lsu_io__in_bits_src2 = io__in_bits_data_imm; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 42:15]
  assign lsu_io__in_bits_func = io__in_bits_ctrl_fuOpType; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 43:15]
  assign lsu_io__out_ready = 1'h1; // @[src/main/scala/nutcore/backend/seq/EXU.scala 61:20]
  assign lsu_io__wdata = io__in_bits_data_src2; // @[src/main/scala/nutcore/backend/seq/EXU.scala 39:34]
  assign lsu_io__instr = io__in_bits_cf_instr[31:0]; // @[src/main/scala/nutcore/backend/seq/EXU.scala 58:16]
  assign lsu_io__dmem_req_ready = io__dmem_req_ready; // @[src/main/scala/nutcore/backend/seq/EXU.scala 60:11]
  assign lsu_io__dmem_resp_valid = io__dmem_resp_valid; // @[src/main/scala/nutcore/backend/seq/EXU.scala 60:11]
  assign lsu_io__dmem_resp_bits_rdata = io__dmem_resp_bits_rdata; // @[src/main/scala/nutcore/backend/seq/EXU.scala 60:11]
  assign lsu_lr_0 = csr_lr_0;
  assign lsu_lr_addr = csr_lrAddr_0;
  assign lsu_DISPLAY_ENABLE = DISPLAY_ENABLE;
  assign lsu_DTLBPF = _WIRE_1_1;
  assign lsu_DTLBENABLE = _WIRE_2_3;
  assign lsu_DTLBFINISH = _WIRE_16;
  assign lsu_lsuMMIO_0 = _WIRE_17;
  assign mdu_clock = clock;
  assign mdu_reset = reset;
  assign mdu_io_in_valid = io__in_bits_ctrl_fuType == 3'h2 & io__in_valid & ~io__flush; // @[src/main/scala/nutcore/backend/seq/EXU.scala 44:81]
  assign mdu_io_in_bits_src1 = io__in_bits_data_src1; // @[src/main/scala/nutcore/backend/seq/EXU.scala 38:34]
  assign mdu_io_in_bits_src2 = io__in_bits_data_src2; // @[src/main/scala/nutcore/backend/seq/EXU.scala 39:34]
  assign mdu_io_in_bits_func = io__in_bits_ctrl_fuOpType; // @[src/main/scala/nutcore/backend/fu/MDU.scala 143:15]
  assign mdu_io_out_ready = 1'h1; // @[src/main/scala/nutcore/backend/seq/EXU.scala 65:20]
  assign mdu_DISPLAY_ENABLE = DISPLAY_ENABLE;
  assign csr_clock = clock;
  assign csr_reset = reset;
  assign csr_io_in_valid = io__in_bits_ctrl_fuType == 3'h3 & io__in_valid & ~io__flush; // @[src/main/scala/nutcore/backend/seq/EXU.scala 44:81]
  assign csr_io_in_bits_src1 = io__in_bits_data_src1; // @[src/main/scala/nutcore/backend/seq/EXU.scala 38:34]
  assign csr_io_in_bits_src2 = io__in_bits_data_src2; // @[src/main/scala/nutcore/backend/seq/EXU.scala 39:34]
  assign csr_io_in_bits_func = io__in_bits_ctrl_fuOpType; // @[src/main/scala/nutcore/backend/fu/CSR.scala 200:15]
  assign csr_io_out_ready = 1'h1; // @[src/main/scala/nutcore/backend/seq/EXU.scala 77:20]
  assign csr_io_cfIn_instr = io__in_bits_cf_instr; // @[src/main/scala/nutcore/backend/seq/EXU.scala 70:15]
  assign csr_io_cfIn_pc = io__in_bits_cf_pc; // @[src/main/scala/nutcore/backend/seq/EXU.scala 70:15]
  assign csr_io_cfIn_exceptionVec_1 = io__in_bits_cf_exceptionVec_1; // @[src/main/scala/nutcore/backend/seq/EXU.scala 70:15]
  assign csr_io_cfIn_exceptionVec_2 = io__in_bits_cf_exceptionVec_2; // @[src/main/scala/nutcore/backend/seq/EXU.scala 70:15]
  assign csr_io_cfIn_exceptionVec_4 = lsu_io__loadAddrMisaligned; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:48]
  assign csr_io_cfIn_exceptionVec_6 = lsu_io__storeAddrMisaligned; // @[src/main/scala/nutcore/backend/seq/EXU.scala 72:49]
  assign csr_io_cfIn_exceptionVec_12 = io__in_bits_cf_exceptionVec_12; // @[src/main/scala/nutcore/backend/seq/EXU.scala 70:15]
  assign csr_io_cfIn_intrVec_0 = io__in_bits_cf_intrVec_0; // @[src/main/scala/nutcore/backend/seq/EXU.scala 70:15]
  assign csr_io_cfIn_intrVec_1 = io__in_bits_cf_intrVec_1; // @[src/main/scala/nutcore/backend/seq/EXU.scala 70:15]
  assign csr_io_cfIn_intrVec_2 = io__in_bits_cf_intrVec_2; // @[src/main/scala/nutcore/backend/seq/EXU.scala 70:15]
  assign csr_io_cfIn_intrVec_3 = io__in_bits_cf_intrVec_3; // @[src/main/scala/nutcore/backend/seq/EXU.scala 70:15]
  assign csr_io_cfIn_intrVec_4 = io__in_bits_cf_intrVec_4; // @[src/main/scala/nutcore/backend/seq/EXU.scala 70:15]
  assign csr_io_cfIn_intrVec_5 = io__in_bits_cf_intrVec_5; // @[src/main/scala/nutcore/backend/seq/EXU.scala 70:15]
  assign csr_io_cfIn_intrVec_6 = io__in_bits_cf_intrVec_6; // @[src/main/scala/nutcore/backend/seq/EXU.scala 70:15]
  assign csr_io_cfIn_intrVec_7 = io__in_bits_cf_intrVec_7; // @[src/main/scala/nutcore/backend/seq/EXU.scala 70:15]
  assign csr_io_cfIn_intrVec_8 = io__in_bits_cf_intrVec_8; // @[src/main/scala/nutcore/backend/seq/EXU.scala 70:15]
  assign csr_io_cfIn_intrVec_9 = io__in_bits_cf_intrVec_9; // @[src/main/scala/nutcore/backend/seq/EXU.scala 70:15]
  assign csr_io_cfIn_intrVec_10 = io__in_bits_cf_intrVec_10; // @[src/main/scala/nutcore/backend/seq/EXU.scala 70:15]
  assign csr_io_cfIn_intrVec_11 = io__in_bits_cf_intrVec_11; // @[src/main/scala/nutcore/backend/seq/EXU.scala 70:15]
  assign csr_io_cfIn_crossPageIPFFix = io__in_bits_cf_crossPageIPFFix; // @[src/main/scala/nutcore/backend/seq/EXU.scala 70:15]
  assign csr_io_instrValid = io__in_valid & _fuValids_0_T_2; // @[src/main/scala/nutcore/backend/seq/EXU.scala 73:36]
  assign csr_io_dmemMMU_loadPF = io__memMMU_dmem_loadPF; // @[src/main/scala/nutcore/backend/seq/EXU.scala 80:18]
  assign csr_io_dmemMMU_storePF = io__memMMU_dmem_storePF; // @[src/main/scala/nutcore/backend/seq/EXU.scala 80:18]
  assign csr_io_dmemMMU_addr = io__memMMU_dmem_addr; // @[src/main/scala/nutcore/backend/seq/EXU.scala 80:18]
  assign csr_set_lr = lsu_setLr_0;
  assign csr_MbpBWrong = alu__WIRE_2_0;
  assign csr_perfCntCondMmulInstr = mdu__WIRE_0;
  assign csr_meip_0 = io_extra_meip_0;
  assign csr_perfCntCondMlsuInstr = _WIRE_2;
  assign csr_perfCntCondMexuBusy = _WIRE_1_0;
  assign csr_perfCntCondMmmioInstr = lsu_io_isMMIO;
  assign csr_perfCntCondMaluInstr = _WIRE;
  assign csr_MbpRRight = alu__WIRE_15_0;
  assign csr_DISPLAY_ENABLE = DISPLAY_ENABLE;
  assign csr_MbpIRight = alu__WIRE_13_0;
  assign csr_perfCntCondMcsrInstr = _WIRE_4;
  assign csr_Custom4 = alu__WIRE_6_0;
  assign csr_Custom3 = alu__WIRE_5_0;
  assign csr_perfCntCondMifuFlush = _WIRE_8;
  assign csr_Custom2 = alu__WIRE_4_1;
  assign csr_Custom1 = alu__WIRE_3_0;
  assign csr_Custom8 = alu__WIRE_10_0;
  assign csr_Custom7 = alu__WIRE_9_0;
  assign csr_perfCntCondMrawStall = _WIRE_11;
  assign csr_perfCntCondMloadStall = lsu_r;
  assign csr_Custom6 = alu__WIRE_8_0;
  assign csr_Custom5 = alu__WIRE_7_0;
  assign csr_perfCntCondISUIssue = _WIRE_2_2;
  assign csr_mtip_0 = io_extra_mtip;
  assign csr_perfCntCondMultiCommit = falseWire;
  assign csr_MbpBRight = alu__WIRE_1_2;
  assign csr_perfCntCondMbruInstr = _WIRE_1;
  assign csr_set_lr_val = lsu_setLrVal_0;
  assign csr_MbpJWrong = alu__WIRE_12_0;
  assign csr_nutcoretrap_0 = nutcoretrap;
  assign csr_LSUADDR = lsu_io_in_bits_src1;
  assign csr_perfCntCondMstoreStall = lsu_r_1;
  assign csr_MbpIWrong = alu__WIRE_14_0;
  assign csr_MbpJRight = alu__WIRE_11_0;
  assign csr_perfCntCondMloadInstr = lsu__WIRE_16;
  assign csr_perfCntCondMmduInstr = _WIRE_3;
  assign csr_set_lr_addr = lsu_setLrAddr_0;
  assign csr_perfCntCondMimemStall = r_0;
  assign csr_MbpRWrong = alu__WIRE_16_0;
  assign csr_msip_0 = io_extra_msip;
  assign csr_perfCntCondMinstret = io_in_valid;
  assign mou_clock = clock;
  assign mou_reset = reset;
  assign mou_io_in_valid = io__in_bits_ctrl_fuType == 3'h4 & io__in_valid & ~io__flush; // @[src/main/scala/nutcore/backend/seq/EXU.scala 44:81]
  assign mou_io_in_bits_func = io__in_bits_ctrl_fuOpType; // @[src/main/scala/nutcore/backend/fu/MOU.scala 45:15]
  assign mou_io_cfIn_pc = io__in_bits_cf_pc; // @[src/main/scala/nutcore/backend/seq/EXU.scala 85:15]
  assign mou_DISPLAY_ENABLE = DISPLAY_ENABLE;
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/utils/GTimer.scala 24:20]
      c <= 64'h0; // @[src/main/scala/utils/GTimer.scala 24:20]
    end else begin
      c <= _c_T_1; // @[src/main/scala/utils/GTimer.scala 25:7]
    end
    if (reset) begin // @[src/main/scala/utils/GTimer.scala 24:20]
      c_1 <= 64'h0; // @[src/main/scala/utils/GTimer.scala 24:20]
    end else begin
      c_1 <= _c_T_3; // @[src/main/scala/utils/GTimer.scala 25:7]
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2 & ~reset) begin
          $fwrite(32'h80000002,"[%d] EXU: ",c); // @[src/main/scala/utils/Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2 & _T_4) begin
          $fwrite(32'h80000002,"[REDIRECT] mou %x csr %x alu %x \n",mou_io_redirect_valid,csr_io_redirect_valid,
            alu_io_redirect_valid); // @[src/main/scala/utils/Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2 & ~reset) begin
          $fwrite(32'h80000002,"[%d] EXU: ",c_1); // @[src/main/scala/utils/Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2 & _T_4) begin
          $fwrite(32'h80000002,"[REDIRECT] flush: %d mou %x csr %x alu %x\n",io__flush,mou_io_redirect_target,
            csr_io_redirect_target,alu_io_redirect_target); // @[src/main/scala/utils/Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  c = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  c_1 = _RAND_1[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module WBU(
  input         clock,
  input         reset,
  input         io__in_valid, // @[src/main/scala/nutcore/backend/seq/WBU.scala 26:14]
  input  [63:0] io__in_bits_decode_cf_instr, // @[src/main/scala/nutcore/backend/seq/WBU.scala 26:14]
  input  [38:0] io__in_bits_decode_cf_pc, // @[src/main/scala/nutcore/backend/seq/WBU.scala 26:14]
  input  [38:0] io__in_bits_decode_cf_redirect_target, // @[src/main/scala/nutcore/backend/seq/WBU.scala 26:14]
  input         io__in_bits_decode_cf_redirect_valid, // @[src/main/scala/nutcore/backend/seq/WBU.scala 26:14]
  input  [2:0]  io__in_bits_decode_ctrl_fuType, // @[src/main/scala/nutcore/backend/seq/WBU.scala 26:14]
  input         io__in_bits_decode_ctrl_rfWen, // @[src/main/scala/nutcore/backend/seq/WBU.scala 26:14]
  input  [4:0]  io__in_bits_decode_ctrl_rfDest, // @[src/main/scala/nutcore/backend/seq/WBU.scala 26:14]
  input         io__in_bits_isMMIO, // @[src/main/scala/nutcore/backend/seq/WBU.scala 26:14]
  input  [63:0] io__in_bits_intrNO, // @[src/main/scala/nutcore/backend/seq/WBU.scala 26:14]
  input  [63:0] io__in_bits_commits_0, // @[src/main/scala/nutcore/backend/seq/WBU.scala 26:14]
  input  [63:0] io__in_bits_commits_1, // @[src/main/scala/nutcore/backend/seq/WBU.scala 26:14]
  input  [63:0] io__in_bits_commits_2, // @[src/main/scala/nutcore/backend/seq/WBU.scala 26:14]
  input  [63:0] io__in_bits_commits_3, // @[src/main/scala/nutcore/backend/seq/WBU.scala 26:14]
  output        io__wb_rfWen, // @[src/main/scala/nutcore/backend/seq/WBU.scala 26:14]
  output [4:0]  io__wb_rfDest, // @[src/main/scala/nutcore/backend/seq/WBU.scala 26:14]
  output [63:0] io__wb_rfData, // @[src/main/scala/nutcore/backend/seq/WBU.scala 26:14]
  output [38:0] io__redirect_target, // @[src/main/scala/nutcore/backend/seq/WBU.scala 26:14]
  output        io__redirect_valid, // @[src/main/scala/nutcore/backend/seq/WBU.scala 26:14]
  input         DISPLAY_ENABLE,
  output        falseWire_0,
  output        io_in_valid
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire [63:0] _GEN_1 = 3'h1 == io__in_bits_decode_ctrl_fuType ? io__in_bits_commits_1 : io__in_bits_commits_0; // @[src/main/scala/nutcore/backend/seq/WBU.scala 34:{16,16}]
  wire [63:0] _GEN_2 = 3'h2 == io__in_bits_decode_ctrl_fuType ? io__in_bits_commits_2 : _GEN_1; // @[src/main/scala/nutcore/backend/seq/WBU.scala 34:{16,16}]
  wire [63:0] _GEN_3 = 3'h3 == io__in_bits_decode_ctrl_fuType ? io__in_bits_commits_3 : _GEN_2; // @[src/main/scala/nutcore/backend/seq/WBU.scala 34:{16,16}]
  reg [63:0] c; // @[src/main/scala/utils/GTimer.scala 24:20]
  wire [63:0] _c_T_1 = c + 64'h1; // @[src/main/scala/utils/GTimer.scala 25:12]
  wire  _T = io__in_valid & DISPLAY_ENABLE; // @[src/main/scala/utils/Debug.scala 55:16]
  wire  _T_2 = ~reset; // @[src/main/scala/utils/Debug.scala 56:24]
  wire  falseWire = 1'h0; // @[src/main/scala/nutcore/backend/seq/WBU.scala 43:{27,27}]
  assign io__wb_rfWen = io__in_bits_decode_ctrl_rfWen & io__in_valid; // @[src/main/scala/nutcore/backend/seq/WBU.scala 32:47]
  assign io__wb_rfDest = io__in_bits_decode_ctrl_rfDest; // @[src/main/scala/nutcore/backend/seq/WBU.scala 33:16]
  assign io__wb_rfData = 3'h4 == io__in_bits_decode_ctrl_fuType ? 64'h0 : _GEN_3; // @[src/main/scala/nutcore/backend/seq/WBU.scala 34:{16,16}]
  assign io__redirect_target = io__in_bits_decode_cf_redirect_target; // @[src/main/scala/nutcore/backend/seq/WBU.scala 38:15]
  assign io__redirect_valid = io__in_bits_decode_cf_redirect_valid & io__in_valid; // @[src/main/scala/nutcore/backend/seq/WBU.scala 39:60]
  assign falseWire_0 = falseWire;
  assign io_in_valid = io__in_valid;
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/utils/GTimer.scala 24:20]
      c <= 64'h0; // @[src/main/scala/utils/GTimer.scala 24:20]
    end else begin
      c <= _c_T_1; // @[src/main/scala/utils/GTimer.scala 25:7]
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T & ~reset) begin
          $fwrite(32'h80000002,"[%d] WBU: ",c); // @[src/main/scala/utils/Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T & _T_2) begin
          $fwrite(32'h80000002,"[COMMIT] pc = 0x%x inst %x wen %x wdst %x wdata %x mmio %x intrNO %x\n",
            io__in_bits_decode_cf_pc,io__in_bits_decode_cf_instr,io__wb_rfWen,io__wb_rfDest,io__wb_rfData,
            io__in_bits_isMMIO,io__in_bits_intrNO); // @[src/main/scala/utils/Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  c = _RAND_0[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Backend_inorder(
  input         clock,
  input         reset,
  output        io_in_0_ready, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  input         io_in_0_valid, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  input  [63:0] io_in_0_bits_cf_instr, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  input  [38:0] io_in_0_bits_cf_pc, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  input  [38:0] io_in_0_bits_cf_pnpc, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  input         io_in_0_bits_cf_exceptionVec_1, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  input         io_in_0_bits_cf_exceptionVec_2, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  input         io_in_0_bits_cf_exceptionVec_12, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  input         io_in_0_bits_cf_intrVec_0, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  input         io_in_0_bits_cf_intrVec_1, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  input         io_in_0_bits_cf_intrVec_2, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  input         io_in_0_bits_cf_intrVec_3, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  input         io_in_0_bits_cf_intrVec_4, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  input         io_in_0_bits_cf_intrVec_5, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  input         io_in_0_bits_cf_intrVec_6, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  input         io_in_0_bits_cf_intrVec_7, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  input         io_in_0_bits_cf_intrVec_8, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  input         io_in_0_bits_cf_intrVec_9, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  input         io_in_0_bits_cf_intrVec_10, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  input         io_in_0_bits_cf_intrVec_11, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  input  [3:0]  io_in_0_bits_cf_brIdx, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  input         io_in_0_bits_cf_crossPageIPFFix, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  input         io_in_0_bits_ctrl_src1Type, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  input         io_in_0_bits_ctrl_src2Type, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  input  [2:0]  io_in_0_bits_ctrl_fuType, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  input  [6:0]  io_in_0_bits_ctrl_fuOpType, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  input  [4:0]  io_in_0_bits_ctrl_rfSrc1, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  input  [4:0]  io_in_0_bits_ctrl_rfSrc2, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  input         io_in_0_bits_ctrl_rfWen, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  input  [4:0]  io_in_0_bits_ctrl_rfDest, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  input         io_in_0_bits_ctrl_isNutCoreTrap, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  input  [63:0] io_in_0_bits_data_imm, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  input  [1:0]  io_flush, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  input         io_dmem_req_ready, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  output        io_dmem_req_valid, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  output [38:0] io_dmem_req_bits_addr, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  output [2:0]  io_dmem_req_bits_size, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  output [3:0]  io_dmem_req_bits_cmd, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  output [7:0]  io_dmem_req_bits_wmask, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  output [63:0] io_dmem_req_bits_wdata, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  input         io_dmem_resp_valid, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  input  [63:0] io_dmem_resp_bits_rdata, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  output [1:0]  io_memMMU_imem_priviledgeMode, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  output [1:0]  io_memMMU_dmem_priviledgeMode, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  output        io_memMMU_dmem_status_sum, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  output        io_memMMU_dmem_status_mxr, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  input         io_memMMU_dmem_loadPF, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  input         io_memMMU_dmem_storePF, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  input  [38:0] io_memMMU_dmem_addr, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  output [38:0] io_redirect_target, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  output        io_redirect_valid, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  input         io_extra_meip_0,
  output        REG_valid,
  output [38:0] REG_pc,
  output        REG_isMissPredict,
  output [38:0] REG_actualTarget,
  output        REG_actualTaken,
  output [6:0]  REG_fuOpType,
  output [1:0]  REG_btbType,
  output        REG_isRVC,
  output        _WIRE_1,
  output [63:0] satp,
  input         _WIRE_4,
  input         _WIRE_1_1,
  input         _WIRE_7,
  input         io_extra_mtip,
  output        _WIRE_11,
  output        _WIRE_1_4,
  output [11:0] _WIRE_14,
  input         _WIRE_2_2,
  input         _WIRE_16,
  input         _WIRE_17,
  input         r_0,
  input         io_extra_msip
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [63:0] _RAND_26;
  reg [63:0] _RAND_27;
  reg [63:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [63:0] _RAND_30;
  reg [63:0] _RAND_31;
  reg [63:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [63:0] _RAND_38;
  reg [63:0] _RAND_39;
  reg [63:0] _RAND_40;
  reg [63:0] _RAND_41;
  reg [63:0] _RAND_42;
`endif // RANDOMIZE_REG_INIT
  wire  isu_clock; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 678:20]
  wire  isu_reset; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 678:20]
  wire  isu_io_in_0_ready; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 678:20]
  wire  isu_io_in_0_valid; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 678:20]
  wire [63:0] isu_io_in_0_bits_cf_instr; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 678:20]
  wire [38:0] isu_io_in_0_bits_cf_pc; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 678:20]
  wire [38:0] isu_io_in_0_bits_cf_pnpc; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 678:20]
  wire  isu_io_in_0_bits_cf_exceptionVec_1; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 678:20]
  wire  isu_io_in_0_bits_cf_exceptionVec_2; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 678:20]
  wire  isu_io_in_0_bits_cf_exceptionVec_12; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 678:20]
  wire  isu_io_in_0_bits_cf_intrVec_0; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 678:20]
  wire  isu_io_in_0_bits_cf_intrVec_1; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 678:20]
  wire  isu_io_in_0_bits_cf_intrVec_2; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 678:20]
  wire  isu_io_in_0_bits_cf_intrVec_3; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 678:20]
  wire  isu_io_in_0_bits_cf_intrVec_4; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 678:20]
  wire  isu_io_in_0_bits_cf_intrVec_5; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 678:20]
  wire  isu_io_in_0_bits_cf_intrVec_6; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 678:20]
  wire  isu_io_in_0_bits_cf_intrVec_7; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 678:20]
  wire  isu_io_in_0_bits_cf_intrVec_8; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 678:20]
  wire  isu_io_in_0_bits_cf_intrVec_9; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 678:20]
  wire  isu_io_in_0_bits_cf_intrVec_10; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 678:20]
  wire  isu_io_in_0_bits_cf_intrVec_11; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 678:20]
  wire [3:0] isu_io_in_0_bits_cf_brIdx; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 678:20]
  wire  isu_io_in_0_bits_cf_crossPageIPFFix; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 678:20]
  wire  isu_io_in_0_bits_ctrl_src1Type; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 678:20]
  wire  isu_io_in_0_bits_ctrl_src2Type; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 678:20]
  wire [2:0] isu_io_in_0_bits_ctrl_fuType; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 678:20]
  wire [6:0] isu_io_in_0_bits_ctrl_fuOpType; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 678:20]
  wire [4:0] isu_io_in_0_bits_ctrl_rfSrc1; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 678:20]
  wire [4:0] isu_io_in_0_bits_ctrl_rfSrc2; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 678:20]
  wire  isu_io_in_0_bits_ctrl_rfWen; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 678:20]
  wire [4:0] isu_io_in_0_bits_ctrl_rfDest; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 678:20]
  wire  isu_io_in_0_bits_ctrl_isNutCoreTrap; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 678:20]
  wire [63:0] isu_io_in_0_bits_data_imm; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 678:20]
  wire  isu_io_out_ready; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 678:20]
  wire  isu_io_out_valid; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 678:20]
  wire [63:0] isu_io_out_bits_cf_instr; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 678:20]
  wire [38:0] isu_io_out_bits_cf_pc; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 678:20]
  wire [38:0] isu_io_out_bits_cf_pnpc; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 678:20]
  wire  isu_io_out_bits_cf_exceptionVec_1; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 678:20]
  wire  isu_io_out_bits_cf_exceptionVec_2; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 678:20]
  wire  isu_io_out_bits_cf_exceptionVec_12; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 678:20]
  wire  isu_io_out_bits_cf_intrVec_0; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 678:20]
  wire  isu_io_out_bits_cf_intrVec_1; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 678:20]
  wire  isu_io_out_bits_cf_intrVec_2; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 678:20]
  wire  isu_io_out_bits_cf_intrVec_3; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 678:20]
  wire  isu_io_out_bits_cf_intrVec_4; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 678:20]
  wire  isu_io_out_bits_cf_intrVec_5; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 678:20]
  wire  isu_io_out_bits_cf_intrVec_6; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 678:20]
  wire  isu_io_out_bits_cf_intrVec_7; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 678:20]
  wire  isu_io_out_bits_cf_intrVec_8; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 678:20]
  wire  isu_io_out_bits_cf_intrVec_9; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 678:20]
  wire  isu_io_out_bits_cf_intrVec_10; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 678:20]
  wire  isu_io_out_bits_cf_intrVec_11; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 678:20]
  wire [3:0] isu_io_out_bits_cf_brIdx; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 678:20]
  wire  isu_io_out_bits_cf_crossPageIPFFix; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 678:20]
  wire [2:0] isu_io_out_bits_ctrl_fuType; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 678:20]
  wire [6:0] isu_io_out_bits_ctrl_fuOpType; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 678:20]
  wire  isu_io_out_bits_ctrl_rfWen; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 678:20]
  wire [4:0] isu_io_out_bits_ctrl_rfDest; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 678:20]
  wire  isu_io_out_bits_ctrl_isNutCoreTrap; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 678:20]
  wire [63:0] isu_io_out_bits_data_src1; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 678:20]
  wire [63:0] isu_io_out_bits_data_src2; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 678:20]
  wire [63:0] isu_io_out_bits_data_imm; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 678:20]
  wire  isu_io_wb_rfWen; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 678:20]
  wire [4:0] isu_io_wb_rfDest; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 678:20]
  wire [63:0] isu_io_wb_rfData; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 678:20]
  wire  isu_io_forward_valid; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 678:20]
  wire  isu_io_forward_wb_rfWen; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 678:20]
  wire [4:0] isu_io_forward_wb_rfDest; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 678:20]
  wire [63:0] isu_io_forward_wb_rfData; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 678:20]
  wire [2:0] isu_io_forward_fuType; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 678:20]
  wire  isu_io_flush; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 678:20]
  wire  isu__WIRE_1_0; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 678:20]
  wire  isu_DISPLAY_ENABLE; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 678:20]
  wire  isu__WIRE_8; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 678:20]
  wire  isu__WIRE_2_2; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 678:20]
  wire  exu_clock; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire  exu_reset; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire  exu_io__in_ready; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire  exu_io__in_valid; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire [63:0] exu_io__in_bits_cf_instr; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire [38:0] exu_io__in_bits_cf_pc; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire [38:0] exu_io__in_bits_cf_pnpc; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire  exu_io__in_bits_cf_exceptionVec_1; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire  exu_io__in_bits_cf_exceptionVec_2; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire  exu_io__in_bits_cf_exceptionVec_12; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire  exu_io__in_bits_cf_intrVec_0; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire  exu_io__in_bits_cf_intrVec_1; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire  exu_io__in_bits_cf_intrVec_2; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire  exu_io__in_bits_cf_intrVec_3; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire  exu_io__in_bits_cf_intrVec_4; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire  exu_io__in_bits_cf_intrVec_5; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire  exu_io__in_bits_cf_intrVec_6; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire  exu_io__in_bits_cf_intrVec_7; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire  exu_io__in_bits_cf_intrVec_8; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire  exu_io__in_bits_cf_intrVec_9; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire  exu_io__in_bits_cf_intrVec_10; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire  exu_io__in_bits_cf_intrVec_11; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire [3:0] exu_io__in_bits_cf_brIdx; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire  exu_io__in_bits_cf_crossPageIPFFix; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire [2:0] exu_io__in_bits_ctrl_fuType; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire [6:0] exu_io__in_bits_ctrl_fuOpType; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire  exu_io__in_bits_ctrl_rfWen; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire [4:0] exu_io__in_bits_ctrl_rfDest; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire  exu_io__in_bits_ctrl_isNutCoreTrap; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire [63:0] exu_io__in_bits_data_src1; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire [63:0] exu_io__in_bits_data_src2; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire [63:0] exu_io__in_bits_data_imm; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire  exu_io__out_ready; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire  exu_io__out_valid; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire [63:0] exu_io__out_bits_decode_cf_instr; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire [38:0] exu_io__out_bits_decode_cf_pc; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire [38:0] exu_io__out_bits_decode_cf_redirect_target; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire  exu_io__out_bits_decode_cf_redirect_valid; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire [2:0] exu_io__out_bits_decode_ctrl_fuType; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire  exu_io__out_bits_decode_ctrl_rfWen; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire [4:0] exu_io__out_bits_decode_ctrl_rfDest; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire  exu_io__out_bits_isMMIO; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire [63:0] exu_io__out_bits_intrNO; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire [63:0] exu_io__out_bits_commits_0; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire [63:0] exu_io__out_bits_commits_1; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire [63:0] exu_io__out_bits_commits_2; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire [63:0] exu_io__out_bits_commits_3; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire  exu_io__flush; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire  exu_io__dmem_req_ready; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire  exu_io__dmem_req_valid; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire [38:0] exu_io__dmem_req_bits_addr; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire [2:0] exu_io__dmem_req_bits_size; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire [3:0] exu_io__dmem_req_bits_cmd; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire [7:0] exu_io__dmem_req_bits_wmask; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire [63:0] exu_io__dmem_req_bits_wdata; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire  exu_io__dmem_resp_valid; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire [63:0] exu_io__dmem_resp_bits_rdata; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire  exu_io__forward_valid; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire  exu_io__forward_wb_rfWen; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire [4:0] exu_io__forward_wb_rfDest; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire [63:0] exu_io__forward_wb_rfData; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire [2:0] exu_io__forward_fuType; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire [1:0] exu_io__memMMU_imem_priviledgeMode; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire [1:0] exu_io__memMMU_dmem_priviledgeMode; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire  exu_io__memMMU_dmem_status_sum; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire  exu_io__memMMU_dmem_status_mxr; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire  exu_io__memMMU_dmem_loadPF; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire  exu_io__memMMU_dmem_storePF; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire [38:0] exu_io__memMMU_dmem_addr; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire  exu_io_extra_meip_0; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire  exu_REG_valid; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire [38:0] exu_REG_pc; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire  exu_REG_isMissPredict; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire [38:0] exu_REG_actualTarget; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire  exu_REG_actualTaken; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire [6:0] exu_REG_fuOpType; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire [1:0] exu_REG_btbType; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire  exu_REG_isRVC; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire  exu__WIRE_6; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire  exu__WIRE_1_0; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire [63:0] exu_satp; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire  exu_DISPLAY_ENABLE; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire  exu__WIRE_1_1; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire  exu__WIRE_8; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire  exu__WIRE_11; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire  exu__WIRE_2_2; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire  exu_io_extra_mtip; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire  exu__WIRE_12; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire  exu_falseWire; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire  exu__WIRE_1_4; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire [11:0] exu__WIRE_14; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire  exu__WIRE_2_3; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire  exu__WIRE_16; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire  exu__WIRE_17; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire  exu_r_0; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire  exu_io_extra_msip; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire  exu_io_in_valid; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire  wbu_clock; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  wbu_reset; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  wbu_io__in_valid; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire [63:0] wbu_io__in_bits_decode_cf_instr; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire [38:0] wbu_io__in_bits_decode_cf_pc; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire [38:0] wbu_io__in_bits_decode_cf_redirect_target; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  wbu_io__in_bits_decode_cf_redirect_valid; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire [2:0] wbu_io__in_bits_decode_ctrl_fuType; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  wbu_io__in_bits_decode_ctrl_rfWen; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire [4:0] wbu_io__in_bits_decode_ctrl_rfDest; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  wbu_io__in_bits_isMMIO; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire [63:0] wbu_io__in_bits_intrNO; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire [63:0] wbu_io__in_bits_commits_0; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire [63:0] wbu_io__in_bits_commits_1; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire [63:0] wbu_io__in_bits_commits_2; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire [63:0] wbu_io__in_bits_commits_3; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  wbu_io__wb_rfWen; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire [4:0] wbu_io__wb_rfDest; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire [63:0] wbu_io__wb_rfData; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire [38:0] wbu_io__redirect_target; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  wbu_io__redirect_valid; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  wbu_DISPLAY_ENABLE; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  wbu_falseWire_0; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  wbu_io_in_valid; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  _T = exu_io__out_ready & exu_io__out_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  reg  valid; // @[src/main/scala/utils/Pipeline.scala 24:24]
  wire  _GEN_0 = _T ? 1'h0 : valid; // @[src/main/scala/utils/Pipeline.scala 24:24 25:{25,33}]
  wire  _T_2 = isu_io_out_valid & exu_io__in_ready; // @[src/main/scala/utils/Pipeline.scala 26:22]
  wire  _GEN_1 = isu_io_out_valid & exu_io__in_ready | _GEN_0; // @[src/main/scala/utils/Pipeline.scala 26:{38,46}]
  reg [63:0] exu_io_in_bits_r_cf_instr; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg [38:0] exu_io_in_bits_r_cf_pc; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg [38:0] exu_io_in_bits_r_cf_pnpc; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg  exu_io_in_bits_r_cf_exceptionVec_1; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg  exu_io_in_bits_r_cf_exceptionVec_2; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg  exu_io_in_bits_r_cf_exceptionVec_12; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg  exu_io_in_bits_r_cf_intrVec_0; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg  exu_io_in_bits_r_cf_intrVec_1; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg  exu_io_in_bits_r_cf_intrVec_2; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg  exu_io_in_bits_r_cf_intrVec_3; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg  exu_io_in_bits_r_cf_intrVec_4; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg  exu_io_in_bits_r_cf_intrVec_5; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg  exu_io_in_bits_r_cf_intrVec_6; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg  exu_io_in_bits_r_cf_intrVec_7; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg  exu_io_in_bits_r_cf_intrVec_8; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg  exu_io_in_bits_r_cf_intrVec_9; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg  exu_io_in_bits_r_cf_intrVec_10; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg  exu_io_in_bits_r_cf_intrVec_11; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg [3:0] exu_io_in_bits_r_cf_brIdx; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg  exu_io_in_bits_r_cf_crossPageIPFFix; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg [2:0] exu_io_in_bits_r_ctrl_fuType; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg [6:0] exu_io_in_bits_r_ctrl_fuOpType; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg  exu_io_in_bits_r_ctrl_rfWen; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg [4:0] exu_io_in_bits_r_ctrl_rfDest; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg  exu_io_in_bits_r_ctrl_isNutCoreTrap; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg [63:0] exu_io_in_bits_r_data_src1; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg [63:0] exu_io_in_bits_r_data_src2; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg [63:0] exu_io_in_bits_r_data_imm; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg  valid_1; // @[src/main/scala/utils/Pipeline.scala 24:24]
  wire  _T_4 = exu_io__out_valid; // @[src/main/scala/utils/Pipeline.scala 26:22]
  reg [63:0] wbu_io_in_bits_r_decode_cf_instr; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg [38:0] wbu_io_in_bits_r_decode_cf_pc; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg [38:0] wbu_io_in_bits_r_decode_cf_redirect_target; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg  wbu_io_in_bits_r_decode_cf_redirect_valid; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg [2:0] wbu_io_in_bits_r_decode_ctrl_fuType; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg  wbu_io_in_bits_r_decode_ctrl_rfWen; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg [4:0] wbu_io_in_bits_r_decode_ctrl_rfDest; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg  wbu_io_in_bits_r_isMMIO; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg [63:0] wbu_io_in_bits_r_intrNO; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg [63:0] wbu_io_in_bits_r_commits_0; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg [63:0] wbu_io_in_bits_r_commits_1; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg [63:0] wbu_io_in_bits_r_commits_2; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg [63:0] wbu_io_in_bits_r_commits_3; // @[src/main/scala/utils/Pipeline.scala 30:28]
  ISU isu ( // @[src/main/scala/nutcore/backend/ooo/Backend.scala 678:20]
    .clock(isu_clock),
    .reset(isu_reset),
    .io_in_0_ready(isu_io_in_0_ready),
    .io_in_0_valid(isu_io_in_0_valid),
    .io_in_0_bits_cf_instr(isu_io_in_0_bits_cf_instr),
    .io_in_0_bits_cf_pc(isu_io_in_0_bits_cf_pc),
    .io_in_0_bits_cf_pnpc(isu_io_in_0_bits_cf_pnpc),
    .io_in_0_bits_cf_exceptionVec_1(isu_io_in_0_bits_cf_exceptionVec_1),
    .io_in_0_bits_cf_exceptionVec_2(isu_io_in_0_bits_cf_exceptionVec_2),
    .io_in_0_bits_cf_exceptionVec_12(isu_io_in_0_bits_cf_exceptionVec_12),
    .io_in_0_bits_cf_intrVec_0(isu_io_in_0_bits_cf_intrVec_0),
    .io_in_0_bits_cf_intrVec_1(isu_io_in_0_bits_cf_intrVec_1),
    .io_in_0_bits_cf_intrVec_2(isu_io_in_0_bits_cf_intrVec_2),
    .io_in_0_bits_cf_intrVec_3(isu_io_in_0_bits_cf_intrVec_3),
    .io_in_0_bits_cf_intrVec_4(isu_io_in_0_bits_cf_intrVec_4),
    .io_in_0_bits_cf_intrVec_5(isu_io_in_0_bits_cf_intrVec_5),
    .io_in_0_bits_cf_intrVec_6(isu_io_in_0_bits_cf_intrVec_6),
    .io_in_0_bits_cf_intrVec_7(isu_io_in_0_bits_cf_intrVec_7),
    .io_in_0_bits_cf_intrVec_8(isu_io_in_0_bits_cf_intrVec_8),
    .io_in_0_bits_cf_intrVec_9(isu_io_in_0_bits_cf_intrVec_9),
    .io_in_0_bits_cf_intrVec_10(isu_io_in_0_bits_cf_intrVec_10),
    .io_in_0_bits_cf_intrVec_11(isu_io_in_0_bits_cf_intrVec_11),
    .io_in_0_bits_cf_brIdx(isu_io_in_0_bits_cf_brIdx),
    .io_in_0_bits_cf_crossPageIPFFix(isu_io_in_0_bits_cf_crossPageIPFFix),
    .io_in_0_bits_ctrl_src1Type(isu_io_in_0_bits_ctrl_src1Type),
    .io_in_0_bits_ctrl_src2Type(isu_io_in_0_bits_ctrl_src2Type),
    .io_in_0_bits_ctrl_fuType(isu_io_in_0_bits_ctrl_fuType),
    .io_in_0_bits_ctrl_fuOpType(isu_io_in_0_bits_ctrl_fuOpType),
    .io_in_0_bits_ctrl_rfSrc1(isu_io_in_0_bits_ctrl_rfSrc1),
    .io_in_0_bits_ctrl_rfSrc2(isu_io_in_0_bits_ctrl_rfSrc2),
    .io_in_0_bits_ctrl_rfWen(isu_io_in_0_bits_ctrl_rfWen),
    .io_in_0_bits_ctrl_rfDest(isu_io_in_0_bits_ctrl_rfDest),
    .io_in_0_bits_ctrl_isNutCoreTrap(isu_io_in_0_bits_ctrl_isNutCoreTrap),
    .io_in_0_bits_data_imm(isu_io_in_0_bits_data_imm),
    .io_out_ready(isu_io_out_ready),
    .io_out_valid(isu_io_out_valid),
    .io_out_bits_cf_instr(isu_io_out_bits_cf_instr),
    .io_out_bits_cf_pc(isu_io_out_bits_cf_pc),
    .io_out_bits_cf_pnpc(isu_io_out_bits_cf_pnpc),
    .io_out_bits_cf_exceptionVec_1(isu_io_out_bits_cf_exceptionVec_1),
    .io_out_bits_cf_exceptionVec_2(isu_io_out_bits_cf_exceptionVec_2),
    .io_out_bits_cf_exceptionVec_12(isu_io_out_bits_cf_exceptionVec_12),
    .io_out_bits_cf_intrVec_0(isu_io_out_bits_cf_intrVec_0),
    .io_out_bits_cf_intrVec_1(isu_io_out_bits_cf_intrVec_1),
    .io_out_bits_cf_intrVec_2(isu_io_out_bits_cf_intrVec_2),
    .io_out_bits_cf_intrVec_3(isu_io_out_bits_cf_intrVec_3),
    .io_out_bits_cf_intrVec_4(isu_io_out_bits_cf_intrVec_4),
    .io_out_bits_cf_intrVec_5(isu_io_out_bits_cf_intrVec_5),
    .io_out_bits_cf_intrVec_6(isu_io_out_bits_cf_intrVec_6),
    .io_out_bits_cf_intrVec_7(isu_io_out_bits_cf_intrVec_7),
    .io_out_bits_cf_intrVec_8(isu_io_out_bits_cf_intrVec_8),
    .io_out_bits_cf_intrVec_9(isu_io_out_bits_cf_intrVec_9),
    .io_out_bits_cf_intrVec_10(isu_io_out_bits_cf_intrVec_10),
    .io_out_bits_cf_intrVec_11(isu_io_out_bits_cf_intrVec_11),
    .io_out_bits_cf_brIdx(isu_io_out_bits_cf_brIdx),
    .io_out_bits_cf_crossPageIPFFix(isu_io_out_bits_cf_crossPageIPFFix),
    .io_out_bits_ctrl_fuType(isu_io_out_bits_ctrl_fuType),
    .io_out_bits_ctrl_fuOpType(isu_io_out_bits_ctrl_fuOpType),
    .io_out_bits_ctrl_rfWen(isu_io_out_bits_ctrl_rfWen),
    .io_out_bits_ctrl_rfDest(isu_io_out_bits_ctrl_rfDest),
    .io_out_bits_ctrl_isNutCoreTrap(isu_io_out_bits_ctrl_isNutCoreTrap),
    .io_out_bits_data_src1(isu_io_out_bits_data_src1),
    .io_out_bits_data_src2(isu_io_out_bits_data_src2),
    .io_out_bits_data_imm(isu_io_out_bits_data_imm),
    .io_wb_rfWen(isu_io_wb_rfWen),
    .io_wb_rfDest(isu_io_wb_rfDest),
    .io_wb_rfData(isu_io_wb_rfData),
    .io_forward_valid(isu_io_forward_valid),
    .io_forward_wb_rfWen(isu_io_forward_wb_rfWen),
    .io_forward_wb_rfDest(isu_io_forward_wb_rfDest),
    .io_forward_wb_rfData(isu_io_forward_wb_rfData),
    .io_forward_fuType(isu_io_forward_fuType),
    .io_flush(isu_io_flush),
    ._WIRE_1_0(isu__WIRE_1_0),
    .DISPLAY_ENABLE(isu_DISPLAY_ENABLE),
    ._WIRE_8(isu__WIRE_8),
    ._WIRE_2_2(isu__WIRE_2_2)
  );
  EXU exu ( // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
    .clock(exu_clock),
    .reset(exu_reset),
    .io__in_ready(exu_io__in_ready),
    .io__in_valid(exu_io__in_valid),
    .io__in_bits_cf_instr(exu_io__in_bits_cf_instr),
    .io__in_bits_cf_pc(exu_io__in_bits_cf_pc),
    .io__in_bits_cf_pnpc(exu_io__in_bits_cf_pnpc),
    .io__in_bits_cf_exceptionVec_1(exu_io__in_bits_cf_exceptionVec_1),
    .io__in_bits_cf_exceptionVec_2(exu_io__in_bits_cf_exceptionVec_2),
    .io__in_bits_cf_exceptionVec_12(exu_io__in_bits_cf_exceptionVec_12),
    .io__in_bits_cf_intrVec_0(exu_io__in_bits_cf_intrVec_0),
    .io__in_bits_cf_intrVec_1(exu_io__in_bits_cf_intrVec_1),
    .io__in_bits_cf_intrVec_2(exu_io__in_bits_cf_intrVec_2),
    .io__in_bits_cf_intrVec_3(exu_io__in_bits_cf_intrVec_3),
    .io__in_bits_cf_intrVec_4(exu_io__in_bits_cf_intrVec_4),
    .io__in_bits_cf_intrVec_5(exu_io__in_bits_cf_intrVec_5),
    .io__in_bits_cf_intrVec_6(exu_io__in_bits_cf_intrVec_6),
    .io__in_bits_cf_intrVec_7(exu_io__in_bits_cf_intrVec_7),
    .io__in_bits_cf_intrVec_8(exu_io__in_bits_cf_intrVec_8),
    .io__in_bits_cf_intrVec_9(exu_io__in_bits_cf_intrVec_9),
    .io__in_bits_cf_intrVec_10(exu_io__in_bits_cf_intrVec_10),
    .io__in_bits_cf_intrVec_11(exu_io__in_bits_cf_intrVec_11),
    .io__in_bits_cf_brIdx(exu_io__in_bits_cf_brIdx),
    .io__in_bits_cf_crossPageIPFFix(exu_io__in_bits_cf_crossPageIPFFix),
    .io__in_bits_ctrl_fuType(exu_io__in_bits_ctrl_fuType),
    .io__in_bits_ctrl_fuOpType(exu_io__in_bits_ctrl_fuOpType),
    .io__in_bits_ctrl_rfWen(exu_io__in_bits_ctrl_rfWen),
    .io__in_bits_ctrl_rfDest(exu_io__in_bits_ctrl_rfDest),
    .io__in_bits_ctrl_isNutCoreTrap(exu_io__in_bits_ctrl_isNutCoreTrap),
    .io__in_bits_data_src1(exu_io__in_bits_data_src1),
    .io__in_bits_data_src2(exu_io__in_bits_data_src2),
    .io__in_bits_data_imm(exu_io__in_bits_data_imm),
    .io__out_ready(exu_io__out_ready),
    .io__out_valid(exu_io__out_valid),
    .io__out_bits_decode_cf_instr(exu_io__out_bits_decode_cf_instr),
    .io__out_bits_decode_cf_pc(exu_io__out_bits_decode_cf_pc),
    .io__out_bits_decode_cf_redirect_target(exu_io__out_bits_decode_cf_redirect_target),
    .io__out_bits_decode_cf_redirect_valid(exu_io__out_bits_decode_cf_redirect_valid),
    .io__out_bits_decode_ctrl_fuType(exu_io__out_bits_decode_ctrl_fuType),
    .io__out_bits_decode_ctrl_rfWen(exu_io__out_bits_decode_ctrl_rfWen),
    .io__out_bits_decode_ctrl_rfDest(exu_io__out_bits_decode_ctrl_rfDest),
    .io__out_bits_isMMIO(exu_io__out_bits_isMMIO),
    .io__out_bits_intrNO(exu_io__out_bits_intrNO),
    .io__out_bits_commits_0(exu_io__out_bits_commits_0),
    .io__out_bits_commits_1(exu_io__out_bits_commits_1),
    .io__out_bits_commits_2(exu_io__out_bits_commits_2),
    .io__out_bits_commits_3(exu_io__out_bits_commits_3),
    .io__flush(exu_io__flush),
    .io__dmem_req_ready(exu_io__dmem_req_ready),
    .io__dmem_req_valid(exu_io__dmem_req_valid),
    .io__dmem_req_bits_addr(exu_io__dmem_req_bits_addr),
    .io__dmem_req_bits_size(exu_io__dmem_req_bits_size),
    .io__dmem_req_bits_cmd(exu_io__dmem_req_bits_cmd),
    .io__dmem_req_bits_wmask(exu_io__dmem_req_bits_wmask),
    .io__dmem_req_bits_wdata(exu_io__dmem_req_bits_wdata),
    .io__dmem_resp_valid(exu_io__dmem_resp_valid),
    .io__dmem_resp_bits_rdata(exu_io__dmem_resp_bits_rdata),
    .io__forward_valid(exu_io__forward_valid),
    .io__forward_wb_rfWen(exu_io__forward_wb_rfWen),
    .io__forward_wb_rfDest(exu_io__forward_wb_rfDest),
    .io__forward_wb_rfData(exu_io__forward_wb_rfData),
    .io__forward_fuType(exu_io__forward_fuType),
    .io__memMMU_imem_priviledgeMode(exu_io__memMMU_imem_priviledgeMode),
    .io__memMMU_dmem_priviledgeMode(exu_io__memMMU_dmem_priviledgeMode),
    .io__memMMU_dmem_status_sum(exu_io__memMMU_dmem_status_sum),
    .io__memMMU_dmem_status_mxr(exu_io__memMMU_dmem_status_mxr),
    .io__memMMU_dmem_loadPF(exu_io__memMMU_dmem_loadPF),
    .io__memMMU_dmem_storePF(exu_io__memMMU_dmem_storePF),
    .io__memMMU_dmem_addr(exu_io__memMMU_dmem_addr),
    .io_extra_meip_0(exu_io_extra_meip_0),
    .REG_valid(exu_REG_valid),
    .REG_pc(exu_REG_pc),
    .REG_isMissPredict(exu_REG_isMissPredict),
    .REG_actualTarget(exu_REG_actualTarget),
    .REG_actualTaken(exu_REG_actualTaken),
    .REG_fuOpType(exu_REG_fuOpType),
    .REG_btbType(exu_REG_btbType),
    .REG_isRVC(exu_REG_isRVC),
    ._WIRE_6(exu__WIRE_6),
    ._WIRE_1_0(exu__WIRE_1_0),
    .satp(exu_satp),
    .DISPLAY_ENABLE(exu_DISPLAY_ENABLE),
    ._WIRE_1_1(exu__WIRE_1_1),
    ._WIRE_8(exu__WIRE_8),
    ._WIRE_11(exu__WIRE_11),
    ._WIRE_2_2(exu__WIRE_2_2),
    .io_extra_mtip(exu_io_extra_mtip),
    ._WIRE_12(exu__WIRE_12),
    .falseWire(exu_falseWire),
    ._WIRE_1_4(exu__WIRE_1_4),
    ._WIRE_14(exu__WIRE_14),
    ._WIRE_2_3(exu__WIRE_2_3),
    ._WIRE_16(exu__WIRE_16),
    ._WIRE_17(exu__WIRE_17),
    .r_0(exu_r_0),
    .io_extra_msip(exu_io_extra_msip),
    .io_in_valid(exu_io_in_valid)
  );
  WBU wbu ( // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
    .clock(wbu_clock),
    .reset(wbu_reset),
    .io__in_valid(wbu_io__in_valid),
    .io__in_bits_decode_cf_instr(wbu_io__in_bits_decode_cf_instr),
    .io__in_bits_decode_cf_pc(wbu_io__in_bits_decode_cf_pc),
    .io__in_bits_decode_cf_redirect_target(wbu_io__in_bits_decode_cf_redirect_target),
    .io__in_bits_decode_cf_redirect_valid(wbu_io__in_bits_decode_cf_redirect_valid),
    .io__in_bits_decode_ctrl_fuType(wbu_io__in_bits_decode_ctrl_fuType),
    .io__in_bits_decode_ctrl_rfWen(wbu_io__in_bits_decode_ctrl_rfWen),
    .io__in_bits_decode_ctrl_rfDest(wbu_io__in_bits_decode_ctrl_rfDest),
    .io__in_bits_isMMIO(wbu_io__in_bits_isMMIO),
    .io__in_bits_intrNO(wbu_io__in_bits_intrNO),
    .io__in_bits_commits_0(wbu_io__in_bits_commits_0),
    .io__in_bits_commits_1(wbu_io__in_bits_commits_1),
    .io__in_bits_commits_2(wbu_io__in_bits_commits_2),
    .io__in_bits_commits_3(wbu_io__in_bits_commits_3),
    .io__wb_rfWen(wbu_io__wb_rfWen),
    .io__wb_rfDest(wbu_io__wb_rfDest),
    .io__wb_rfData(wbu_io__wb_rfData),
    .io__redirect_target(wbu_io__redirect_target),
    .io__redirect_valid(wbu_io__redirect_valid),
    .DISPLAY_ENABLE(wbu_DISPLAY_ENABLE),
    .falseWire_0(wbu_falseWire_0),
    .io_in_valid(wbu_io_in_valid)
  );
  assign io_in_0_ready = isu_io_in_0_ready; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 685:13]
  assign io_dmem_req_valid = exu_io__dmem_req_valid; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 697:11]
  assign io_dmem_req_bits_addr = exu_io__dmem_req_bits_addr; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 697:11]
  assign io_dmem_req_bits_size = exu_io__dmem_req_bits_size; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 697:11]
  assign io_dmem_req_bits_cmd = exu_io__dmem_req_bits_cmd; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 697:11]
  assign io_dmem_req_bits_wmask = exu_io__dmem_req_bits_wmask; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 697:11]
  assign io_dmem_req_bits_wdata = exu_io__dmem_req_bits_wdata; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 697:11]
  assign io_memMMU_imem_priviledgeMode = exu_io__memMMU_imem_priviledgeMode; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 695:18]
  assign io_memMMU_dmem_priviledgeMode = exu_io__memMMU_dmem_priviledgeMode; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 696:18]
  assign io_memMMU_dmem_status_sum = exu_io__memMMU_dmem_status_sum; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 696:18]
  assign io_memMMU_dmem_status_mxr = exu_io__memMMU_dmem_status_mxr; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 696:18]
  assign io_redirect_target = wbu_io__redirect_target; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 691:15]
  assign io_redirect_valid = wbu_io__redirect_valid; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 691:15]
  assign REG_valid = exu_REG_valid;
  assign REG_pc = exu_REG_pc;
  assign REG_isMissPredict = exu_REG_isMissPredict;
  assign REG_actualTarget = exu_REG_actualTarget;
  assign REG_actualTaken = exu_REG_actualTaken;
  assign REG_fuOpType = exu_REG_fuOpType;
  assign REG_btbType = exu_REG_btbType;
  assign REG_isRVC = exu_REG_isRVC;
  assign _WIRE_1 = exu__WIRE_6;
  assign satp = exu_satp;
  assign _WIRE_11 = exu__WIRE_12;
  assign _WIRE_1_4 = exu__WIRE_1_4;
  assign _WIRE_14 = exu__WIRE_14;
  assign isu_clock = clock;
  assign isu_reset = reset;
  assign isu_io_in_0_valid = io_in_0_valid; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 685:13]
  assign isu_io_in_0_bits_cf_instr = io_in_0_bits_cf_instr; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 685:13]
  assign isu_io_in_0_bits_cf_pc = io_in_0_bits_cf_pc; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 685:13]
  assign isu_io_in_0_bits_cf_pnpc = io_in_0_bits_cf_pnpc; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 685:13]
  assign isu_io_in_0_bits_cf_exceptionVec_1 = io_in_0_bits_cf_exceptionVec_1; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 685:13]
  assign isu_io_in_0_bits_cf_exceptionVec_2 = io_in_0_bits_cf_exceptionVec_2; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 685:13]
  assign isu_io_in_0_bits_cf_exceptionVec_12 = io_in_0_bits_cf_exceptionVec_12; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 685:13]
  assign isu_io_in_0_bits_cf_intrVec_0 = io_in_0_bits_cf_intrVec_0; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 685:13]
  assign isu_io_in_0_bits_cf_intrVec_1 = io_in_0_bits_cf_intrVec_1; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 685:13]
  assign isu_io_in_0_bits_cf_intrVec_2 = io_in_0_bits_cf_intrVec_2; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 685:13]
  assign isu_io_in_0_bits_cf_intrVec_3 = io_in_0_bits_cf_intrVec_3; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 685:13]
  assign isu_io_in_0_bits_cf_intrVec_4 = io_in_0_bits_cf_intrVec_4; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 685:13]
  assign isu_io_in_0_bits_cf_intrVec_5 = io_in_0_bits_cf_intrVec_5; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 685:13]
  assign isu_io_in_0_bits_cf_intrVec_6 = io_in_0_bits_cf_intrVec_6; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 685:13]
  assign isu_io_in_0_bits_cf_intrVec_7 = io_in_0_bits_cf_intrVec_7; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 685:13]
  assign isu_io_in_0_bits_cf_intrVec_8 = io_in_0_bits_cf_intrVec_8; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 685:13]
  assign isu_io_in_0_bits_cf_intrVec_9 = io_in_0_bits_cf_intrVec_9; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 685:13]
  assign isu_io_in_0_bits_cf_intrVec_10 = io_in_0_bits_cf_intrVec_10; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 685:13]
  assign isu_io_in_0_bits_cf_intrVec_11 = io_in_0_bits_cf_intrVec_11; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 685:13]
  assign isu_io_in_0_bits_cf_brIdx = io_in_0_bits_cf_brIdx; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 685:13]
  assign isu_io_in_0_bits_cf_crossPageIPFFix = io_in_0_bits_cf_crossPageIPFFix; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 685:13]
  assign isu_io_in_0_bits_ctrl_src1Type = io_in_0_bits_ctrl_src1Type; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 685:13]
  assign isu_io_in_0_bits_ctrl_src2Type = io_in_0_bits_ctrl_src2Type; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 685:13]
  assign isu_io_in_0_bits_ctrl_fuType = io_in_0_bits_ctrl_fuType; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 685:13]
  assign isu_io_in_0_bits_ctrl_fuOpType = io_in_0_bits_ctrl_fuOpType; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 685:13]
  assign isu_io_in_0_bits_ctrl_rfSrc1 = io_in_0_bits_ctrl_rfSrc1; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 685:13]
  assign isu_io_in_0_bits_ctrl_rfSrc2 = io_in_0_bits_ctrl_rfSrc2; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 685:13]
  assign isu_io_in_0_bits_ctrl_rfWen = io_in_0_bits_ctrl_rfWen; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 685:13]
  assign isu_io_in_0_bits_ctrl_rfDest = io_in_0_bits_ctrl_rfDest; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 685:13]
  assign isu_io_in_0_bits_ctrl_isNutCoreTrap = io_in_0_bits_ctrl_isNutCoreTrap; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 685:13]
  assign isu_io_in_0_bits_data_imm = io_in_0_bits_data_imm; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 685:13]
  assign isu_io_out_ready = exu_io__in_ready; // @[src/main/scala/utils/Pipeline.scala 29:16]
  assign isu_io_wb_rfWen = wbu_io__wb_rfWen; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 690:13]
  assign isu_io_wb_rfDest = wbu_io__wb_rfDest; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 690:13]
  assign isu_io_wb_rfData = wbu_io__wb_rfData; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 690:13]
  assign isu_io_forward_valid = exu_io__forward_valid; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 693:18]
  assign isu_io_forward_wb_rfWen = exu_io__forward_wb_rfWen; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 693:18]
  assign isu_io_forward_wb_rfDest = exu_io__forward_wb_rfDest; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 693:18]
  assign isu_io_forward_wb_rfData = exu_io__forward_wb_rfData; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 693:18]
  assign isu_io_forward_fuType = exu_io__forward_fuType; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 693:18]
  assign isu_io_flush = io_flush[0]; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 687:27]
  assign isu_DISPLAY_ENABLE = _WIRE_4;
  assign exu_clock = clock;
  assign exu_reset = reset;
  assign exu_io__in_valid = valid; // @[src/main/scala/utils/Pipeline.scala 31:17]
  assign exu_io__in_bits_cf_instr = exu_io_in_bits_r_cf_instr; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign exu_io__in_bits_cf_pc = exu_io_in_bits_r_cf_pc; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign exu_io__in_bits_cf_pnpc = exu_io_in_bits_r_cf_pnpc; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign exu_io__in_bits_cf_exceptionVec_1 = exu_io_in_bits_r_cf_exceptionVec_1; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign exu_io__in_bits_cf_exceptionVec_2 = exu_io_in_bits_r_cf_exceptionVec_2; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign exu_io__in_bits_cf_exceptionVec_12 = exu_io_in_bits_r_cf_exceptionVec_12; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign exu_io__in_bits_cf_intrVec_0 = exu_io_in_bits_r_cf_intrVec_0; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign exu_io__in_bits_cf_intrVec_1 = exu_io_in_bits_r_cf_intrVec_1; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign exu_io__in_bits_cf_intrVec_2 = exu_io_in_bits_r_cf_intrVec_2; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign exu_io__in_bits_cf_intrVec_3 = exu_io_in_bits_r_cf_intrVec_3; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign exu_io__in_bits_cf_intrVec_4 = exu_io_in_bits_r_cf_intrVec_4; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign exu_io__in_bits_cf_intrVec_5 = exu_io_in_bits_r_cf_intrVec_5; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign exu_io__in_bits_cf_intrVec_6 = exu_io_in_bits_r_cf_intrVec_6; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign exu_io__in_bits_cf_intrVec_7 = exu_io_in_bits_r_cf_intrVec_7; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign exu_io__in_bits_cf_intrVec_8 = exu_io_in_bits_r_cf_intrVec_8; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign exu_io__in_bits_cf_intrVec_9 = exu_io_in_bits_r_cf_intrVec_9; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign exu_io__in_bits_cf_intrVec_10 = exu_io_in_bits_r_cf_intrVec_10; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign exu_io__in_bits_cf_intrVec_11 = exu_io_in_bits_r_cf_intrVec_11; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign exu_io__in_bits_cf_brIdx = exu_io_in_bits_r_cf_brIdx; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign exu_io__in_bits_cf_crossPageIPFFix = exu_io_in_bits_r_cf_crossPageIPFFix; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign exu_io__in_bits_ctrl_fuType = exu_io_in_bits_r_ctrl_fuType; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign exu_io__in_bits_ctrl_fuOpType = exu_io_in_bits_r_ctrl_fuOpType; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign exu_io__in_bits_ctrl_rfWen = exu_io_in_bits_r_ctrl_rfWen; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign exu_io__in_bits_ctrl_rfDest = exu_io_in_bits_r_ctrl_rfDest; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign exu_io__in_bits_ctrl_isNutCoreTrap = exu_io_in_bits_r_ctrl_isNutCoreTrap; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign exu_io__in_bits_data_src1 = exu_io_in_bits_r_data_src1; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign exu_io__in_bits_data_src2 = exu_io_in_bits_r_data_src2; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign exu_io__in_bits_data_imm = exu_io_in_bits_r_data_imm; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign exu_io__out_ready = 1'h1; // @[src/main/scala/utils/Pipeline.scala 29:16]
  assign exu_io__flush = io_flush[1]; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 688:27]
  assign exu_io__dmem_req_ready = io_dmem_req_ready; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 697:11]
  assign exu_io__dmem_resp_valid = io_dmem_resp_valid; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 697:11]
  assign exu_io__dmem_resp_bits_rdata = io_dmem_resp_bits_rdata; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 697:11]
  assign exu_io__memMMU_dmem_loadPF = io_memMMU_dmem_loadPF; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 696:18]
  assign exu_io__memMMU_dmem_storePF = io_memMMU_dmem_storePF; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 696:18]
  assign exu_io__memMMU_dmem_addr = io_memMMU_dmem_addr; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 696:18]
  assign exu_io_extra_meip_0 = io_extra_meip_0;
  assign exu__WIRE_1_0 = isu__WIRE_1_0;
  assign exu_DISPLAY_ENABLE = _WIRE_4;
  assign exu__WIRE_1_1 = _WIRE_1_1;
  assign exu__WIRE_8 = _WIRE_7;
  assign exu__WIRE_11 = isu__WIRE_8;
  assign exu__WIRE_2_2 = isu__WIRE_2_2;
  assign exu_io_extra_mtip = io_extra_mtip;
  assign exu_falseWire = wbu_falseWire_0;
  assign exu__WIRE_2_3 = _WIRE_2_2;
  assign exu__WIRE_16 = _WIRE_16;
  assign exu__WIRE_17 = _WIRE_17;
  assign exu_r_0 = r_0;
  assign exu_io_extra_msip = io_extra_msip;
  assign exu_io_in_valid = wbu_io_in_valid;
  assign wbu_clock = clock;
  assign wbu_reset = reset;
  assign wbu_io__in_valid = valid_1; // @[src/main/scala/utils/Pipeline.scala 31:17]
  assign wbu_io__in_bits_decode_cf_instr = wbu_io_in_bits_r_decode_cf_instr; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign wbu_io__in_bits_decode_cf_pc = wbu_io_in_bits_r_decode_cf_pc; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign wbu_io__in_bits_decode_cf_redirect_target = wbu_io_in_bits_r_decode_cf_redirect_target; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign wbu_io__in_bits_decode_cf_redirect_valid = wbu_io_in_bits_r_decode_cf_redirect_valid; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign wbu_io__in_bits_decode_ctrl_fuType = wbu_io_in_bits_r_decode_ctrl_fuType; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign wbu_io__in_bits_decode_ctrl_rfWen = wbu_io_in_bits_r_decode_ctrl_rfWen; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign wbu_io__in_bits_decode_ctrl_rfDest = wbu_io_in_bits_r_decode_ctrl_rfDest; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign wbu_io__in_bits_isMMIO = wbu_io_in_bits_r_isMMIO; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign wbu_io__in_bits_intrNO = wbu_io_in_bits_r_intrNO; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign wbu_io__in_bits_commits_0 = wbu_io_in_bits_r_commits_0; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign wbu_io__in_bits_commits_1 = wbu_io_in_bits_r_commits_1; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign wbu_io__in_bits_commits_2 = wbu_io_in_bits_r_commits_2; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign wbu_io__in_bits_commits_3 = wbu_io_in_bits_r_commits_3; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign wbu_DISPLAY_ENABLE = _WIRE_4;
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/utils/Pipeline.scala 24:24]
      valid <= 1'h0; // @[src/main/scala/utils/Pipeline.scala 24:24]
    end else if (io_flush[0]) begin // @[src/main/scala/utils/Pipeline.scala 27:20]
      valid <= 1'h0; // @[src/main/scala/utils/Pipeline.scala 27:28]
    end else begin
      valid <= _GEN_1;
    end
    if (_T_2) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      exu_io_in_bits_r_cf_instr <= isu_io_out_bits_cf_instr; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_2) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      exu_io_in_bits_r_cf_pc <= isu_io_out_bits_cf_pc; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_2) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      exu_io_in_bits_r_cf_pnpc <= isu_io_out_bits_cf_pnpc; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_2) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      exu_io_in_bits_r_cf_exceptionVec_1 <= isu_io_out_bits_cf_exceptionVec_1; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_2) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      exu_io_in_bits_r_cf_exceptionVec_2 <= isu_io_out_bits_cf_exceptionVec_2; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_2) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      exu_io_in_bits_r_cf_exceptionVec_12 <= isu_io_out_bits_cf_exceptionVec_12; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_2) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      exu_io_in_bits_r_cf_intrVec_0 <= isu_io_out_bits_cf_intrVec_0; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_2) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      exu_io_in_bits_r_cf_intrVec_1 <= isu_io_out_bits_cf_intrVec_1; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_2) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      exu_io_in_bits_r_cf_intrVec_2 <= isu_io_out_bits_cf_intrVec_2; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_2) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      exu_io_in_bits_r_cf_intrVec_3 <= isu_io_out_bits_cf_intrVec_3; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_2) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      exu_io_in_bits_r_cf_intrVec_4 <= isu_io_out_bits_cf_intrVec_4; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_2) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      exu_io_in_bits_r_cf_intrVec_5 <= isu_io_out_bits_cf_intrVec_5; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_2) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      exu_io_in_bits_r_cf_intrVec_6 <= isu_io_out_bits_cf_intrVec_6; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_2) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      exu_io_in_bits_r_cf_intrVec_7 <= isu_io_out_bits_cf_intrVec_7; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_2) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      exu_io_in_bits_r_cf_intrVec_8 <= isu_io_out_bits_cf_intrVec_8; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_2) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      exu_io_in_bits_r_cf_intrVec_9 <= isu_io_out_bits_cf_intrVec_9; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_2) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      exu_io_in_bits_r_cf_intrVec_10 <= isu_io_out_bits_cf_intrVec_10; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_2) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      exu_io_in_bits_r_cf_intrVec_11 <= isu_io_out_bits_cf_intrVec_11; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_2) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      exu_io_in_bits_r_cf_brIdx <= isu_io_out_bits_cf_brIdx; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_2) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      exu_io_in_bits_r_cf_crossPageIPFFix <= isu_io_out_bits_cf_crossPageIPFFix; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_2) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      exu_io_in_bits_r_ctrl_fuType <= isu_io_out_bits_ctrl_fuType; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_2) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      exu_io_in_bits_r_ctrl_fuOpType <= isu_io_out_bits_ctrl_fuOpType; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_2) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      exu_io_in_bits_r_ctrl_rfWen <= isu_io_out_bits_ctrl_rfWen; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_2) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      exu_io_in_bits_r_ctrl_rfDest <= isu_io_out_bits_ctrl_rfDest; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_2) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      exu_io_in_bits_r_ctrl_isNutCoreTrap <= isu_io_out_bits_ctrl_isNutCoreTrap; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_2) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      exu_io_in_bits_r_data_src1 <= isu_io_out_bits_data_src1; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_2) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      exu_io_in_bits_r_data_src2 <= isu_io_out_bits_data_src2; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_2) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      exu_io_in_bits_r_data_imm <= isu_io_out_bits_data_imm; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (reset) begin // @[src/main/scala/utils/Pipeline.scala 24:24]
      valid_1 <= 1'h0; // @[src/main/scala/utils/Pipeline.scala 24:24]
    end else if (io_flush[1]) begin // @[src/main/scala/utils/Pipeline.scala 27:20]
      valid_1 <= 1'h0; // @[src/main/scala/utils/Pipeline.scala 27:28]
    end else begin
      valid_1 <= _T_4;
    end
    if (_T_4) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      wbu_io_in_bits_r_decode_cf_instr <= exu_io__out_bits_decode_cf_instr; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_4) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      wbu_io_in_bits_r_decode_cf_pc <= exu_io__out_bits_decode_cf_pc; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_4) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      wbu_io_in_bits_r_decode_cf_redirect_target <= exu_io__out_bits_decode_cf_redirect_target; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_4) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      wbu_io_in_bits_r_decode_cf_redirect_valid <= exu_io__out_bits_decode_cf_redirect_valid; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_4) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      wbu_io_in_bits_r_decode_ctrl_fuType <= exu_io__out_bits_decode_ctrl_fuType; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_4) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      wbu_io_in_bits_r_decode_ctrl_rfWen <= exu_io__out_bits_decode_ctrl_rfWen; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_4) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      wbu_io_in_bits_r_decode_ctrl_rfDest <= exu_io__out_bits_decode_ctrl_rfDest; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_4) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      wbu_io_in_bits_r_isMMIO <= exu_io__out_bits_isMMIO; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_4) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      wbu_io_in_bits_r_intrNO <= exu_io__out_bits_intrNO; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_4) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      wbu_io_in_bits_r_commits_0 <= exu_io__out_bits_commits_0; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_4) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      wbu_io_in_bits_r_commits_1 <= exu_io__out_bits_commits_1; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_4) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      wbu_io_in_bits_r_commits_2 <= exu_io__out_bits_commits_2; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_4) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      wbu_io_in_bits_r_commits_3 <= exu_io__out_bits_commits_3; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  valid = _RAND_0[0:0];
  _RAND_1 = {2{`RANDOM}};
  exu_io_in_bits_r_cf_instr = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  exu_io_in_bits_r_cf_pc = _RAND_2[38:0];
  _RAND_3 = {2{`RANDOM}};
  exu_io_in_bits_r_cf_pnpc = _RAND_3[38:0];
  _RAND_4 = {1{`RANDOM}};
  exu_io_in_bits_r_cf_exceptionVec_1 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  exu_io_in_bits_r_cf_exceptionVec_2 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  exu_io_in_bits_r_cf_exceptionVec_12 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  exu_io_in_bits_r_cf_intrVec_0 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  exu_io_in_bits_r_cf_intrVec_1 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  exu_io_in_bits_r_cf_intrVec_2 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  exu_io_in_bits_r_cf_intrVec_3 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  exu_io_in_bits_r_cf_intrVec_4 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  exu_io_in_bits_r_cf_intrVec_5 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  exu_io_in_bits_r_cf_intrVec_6 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  exu_io_in_bits_r_cf_intrVec_7 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  exu_io_in_bits_r_cf_intrVec_8 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  exu_io_in_bits_r_cf_intrVec_9 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  exu_io_in_bits_r_cf_intrVec_10 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  exu_io_in_bits_r_cf_intrVec_11 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  exu_io_in_bits_r_cf_brIdx = _RAND_19[3:0];
  _RAND_20 = {1{`RANDOM}};
  exu_io_in_bits_r_cf_crossPageIPFFix = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  exu_io_in_bits_r_ctrl_fuType = _RAND_21[2:0];
  _RAND_22 = {1{`RANDOM}};
  exu_io_in_bits_r_ctrl_fuOpType = _RAND_22[6:0];
  _RAND_23 = {1{`RANDOM}};
  exu_io_in_bits_r_ctrl_rfWen = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  exu_io_in_bits_r_ctrl_rfDest = _RAND_24[4:0];
  _RAND_25 = {1{`RANDOM}};
  exu_io_in_bits_r_ctrl_isNutCoreTrap = _RAND_25[0:0];
  _RAND_26 = {2{`RANDOM}};
  exu_io_in_bits_r_data_src1 = _RAND_26[63:0];
  _RAND_27 = {2{`RANDOM}};
  exu_io_in_bits_r_data_src2 = _RAND_27[63:0];
  _RAND_28 = {2{`RANDOM}};
  exu_io_in_bits_r_data_imm = _RAND_28[63:0];
  _RAND_29 = {1{`RANDOM}};
  valid_1 = _RAND_29[0:0];
  _RAND_30 = {2{`RANDOM}};
  wbu_io_in_bits_r_decode_cf_instr = _RAND_30[63:0];
  _RAND_31 = {2{`RANDOM}};
  wbu_io_in_bits_r_decode_cf_pc = _RAND_31[38:0];
  _RAND_32 = {2{`RANDOM}};
  wbu_io_in_bits_r_decode_cf_redirect_target = _RAND_32[38:0];
  _RAND_33 = {1{`RANDOM}};
  wbu_io_in_bits_r_decode_cf_redirect_valid = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  wbu_io_in_bits_r_decode_ctrl_fuType = _RAND_34[2:0];
  _RAND_35 = {1{`RANDOM}};
  wbu_io_in_bits_r_decode_ctrl_rfWen = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  wbu_io_in_bits_r_decode_ctrl_rfDest = _RAND_36[4:0];
  _RAND_37 = {1{`RANDOM}};
  wbu_io_in_bits_r_isMMIO = _RAND_37[0:0];
  _RAND_38 = {2{`RANDOM}};
  wbu_io_in_bits_r_intrNO = _RAND_38[63:0];
  _RAND_39 = {2{`RANDOM}};
  wbu_io_in_bits_r_commits_0 = _RAND_39[63:0];
  _RAND_40 = {2{`RANDOM}};
  wbu_io_in_bits_r_commits_1 = _RAND_40[63:0];
  _RAND_41 = {2{`RANDOM}};
  wbu_io_in_bits_r_commits_2 = _RAND_41[63:0];
  _RAND_42 = {2{`RANDOM}};
  wbu_io_in_bits_r_commits_3 = _RAND_42[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module LockingArbiter(
  input         clock,
  input         reset,
  output        io_in_0_ready, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  input         io_in_0_valid, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  input  [31:0] io_in_0_bits_addr, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  input  [3:0]  io_in_0_bits_cmd, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  input  [7:0]  io_in_0_bits_wmask, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  input  [63:0] io_in_0_bits_wdata, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  output        io_in_1_ready, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  input         io_in_1_valid, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  input  [31:0] io_in_1_bits_addr, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  input  [2:0]  io_in_1_bits_size, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  input  [3:0]  io_in_1_bits_cmd, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  input  [7:0]  io_in_1_bits_wmask, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  input  [63:0] io_in_1_bits_wdata, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  input         io_out_ready, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  output        io_out_valid, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  output [31:0] io_out_bits_addr, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  output [2:0]  io_out_bits_size, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  output [3:0]  io_out_bits_cmd, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  output [7:0]  io_out_bits_wmask, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  output [63:0] io_out_bits_wdata, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  output        io_chosen // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg [2:0] lockCount_value; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
  reg  lockIdx; // @[src/main/scala/chisel3/util/Arbiter.scala 60:22]
  wire  locked = lockCount_value != 3'h0; // @[src/main/scala/chisel3/util/Arbiter.scala 61:34]
  wire  wantsLock = io_out_bits_cmd[0] & io_out_bits_cmd[1]; // @[src/main/scala/bus/simplebus/Crossbar.scala 94:62]
  wire  _T = io_out_ready & io_out_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  wire [2:0] _value_T_1 = lockCount_value + 3'h1; // @[src/main/scala/chisel3/util/Counter.scala 77:24]
  wire  io_chosen_choice = io_in_0_valid ? 1'h0 : 1'h1; // @[src/main/scala/chisel3/util/Arbiter.scala 103:{26,35} 101:41]
  wire  _T_2 = ~io_in_0_valid; // @[src/main/scala/chisel3/util/Arbiter.scala 45:78]
  wire  _io_in_0_ready_T_1 = locked ? ~lockIdx : 1'h1; // @[src/main/scala/chisel3/util/Arbiter.scala 71:22]
  wire  _io_in_1_ready_T_1 = locked ? lockIdx : _T_2; // @[src/main/scala/chisel3/util/Arbiter.scala 71:22]
  assign io_in_0_ready = _io_in_0_ready_T_1 & io_out_ready; // @[src/main/scala/chisel3/util/Arbiter.scala 71:56]
  assign io_in_1_ready = _io_in_1_ready_T_1 & io_out_ready; // @[src/main/scala/chisel3/util/Arbiter.scala 71:56]
  assign io_out_valid = io_chosen ? io_in_1_valid : io_in_0_valid; // @[src/main/scala/chisel3/util/Arbiter.scala 55:{16,16}]
  assign io_out_bits_addr = io_chosen ? io_in_1_bits_addr : io_in_0_bits_addr; // @[src/main/scala/chisel3/util/Arbiter.scala 56:{15,15}]
  assign io_out_bits_size = io_chosen ? io_in_1_bits_size : 3'h3; // @[src/main/scala/chisel3/util/Arbiter.scala 56:{15,15}]
  assign io_out_bits_cmd = io_chosen ? io_in_1_bits_cmd : io_in_0_bits_cmd; // @[src/main/scala/chisel3/util/Arbiter.scala 56:{15,15}]
  assign io_out_bits_wmask = io_chosen ? io_in_1_bits_wmask : io_in_0_bits_wmask; // @[src/main/scala/chisel3/util/Arbiter.scala 56:{15,15}]
  assign io_out_bits_wdata = io_chosen ? io_in_1_bits_wdata : io_in_0_bits_wdata; // @[src/main/scala/chisel3/util/Arbiter.scala 56:{15,15}]
  assign io_chosen = locked ? lockIdx : io_chosen_choice; // @[src/main/scala/chisel3/util/Arbiter.scala 54:13 69:{18,30}]
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/chisel3/util/Counter.scala 61:40]
      lockCount_value <= 3'h0; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end else if (_T & wantsLock) begin // @[src/main/scala/chisel3/util/Arbiter.scala 64:36]
      lockCount_value <= _value_T_1; // @[src/main/scala/chisel3/util/Counter.scala 77:15]
    end
    if (_T & wantsLock) begin // @[src/main/scala/chisel3/util/Arbiter.scala 64:36]
      lockIdx <= io_chosen; // @[src/main/scala/chisel3/util/Arbiter.scala 65:15]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  lockCount_value = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  lockIdx = _RAND_1[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module SimpleBusCrossbarNto1(
  input         clock,
  input         reset,
  output        io_in_0_req_ready, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  input         io_in_0_req_valid, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  input  [31:0] io_in_0_req_bits_addr, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  input  [3:0]  io_in_0_req_bits_cmd, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  input  [7:0]  io_in_0_req_bits_wmask, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  input  [63:0] io_in_0_req_bits_wdata, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  output        io_in_0_resp_valid, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  output [3:0]  io_in_0_resp_bits_cmd, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  output [63:0] io_in_0_resp_bits_rdata, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  output        io_in_1_req_ready, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  input         io_in_1_req_valid, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  input  [31:0] io_in_1_req_bits_addr, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  input  [2:0]  io_in_1_req_bits_size, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  input  [3:0]  io_in_1_req_bits_cmd, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  input  [7:0]  io_in_1_req_bits_wmask, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  input  [63:0] io_in_1_req_bits_wdata, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  output        io_in_1_resp_valid, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  output [3:0]  io_in_1_resp_bits_cmd, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  output [63:0] io_in_1_resp_bits_rdata, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  input         io_out_req_ready, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  output        io_out_req_valid, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  output [31:0] io_out_req_bits_addr, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  output [2:0]  io_out_req_bits_size, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  output [3:0]  io_out_req_bits_cmd, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  output [7:0]  io_out_req_bits_wmask, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  output [63:0] io_out_req_bits_wdata, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  output        io_out_resp_ready, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  input         io_out_resp_valid, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  input  [3:0]  io_out_resp_bits_cmd, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  input  [63:0] io_out_resp_bits_rdata // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  wire  inputArb_clock; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire  inputArb_reset; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire  inputArb_io_in_0_ready; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire  inputArb_io_in_0_valid; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire [31:0] inputArb_io_in_0_bits_addr; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire [3:0] inputArb_io_in_0_bits_cmd; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire [7:0] inputArb_io_in_0_bits_wmask; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire [63:0] inputArb_io_in_0_bits_wdata; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire  inputArb_io_in_1_ready; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire  inputArb_io_in_1_valid; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire [31:0] inputArb_io_in_1_bits_addr; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire [2:0] inputArb_io_in_1_bits_size; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire [3:0] inputArb_io_in_1_bits_cmd; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire [7:0] inputArb_io_in_1_bits_wmask; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire [63:0] inputArb_io_in_1_bits_wdata; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire  inputArb_io_out_ready; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire  inputArb_io_out_valid; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire [31:0] inputArb_io_out_bits_addr; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire [2:0] inputArb_io_out_bits_size; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire [3:0] inputArb_io_out_bits_cmd; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire [7:0] inputArb_io_out_bits_wmask; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire [63:0] inputArb_io_out_bits_wdata; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire  inputArb_io_chosen; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  reg [1:0] state; // @[src/main/scala/bus/simplebus/Crossbar.scala 92:22]
  wire  _T_1 = ~inputArb_io_out_bits_cmd[0]; // @[src/main/scala/bus/simplebus/SimpleBus.scala 73:18]
  wire  _T_4 = ~inputArb_io_out_bits_cmd[0] & ~inputArb_io_out_bits_cmd[3]; // @[src/main/scala/bus/simplebus/SimpleBus.scala 73:26]
  reg  inflightSrc; // @[src/main/scala/bus/simplebus/Crossbar.scala 99:28]
  wire  _io_out_req_valid_T = state == 2'h0; // @[src/main/scala/bus/simplebus/Crossbar.scala 103:47]
  wire  _T_15 = inputArb_io_out_ready & inputArb_io_out_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  wire  _T_21 = inputArb_io_out_bits_cmd == 4'h7; // @[src/main/scala/bus/simplebus/SimpleBus.scala 78:27]
  wire  _T_22 = inputArb_io_out_bits_cmd == 4'h1; // @[src/main/scala/bus/simplebus/SimpleBus.scala 77:29]
  wire [1:0] _GEN_4 = _T_21 | _T_22 ? 2'h2 : state; // @[src/main/scala/bus/simplebus/Crossbar.scala 118:{80,88} 92:22]
  wire  _T_25 = io_out_resp_ready & io_out_resp_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  wire  _T_26 = io_out_resp_bits_cmd == 4'h6; // @[src/main/scala/bus/simplebus/SimpleBus.scala 91:24]
  wire [1:0] _GEN_9 = _T_25 ? 2'h0 : state; // @[src/main/scala/bus/simplebus/Crossbar.scala 122:{48,56} 92:22]
  LockingArbiter inputArb ( // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
    .clock(inputArb_clock),
    .reset(inputArb_reset),
    .io_in_0_ready(inputArb_io_in_0_ready),
    .io_in_0_valid(inputArb_io_in_0_valid),
    .io_in_0_bits_addr(inputArb_io_in_0_bits_addr),
    .io_in_0_bits_cmd(inputArb_io_in_0_bits_cmd),
    .io_in_0_bits_wmask(inputArb_io_in_0_bits_wmask),
    .io_in_0_bits_wdata(inputArb_io_in_0_bits_wdata),
    .io_in_1_ready(inputArb_io_in_1_ready),
    .io_in_1_valid(inputArb_io_in_1_valid),
    .io_in_1_bits_addr(inputArb_io_in_1_bits_addr),
    .io_in_1_bits_size(inputArb_io_in_1_bits_size),
    .io_in_1_bits_cmd(inputArb_io_in_1_bits_cmd),
    .io_in_1_bits_wmask(inputArb_io_in_1_bits_wmask),
    .io_in_1_bits_wdata(inputArb_io_in_1_bits_wdata),
    .io_out_ready(inputArb_io_out_ready),
    .io_out_valid(inputArb_io_out_valid),
    .io_out_bits_addr(inputArb_io_out_bits_addr),
    .io_out_bits_size(inputArb_io_out_bits_size),
    .io_out_bits_cmd(inputArb_io_out_bits_cmd),
    .io_out_bits_wmask(inputArb_io_out_bits_wmask),
    .io_out_bits_wdata(inputArb_io_out_bits_wdata),
    .io_chosen(inputArb_io_chosen)
  );
  assign io_in_0_req_ready = inputArb_io_in_0_ready; // @[src/main/scala/bus/simplebus/Crossbar.scala 96:68]
  assign io_in_0_resp_valid = ~inflightSrc & io_out_resp_valid; // @[src/main/scala/bus/simplebus/Crossbar.scala 109:{13,13} 107:26]
  assign io_in_0_resp_bits_cmd = io_out_resp_bits_cmd; // @[src/main/scala/bus/simplebus/Crossbar.scala 106:25]
  assign io_in_0_resp_bits_rdata = io_out_resp_bits_rdata; // @[src/main/scala/bus/simplebus/Crossbar.scala 106:25]
  assign io_in_1_req_ready = inputArb_io_in_1_ready; // @[src/main/scala/bus/simplebus/Crossbar.scala 96:68]
  assign io_in_1_resp_valid = inflightSrc & io_out_resp_valid; // @[src/main/scala/bus/simplebus/Crossbar.scala 109:{13,13} 107:26]
  assign io_in_1_resp_bits_cmd = io_out_resp_bits_cmd; // @[src/main/scala/bus/simplebus/Crossbar.scala 106:25]
  assign io_in_1_resp_bits_rdata = io_out_resp_bits_rdata; // @[src/main/scala/bus/simplebus/Crossbar.scala 106:25]
  assign io_out_req_valid = inputArb_io_out_valid & state == 2'h0; // @[src/main/scala/bus/simplebus/Crossbar.scala 103:37]
  assign io_out_req_bits_addr = inputArb_io_out_bits_addr; // @[src/main/scala/bus/simplebus/Crossbar.scala 101:19]
  assign io_out_req_bits_size = inputArb_io_out_bits_size; // @[src/main/scala/bus/simplebus/Crossbar.scala 101:19]
  assign io_out_req_bits_cmd = inputArb_io_out_bits_cmd; // @[src/main/scala/bus/simplebus/Crossbar.scala 101:19]
  assign io_out_req_bits_wmask = inputArb_io_out_bits_wmask; // @[src/main/scala/bus/simplebus/Crossbar.scala 101:19]
  assign io_out_req_bits_wdata = inputArb_io_out_bits_wdata; // @[src/main/scala/bus/simplebus/Crossbar.scala 101:19]
  assign io_out_resp_ready = 1'h1; // @[src/main/scala/bus/simplebus/Crossbar.scala 110:{13,13}]
  assign inputArb_clock = clock;
  assign inputArb_reset = reset;
  assign inputArb_io_in_0_valid = io_in_0_req_valid; // @[src/main/scala/bus/simplebus/Crossbar.scala 96:68]
  assign inputArb_io_in_0_bits_addr = io_in_0_req_bits_addr; // @[src/main/scala/bus/simplebus/Crossbar.scala 96:68]
  assign inputArb_io_in_0_bits_cmd = io_in_0_req_bits_cmd; // @[src/main/scala/bus/simplebus/Crossbar.scala 96:68]
  assign inputArb_io_in_0_bits_wmask = io_in_0_req_bits_wmask; // @[src/main/scala/bus/simplebus/Crossbar.scala 96:68]
  assign inputArb_io_in_0_bits_wdata = io_in_0_req_bits_wdata; // @[src/main/scala/bus/simplebus/Crossbar.scala 96:68]
  assign inputArb_io_in_1_valid = io_in_1_req_valid; // @[src/main/scala/bus/simplebus/Crossbar.scala 96:68]
  assign inputArb_io_in_1_bits_addr = io_in_1_req_bits_addr; // @[src/main/scala/bus/simplebus/Crossbar.scala 96:68]
  assign inputArb_io_in_1_bits_size = io_in_1_req_bits_size; // @[src/main/scala/bus/simplebus/Crossbar.scala 96:68]
  assign inputArb_io_in_1_bits_cmd = io_in_1_req_bits_cmd; // @[src/main/scala/bus/simplebus/Crossbar.scala 96:68]
  assign inputArb_io_in_1_bits_wmask = io_in_1_req_bits_wmask; // @[src/main/scala/bus/simplebus/Crossbar.scala 96:68]
  assign inputArb_io_in_1_bits_wdata = io_in_1_req_bits_wdata; // @[src/main/scala/bus/simplebus/Crossbar.scala 96:68]
  assign inputArb_io_out_ready = io_out_req_ready & _io_out_req_valid_T; // @[src/main/scala/bus/simplebus/Crossbar.scala 104:37]
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 92:22]
      state <= 2'h0; // @[src/main/scala/bus/simplebus/Crossbar.scala 92:22]
    end else if (2'h0 == state) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 113:18]
      if (_T_15) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 115:27]
        if (_T_4) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 117:38]
          state <= 2'h1; // @[src/main/scala/bus/simplebus/Crossbar.scala 117:46]
        end else begin
          state <= _GEN_4;
        end
      end
    end else if (2'h1 == state) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 113:18]
      if (_T_25 & _T_26) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 121:78]
        state <= 2'h0; // @[src/main/scala/bus/simplebus/Crossbar.scala 121:86]
      end
    end else if (2'h2 == state) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 113:18]
      state <= _GEN_9;
    end
    if (reset) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 99:28]
      inflightSrc <= 1'h0; // @[src/main/scala/bus/simplebus/Crossbar.scala 99:28]
    end else if (2'h0 == state) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 113:18]
      if (_T_15) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 115:27]
        inflightSrc <= inputArb_io_chosen; // @[src/main/scala/bus/simplebus/Crossbar.scala 116:21]
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~(inputArb_io_out_valid & ~_T_4 & _T_1))) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Crossbar.scala:98 assert(!(thisReq.valid && !thisReq.bits.isRead() && !thisReq.bits.isWrite()))\n"
            ); // @[src/main/scala/bus/simplebus/Crossbar.scala 98:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~(inputArb_io_out_valid & ~_T_4 & _T_1)) & ~reset) begin
          $fatal; // @[src/main/scala/bus/simplebus/Crossbar.scala 98:9]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  inflightSrc = _RAND_1[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module LockingArbiter_1(
  input         clock,
  input         reset,
  output        io_in_0_ready, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  input         io_in_0_valid, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  input  [31:0] io_in_0_bits_addr, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  input  [2:0]  io_in_0_bits_size, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  input  [3:0]  io_in_0_bits_cmd, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  input  [7:0]  io_in_0_bits_wmask, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  input  [63:0] io_in_0_bits_wdata, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  output        io_in_1_ready, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  input         io_in_1_valid, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  input  [31:0] io_in_1_bits_addr, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  input  [3:0]  io_in_1_bits_cmd, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  input  [63:0] io_in_1_bits_wdata, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  output        io_in_2_ready, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  input         io_in_2_valid, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  input  [31:0] io_in_2_bits_addr, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  input  [3:0]  io_in_2_bits_cmd, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  input  [63:0] io_in_2_bits_wdata, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  output        io_in_3_ready, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  input         io_in_3_valid, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  input  [31:0] io_in_3_bits_addr, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  input  [2:0]  io_in_3_bits_size, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  input  [3:0]  io_in_3_bits_cmd, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  input  [7:0]  io_in_3_bits_wmask, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  input  [63:0] io_in_3_bits_wdata, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  input         io_out_ready, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  output        io_out_valid, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  output [31:0] io_out_bits_addr, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  output [2:0]  io_out_bits_size, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  output [3:0]  io_out_bits_cmd, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  output [7:0]  io_out_bits_wmask, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  output [63:0] io_out_bits_wdata, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  output [1:0]  io_chosen // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  wire  _GEN_1 = 2'h1 == io_chosen ? io_in_1_valid : io_in_0_valid; // @[src/main/scala/chisel3/util/Arbiter.scala 55:{16,16}]
  wire  _GEN_2 = 2'h2 == io_chosen ? io_in_2_valid : _GEN_1; // @[src/main/scala/chisel3/util/Arbiter.scala 55:{16,16}]
  wire [31:0] _GEN_5 = 2'h1 == io_chosen ? io_in_1_bits_addr : io_in_0_bits_addr; // @[src/main/scala/chisel3/util/Arbiter.scala 56:{15,15}]
  wire [31:0] _GEN_6 = 2'h2 == io_chosen ? io_in_2_bits_addr : _GEN_5; // @[src/main/scala/chisel3/util/Arbiter.scala 56:{15,15}]
  wire [2:0] _GEN_9 = 2'h1 == io_chosen ? 3'h3 : io_in_0_bits_size; // @[src/main/scala/chisel3/util/Arbiter.scala 56:{15,15}]
  wire [2:0] _GEN_10 = 2'h2 == io_chosen ? 3'h3 : _GEN_9; // @[src/main/scala/chisel3/util/Arbiter.scala 56:{15,15}]
  wire [3:0] _GEN_13 = 2'h1 == io_chosen ? io_in_1_bits_cmd : io_in_0_bits_cmd; // @[src/main/scala/chisel3/util/Arbiter.scala 56:{15,15}]
  wire [3:0] _GEN_14 = 2'h2 == io_chosen ? io_in_2_bits_cmd : _GEN_13; // @[src/main/scala/chisel3/util/Arbiter.scala 56:{15,15}]
  wire [7:0] _GEN_17 = 2'h1 == io_chosen ? 8'hff : io_in_0_bits_wmask; // @[src/main/scala/chisel3/util/Arbiter.scala 56:{15,15}]
  wire [7:0] _GEN_18 = 2'h2 == io_chosen ? 8'hff : _GEN_17; // @[src/main/scala/chisel3/util/Arbiter.scala 56:{15,15}]
  wire [63:0] _GEN_21 = 2'h1 == io_chosen ? io_in_1_bits_wdata : io_in_0_bits_wdata; // @[src/main/scala/chisel3/util/Arbiter.scala 56:{15,15}]
  wire [63:0] _GEN_22 = 2'h2 == io_chosen ? io_in_2_bits_wdata : _GEN_21; // @[src/main/scala/chisel3/util/Arbiter.scala 56:{15,15}]
  reg [2:0] lockCount_value; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
  reg [1:0] lockIdx; // @[src/main/scala/chisel3/util/Arbiter.scala 60:22]
  wire  locked = lockCount_value != 3'h0; // @[src/main/scala/chisel3/util/Arbiter.scala 61:34]
  wire  wantsLock = io_out_bits_cmd[0] & io_out_bits_cmd[1]; // @[src/main/scala/bus/simplebus/Crossbar.scala 94:62]
  wire  _T = io_out_ready & io_out_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  wire [2:0] _value_T_1 = lockCount_value + 3'h1; // @[src/main/scala/chisel3/util/Counter.scala 77:24]
  wire [1:0] _GEN_27 = io_in_2_valid ? 2'h2 : 2'h3; // @[src/main/scala/chisel3/util/Arbiter.scala 103:{26,35} 101:41]
  wire [1:0] _GEN_28 = io_in_1_valid ? 2'h1 : _GEN_27; // @[src/main/scala/chisel3/util/Arbiter.scala 103:{26,35}]
  wire [1:0] io_chosen_choice = io_in_0_valid ? 2'h0 : _GEN_28; // @[src/main/scala/chisel3/util/Arbiter.scala 103:{26,35}]
  wire  _T_4 = ~io_in_0_valid; // @[src/main/scala/chisel3/util/Arbiter.scala 45:78]
  wire  _T_5 = ~(io_in_0_valid | io_in_1_valid); // @[src/main/scala/chisel3/util/Arbiter.scala 45:78]
  wire  _T_6 = ~(io_in_0_valid | io_in_1_valid | io_in_2_valid); // @[src/main/scala/chisel3/util/Arbiter.scala 45:78]
  wire  _io_in_0_ready_T_1 = locked ? lockIdx == 2'h0 : 1'h1; // @[src/main/scala/chisel3/util/Arbiter.scala 71:22]
  wire  _io_in_1_ready_T_1 = locked ? lockIdx == 2'h1 : _T_4; // @[src/main/scala/chisel3/util/Arbiter.scala 71:22]
  wire  _io_in_2_ready_T_1 = locked ? lockIdx == 2'h2 : _T_5; // @[src/main/scala/chisel3/util/Arbiter.scala 71:22]
  wire  _io_in_3_ready_T_1 = locked ? lockIdx == 2'h3 : _T_6; // @[src/main/scala/chisel3/util/Arbiter.scala 71:22]
  assign io_in_0_ready = _io_in_0_ready_T_1 & io_out_ready; // @[src/main/scala/chisel3/util/Arbiter.scala 71:56]
  assign io_in_1_ready = _io_in_1_ready_T_1 & io_out_ready; // @[src/main/scala/chisel3/util/Arbiter.scala 71:56]
  assign io_in_2_ready = _io_in_2_ready_T_1 & io_out_ready; // @[src/main/scala/chisel3/util/Arbiter.scala 71:56]
  assign io_in_3_ready = _io_in_3_ready_T_1 & io_out_ready; // @[src/main/scala/chisel3/util/Arbiter.scala 71:56]
  assign io_out_valid = 2'h3 == io_chosen ? io_in_3_valid : _GEN_2; // @[src/main/scala/chisel3/util/Arbiter.scala 55:{16,16}]
  assign io_out_bits_addr = 2'h3 == io_chosen ? io_in_3_bits_addr : _GEN_6; // @[src/main/scala/chisel3/util/Arbiter.scala 56:{15,15}]
  assign io_out_bits_size = 2'h3 == io_chosen ? io_in_3_bits_size : _GEN_10; // @[src/main/scala/chisel3/util/Arbiter.scala 56:{15,15}]
  assign io_out_bits_cmd = 2'h3 == io_chosen ? io_in_3_bits_cmd : _GEN_14; // @[src/main/scala/chisel3/util/Arbiter.scala 56:{15,15}]
  assign io_out_bits_wmask = 2'h3 == io_chosen ? io_in_3_bits_wmask : _GEN_18; // @[src/main/scala/chisel3/util/Arbiter.scala 56:{15,15}]
  assign io_out_bits_wdata = 2'h3 == io_chosen ? io_in_3_bits_wdata : _GEN_22; // @[src/main/scala/chisel3/util/Arbiter.scala 56:{15,15}]
  assign io_chosen = locked ? lockIdx : io_chosen_choice; // @[src/main/scala/chisel3/util/Arbiter.scala 54:13 69:{18,30}]
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/chisel3/util/Counter.scala 61:40]
      lockCount_value <= 3'h0; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end else if (_T & wantsLock) begin // @[src/main/scala/chisel3/util/Arbiter.scala 64:36]
      lockCount_value <= _value_T_1; // @[src/main/scala/chisel3/util/Counter.scala 77:15]
    end
    if (_T & wantsLock) begin // @[src/main/scala/chisel3/util/Arbiter.scala 64:36]
      lockIdx <= io_chosen; // @[src/main/scala/chisel3/util/Arbiter.scala 65:15]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  lockCount_value = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  lockIdx = _RAND_1[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module SimpleBusCrossbarNto1_1(
  input         clock,
  input         reset,
  output        io_in_0_req_ready, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  input         io_in_0_req_valid, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  input  [31:0] io_in_0_req_bits_addr, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  input  [2:0]  io_in_0_req_bits_size, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  input  [3:0]  io_in_0_req_bits_cmd, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  input  [7:0]  io_in_0_req_bits_wmask, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  input  [63:0] io_in_0_req_bits_wdata, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  output        io_in_0_resp_valid, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  output [3:0]  io_in_0_resp_bits_cmd, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  output [63:0] io_in_0_resp_bits_rdata, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  output        io_in_1_req_ready, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  input         io_in_1_req_valid, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  input  [31:0] io_in_1_req_bits_addr, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  input  [3:0]  io_in_1_req_bits_cmd, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  input  [63:0] io_in_1_req_bits_wdata, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  output        io_in_1_resp_valid, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  output [3:0]  io_in_1_resp_bits_cmd, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  output [63:0] io_in_1_resp_bits_rdata, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  output        io_in_2_req_ready, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  input         io_in_2_req_valid, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  input  [31:0] io_in_2_req_bits_addr, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  input  [3:0]  io_in_2_req_bits_cmd, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  input  [63:0] io_in_2_req_bits_wdata, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  output        io_in_2_resp_valid, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  output [3:0]  io_in_2_resp_bits_cmd, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  output [63:0] io_in_2_resp_bits_rdata, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  output        io_in_3_req_ready, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  input         io_in_3_req_valid, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  input  [31:0] io_in_3_req_bits_addr, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  input  [2:0]  io_in_3_req_bits_size, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  input  [3:0]  io_in_3_req_bits_cmd, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  input  [7:0]  io_in_3_req_bits_wmask, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  input  [63:0] io_in_3_req_bits_wdata, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  input         io_in_3_resp_ready, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  output        io_in_3_resp_valid, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  output [3:0]  io_in_3_resp_bits_cmd, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  output [63:0] io_in_3_resp_bits_rdata, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  input         io_out_req_ready, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  output        io_out_req_valid, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  output [31:0] io_out_req_bits_addr, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  output [2:0]  io_out_req_bits_size, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  output [3:0]  io_out_req_bits_cmd, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  output [7:0]  io_out_req_bits_wmask, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  output [63:0] io_out_req_bits_wdata, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  output        io_out_resp_ready, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  input         io_out_resp_valid, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  input  [3:0]  io_out_resp_bits_cmd, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  input  [63:0] io_out_resp_bits_rdata // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  wire  inputArb_clock; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire  inputArb_reset; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire  inputArb_io_in_0_ready; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire  inputArb_io_in_0_valid; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire [31:0] inputArb_io_in_0_bits_addr; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire [2:0] inputArb_io_in_0_bits_size; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire [3:0] inputArb_io_in_0_bits_cmd; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire [7:0] inputArb_io_in_0_bits_wmask; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire [63:0] inputArb_io_in_0_bits_wdata; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire  inputArb_io_in_1_ready; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire  inputArb_io_in_1_valid; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire [31:0] inputArb_io_in_1_bits_addr; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire [3:0] inputArb_io_in_1_bits_cmd; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire [63:0] inputArb_io_in_1_bits_wdata; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire  inputArb_io_in_2_ready; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire  inputArb_io_in_2_valid; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire [31:0] inputArb_io_in_2_bits_addr; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire [3:0] inputArb_io_in_2_bits_cmd; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire [63:0] inputArb_io_in_2_bits_wdata; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire  inputArb_io_in_3_ready; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire  inputArb_io_in_3_valid; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire [31:0] inputArb_io_in_3_bits_addr; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire [2:0] inputArb_io_in_3_bits_size; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire [3:0] inputArb_io_in_3_bits_cmd; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire [7:0] inputArb_io_in_3_bits_wmask; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire [63:0] inputArb_io_in_3_bits_wdata; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire  inputArb_io_out_ready; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire  inputArb_io_out_valid; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire [31:0] inputArb_io_out_bits_addr; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire [2:0] inputArb_io_out_bits_size; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire [3:0] inputArb_io_out_bits_cmd; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire [7:0] inputArb_io_out_bits_wmask; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire [63:0] inputArb_io_out_bits_wdata; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire [1:0] inputArb_io_chosen; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  reg [1:0] state; // @[src/main/scala/bus/simplebus/Crossbar.scala 92:22]
  wire  _T_1 = ~inputArb_io_out_bits_cmd[0]; // @[src/main/scala/bus/simplebus/SimpleBus.scala 73:18]
  wire  _T_4 = ~inputArb_io_out_bits_cmd[0] & ~inputArb_io_out_bits_cmd[3]; // @[src/main/scala/bus/simplebus/SimpleBus.scala 73:26]
  reg [1:0] inflightSrc; // @[src/main/scala/bus/simplebus/Crossbar.scala 99:28]
  wire  _io_out_req_valid_T = state == 2'h0; // @[src/main/scala/bus/simplebus/Crossbar.scala 103:47]
  wire  _T_15 = inputArb_io_out_ready & inputArb_io_out_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  wire  _T_21 = inputArb_io_out_bits_cmd == 4'h7; // @[src/main/scala/bus/simplebus/SimpleBus.scala 78:27]
  wire  _T_22 = inputArb_io_out_bits_cmd == 4'h1; // @[src/main/scala/bus/simplebus/SimpleBus.scala 77:29]
  wire [1:0] _GEN_8 = _T_21 | _T_22 ? 2'h2 : state; // @[src/main/scala/bus/simplebus/Crossbar.scala 118:{80,88} 92:22]
  wire  _T_25 = io_out_resp_ready & io_out_resp_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  wire  _T_26 = io_out_resp_bits_cmd == 4'h6; // @[src/main/scala/bus/simplebus/SimpleBus.scala 91:24]
  wire [1:0] _GEN_13 = _T_25 ? 2'h0 : state; // @[src/main/scala/bus/simplebus/Crossbar.scala 122:{48,56} 92:22]
  LockingArbiter_1 inputArb ( // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
    .clock(inputArb_clock),
    .reset(inputArb_reset),
    .io_in_0_ready(inputArb_io_in_0_ready),
    .io_in_0_valid(inputArb_io_in_0_valid),
    .io_in_0_bits_addr(inputArb_io_in_0_bits_addr),
    .io_in_0_bits_size(inputArb_io_in_0_bits_size),
    .io_in_0_bits_cmd(inputArb_io_in_0_bits_cmd),
    .io_in_0_bits_wmask(inputArb_io_in_0_bits_wmask),
    .io_in_0_bits_wdata(inputArb_io_in_0_bits_wdata),
    .io_in_1_ready(inputArb_io_in_1_ready),
    .io_in_1_valid(inputArb_io_in_1_valid),
    .io_in_1_bits_addr(inputArb_io_in_1_bits_addr),
    .io_in_1_bits_cmd(inputArb_io_in_1_bits_cmd),
    .io_in_1_bits_wdata(inputArb_io_in_1_bits_wdata),
    .io_in_2_ready(inputArb_io_in_2_ready),
    .io_in_2_valid(inputArb_io_in_2_valid),
    .io_in_2_bits_addr(inputArb_io_in_2_bits_addr),
    .io_in_2_bits_cmd(inputArb_io_in_2_bits_cmd),
    .io_in_2_bits_wdata(inputArb_io_in_2_bits_wdata),
    .io_in_3_ready(inputArb_io_in_3_ready),
    .io_in_3_valid(inputArb_io_in_3_valid),
    .io_in_3_bits_addr(inputArb_io_in_3_bits_addr),
    .io_in_3_bits_size(inputArb_io_in_3_bits_size),
    .io_in_3_bits_cmd(inputArb_io_in_3_bits_cmd),
    .io_in_3_bits_wmask(inputArb_io_in_3_bits_wmask),
    .io_in_3_bits_wdata(inputArb_io_in_3_bits_wdata),
    .io_out_ready(inputArb_io_out_ready),
    .io_out_valid(inputArb_io_out_valid),
    .io_out_bits_addr(inputArb_io_out_bits_addr),
    .io_out_bits_size(inputArb_io_out_bits_size),
    .io_out_bits_cmd(inputArb_io_out_bits_cmd),
    .io_out_bits_wmask(inputArb_io_out_bits_wmask),
    .io_out_bits_wdata(inputArb_io_out_bits_wdata),
    .io_chosen(inputArb_io_chosen)
  );
  assign io_in_0_req_ready = inputArb_io_in_0_ready; // @[src/main/scala/bus/simplebus/Crossbar.scala 96:68]
  assign io_in_0_resp_valid = 2'h0 == inflightSrc & io_out_resp_valid; // @[src/main/scala/bus/simplebus/Crossbar.scala 109:{13,13} 107:26]
  assign io_in_0_resp_bits_cmd = io_out_resp_bits_cmd; // @[src/main/scala/bus/simplebus/Crossbar.scala 106:25]
  assign io_in_0_resp_bits_rdata = io_out_resp_bits_rdata; // @[src/main/scala/bus/simplebus/Crossbar.scala 106:25]
  assign io_in_1_req_ready = inputArb_io_in_1_ready; // @[src/main/scala/bus/simplebus/Crossbar.scala 96:68]
  assign io_in_1_resp_valid = 2'h1 == inflightSrc & io_out_resp_valid; // @[src/main/scala/bus/simplebus/Crossbar.scala 109:{13,13} 107:26]
  assign io_in_1_resp_bits_cmd = io_out_resp_bits_cmd; // @[src/main/scala/bus/simplebus/Crossbar.scala 106:25]
  assign io_in_1_resp_bits_rdata = io_out_resp_bits_rdata; // @[src/main/scala/bus/simplebus/Crossbar.scala 106:25]
  assign io_in_2_req_ready = inputArb_io_in_2_ready; // @[src/main/scala/bus/simplebus/Crossbar.scala 96:68]
  assign io_in_2_resp_valid = 2'h2 == inflightSrc & io_out_resp_valid; // @[src/main/scala/bus/simplebus/Crossbar.scala 109:{13,13} 107:26]
  assign io_in_2_resp_bits_cmd = io_out_resp_bits_cmd; // @[src/main/scala/bus/simplebus/Crossbar.scala 106:25]
  assign io_in_2_resp_bits_rdata = io_out_resp_bits_rdata; // @[src/main/scala/bus/simplebus/Crossbar.scala 106:25]
  assign io_in_3_req_ready = inputArb_io_in_3_ready; // @[src/main/scala/bus/simplebus/Crossbar.scala 96:68]
  assign io_in_3_resp_valid = 2'h3 == inflightSrc & io_out_resp_valid; // @[src/main/scala/bus/simplebus/Crossbar.scala 109:{13,13} 107:26]
  assign io_in_3_resp_bits_cmd = io_out_resp_bits_cmd; // @[src/main/scala/bus/simplebus/Crossbar.scala 106:25]
  assign io_in_3_resp_bits_rdata = io_out_resp_bits_rdata; // @[src/main/scala/bus/simplebus/Crossbar.scala 106:25]
  assign io_out_req_valid = inputArb_io_out_valid & state == 2'h0; // @[src/main/scala/bus/simplebus/Crossbar.scala 103:37]
  assign io_out_req_bits_addr = inputArb_io_out_bits_addr; // @[src/main/scala/bus/simplebus/Crossbar.scala 101:19]
  assign io_out_req_bits_size = inputArb_io_out_bits_size; // @[src/main/scala/bus/simplebus/Crossbar.scala 101:19]
  assign io_out_req_bits_cmd = inputArb_io_out_bits_cmd; // @[src/main/scala/bus/simplebus/Crossbar.scala 101:19]
  assign io_out_req_bits_wmask = inputArb_io_out_bits_wmask; // @[src/main/scala/bus/simplebus/Crossbar.scala 101:19]
  assign io_out_req_bits_wdata = inputArb_io_out_bits_wdata; // @[src/main/scala/bus/simplebus/Crossbar.scala 101:19]
  assign io_out_resp_ready = 2'h3 == inflightSrc ? io_in_3_resp_ready : 1'h1; // @[src/main/scala/bus/simplebus/Crossbar.scala 110:{13,13}]
  assign inputArb_clock = clock;
  assign inputArb_reset = reset;
  assign inputArb_io_in_0_valid = io_in_0_req_valid; // @[src/main/scala/bus/simplebus/Crossbar.scala 96:68]
  assign inputArb_io_in_0_bits_addr = io_in_0_req_bits_addr; // @[src/main/scala/bus/simplebus/Crossbar.scala 96:68]
  assign inputArb_io_in_0_bits_size = io_in_0_req_bits_size; // @[src/main/scala/bus/simplebus/Crossbar.scala 96:68]
  assign inputArb_io_in_0_bits_cmd = io_in_0_req_bits_cmd; // @[src/main/scala/bus/simplebus/Crossbar.scala 96:68]
  assign inputArb_io_in_0_bits_wmask = io_in_0_req_bits_wmask; // @[src/main/scala/bus/simplebus/Crossbar.scala 96:68]
  assign inputArb_io_in_0_bits_wdata = io_in_0_req_bits_wdata; // @[src/main/scala/bus/simplebus/Crossbar.scala 96:68]
  assign inputArb_io_in_1_valid = io_in_1_req_valid; // @[src/main/scala/bus/simplebus/Crossbar.scala 96:68]
  assign inputArb_io_in_1_bits_addr = io_in_1_req_bits_addr; // @[src/main/scala/bus/simplebus/Crossbar.scala 96:68]
  assign inputArb_io_in_1_bits_cmd = io_in_1_req_bits_cmd; // @[src/main/scala/bus/simplebus/Crossbar.scala 96:68]
  assign inputArb_io_in_1_bits_wdata = io_in_1_req_bits_wdata; // @[src/main/scala/bus/simplebus/Crossbar.scala 96:68]
  assign inputArb_io_in_2_valid = io_in_2_req_valid; // @[src/main/scala/bus/simplebus/Crossbar.scala 96:68]
  assign inputArb_io_in_2_bits_addr = io_in_2_req_bits_addr; // @[src/main/scala/bus/simplebus/Crossbar.scala 96:68]
  assign inputArb_io_in_2_bits_cmd = io_in_2_req_bits_cmd; // @[src/main/scala/bus/simplebus/Crossbar.scala 96:68]
  assign inputArb_io_in_2_bits_wdata = io_in_2_req_bits_wdata; // @[src/main/scala/bus/simplebus/Crossbar.scala 96:68]
  assign inputArb_io_in_3_valid = io_in_3_req_valid; // @[src/main/scala/bus/simplebus/Crossbar.scala 96:68]
  assign inputArb_io_in_3_bits_addr = io_in_3_req_bits_addr; // @[src/main/scala/bus/simplebus/Crossbar.scala 96:68]
  assign inputArb_io_in_3_bits_size = io_in_3_req_bits_size; // @[src/main/scala/bus/simplebus/Crossbar.scala 96:68]
  assign inputArb_io_in_3_bits_cmd = io_in_3_req_bits_cmd; // @[src/main/scala/bus/simplebus/Crossbar.scala 96:68]
  assign inputArb_io_in_3_bits_wmask = io_in_3_req_bits_wmask; // @[src/main/scala/bus/simplebus/Crossbar.scala 96:68]
  assign inputArb_io_in_3_bits_wdata = io_in_3_req_bits_wdata; // @[src/main/scala/bus/simplebus/Crossbar.scala 96:68]
  assign inputArb_io_out_ready = io_out_req_ready & _io_out_req_valid_T; // @[src/main/scala/bus/simplebus/Crossbar.scala 104:37]
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 92:22]
      state <= 2'h0; // @[src/main/scala/bus/simplebus/Crossbar.scala 92:22]
    end else if (2'h0 == state) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 113:18]
      if (_T_15) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 115:27]
        if (_T_4) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 117:38]
          state <= 2'h1; // @[src/main/scala/bus/simplebus/Crossbar.scala 117:46]
        end else begin
          state <= _GEN_8;
        end
      end
    end else if (2'h1 == state) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 113:18]
      if (_T_25 & _T_26) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 121:78]
        state <= 2'h0; // @[src/main/scala/bus/simplebus/Crossbar.scala 121:86]
      end
    end else if (2'h2 == state) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 113:18]
      state <= _GEN_13;
    end
    if (reset) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 99:28]
      inflightSrc <= 2'h0; // @[src/main/scala/bus/simplebus/Crossbar.scala 99:28]
    end else if (2'h0 == state) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 113:18]
      if (_T_15) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 115:27]
        inflightSrc <= inputArb_io_chosen; // @[src/main/scala/bus/simplebus/Crossbar.scala 116:21]
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~(inputArb_io_out_valid & ~_T_4 & _T_1))) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Crossbar.scala:98 assert(!(thisReq.valid && !thisReq.bits.isRead() && !thisReq.bits.isWrite()))\n"
            ); // @[src/main/scala/bus/simplebus/Crossbar.scala 98:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~(inputArb_io_out_valid & ~_T_4 & _T_1)) & ~reset) begin
          $fatal; // @[src/main/scala/bus/simplebus/Crossbar.scala 98:9]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  inflightSrc = _RAND_1[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module EmbeddedTLBExec(
  input          clock,
  input          reset,
  output         io_in_ready, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 178:14]
  input          io_in_valid, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 178:14]
  input  [38:0]  io_in_bits_addr, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 178:14]
  input  [86:0]  io_in_bits_user, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 178:14]
  input          io_out_ready, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 178:14]
  output         io_out_valid, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 178:14]
  output [31:0]  io_out_bits_addr, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 178:14]
  output [86:0]  io_out_bits_user, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 178:14]
  input  [120:0] io_md_0, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 178:14]
  input  [120:0] io_md_1, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 178:14]
  input  [120:0] io_md_2, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 178:14]
  input  [120:0] io_md_3, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 178:14]
  output         io_mdWrite_wen, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 178:14]
  output         io_mdWrite_windex, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 178:14]
  output [3:0]   io_mdWrite_waymask, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 178:14]
  output [120:0] io_mdWrite_wdata, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 178:14]
  input          io_mdReady, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 178:14]
  input          io_mem_req_ready, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 178:14]
  output         io_mem_req_valid, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 178:14]
  output [31:0]  io_mem_req_bits_addr, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 178:14]
  output [2:0]   io_mem_req_bits_size, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 178:14]
  output [3:0]   io_mem_req_bits_cmd, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 178:14]
  output [7:0]   io_mem_req_bits_wmask, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 178:14]
  output [63:0]  io_mem_req_bits_wdata, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 178:14]
  output         io_mem_resp_ready, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 178:14]
  input          io_mem_resp_valid, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 178:14]
  input  [3:0]   io_mem_resp_bits_cmd, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 178:14]
  input  [63:0]  io_mem_resp_bits_rdata, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 178:14]
  input          io_flush, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 178:14]
  input  [63:0]  io_satp, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 178:14]
  input  [1:0]   io_pf_priviledgeMode, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 178:14]
  output         io_pf_loadPF, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 178:14]
  output         io_pf_storePF, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 178:14]
  output         io_ipf, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 178:14]
  output         io_isFinish, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 178:14]
  input          DISPLAY_ENABLE
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [63:0] _RAND_20;
  reg [63:0] _RAND_21;
  reg [63:0] _RAND_22;
  reg [63:0] _RAND_23;
  reg [63:0] _RAND_24;
  reg [63:0] _RAND_25;
  reg [63:0] _RAND_26;
  reg [63:0] _RAND_27;
`endif // RANDOMIZE_REG_INIT
  wire [8:0] vpn_vpn0 = io_in_bits_addr[20:12]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 198:54]
  wire [8:0] vpn_vpn1 = io_in_bits_addr[29:21]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 198:54]
  wire [8:0] vpn_vpn2 = io_in_bits_addr[38:30]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 198:54]
  wire [19:0] satp_ppn = io_satp[19:0]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 200:30]
  wire [15:0] satp_asid = io_satp[59:44]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 200:30]
  wire [17:0] hitVec_hi = {vpn_vpn2,vpn_vpn1}; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 209:201]
  wire [26:0] _hitVec_T_34 = {vpn_vpn2,vpn_vpn1,vpn_vpn0}; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 209:201]
  wire [26:0] _hitVec_T_35 = {9'h1ff,io_md_0[77:60]}; // @[src/main/scala/nutcore/mem/TLB.scala 131:9]
  wire [26:0] _hitVec_T_36 = _hitVec_T_35 & io_md_0[120:94]; // @[src/main/scala/nutcore/mem/TLB.scala 131:37]
  wire [26:0] _hitVec_T_38 = _hitVec_T_35 & _hitVec_T_34; // @[src/main/scala/nutcore/mem/TLB.scala 131:84]
  wire  _hitVec_T_39 = _hitVec_T_36 == _hitVec_T_38; // @[src/main/scala/nutcore/mem/TLB.scala 131:48]
  wire  _hitVec_T_40 = io_md_0[52] & io_md_0[93:78] == satp_asid & _hitVec_T_39; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 209:132]
  wire [26:0] _hitVec_T_76 = {9'h1ff,io_md_1[77:60]}; // @[src/main/scala/nutcore/mem/TLB.scala 131:9]
  wire [26:0] _hitVec_T_77 = _hitVec_T_76 & io_md_1[120:94]; // @[src/main/scala/nutcore/mem/TLB.scala 131:37]
  wire [26:0] _hitVec_T_79 = _hitVec_T_76 & _hitVec_T_34; // @[src/main/scala/nutcore/mem/TLB.scala 131:84]
  wire  _hitVec_T_80 = _hitVec_T_77 == _hitVec_T_79; // @[src/main/scala/nutcore/mem/TLB.scala 131:48]
  wire  _hitVec_T_81 = io_md_1[52] & io_md_1[93:78] == satp_asid & _hitVec_T_80; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 209:132]
  wire [26:0] _hitVec_T_117 = {9'h1ff,io_md_2[77:60]}; // @[src/main/scala/nutcore/mem/TLB.scala 131:9]
  wire [26:0] _hitVec_T_118 = _hitVec_T_117 & io_md_2[120:94]; // @[src/main/scala/nutcore/mem/TLB.scala 131:37]
  wire [26:0] _hitVec_T_120 = _hitVec_T_117 & _hitVec_T_34; // @[src/main/scala/nutcore/mem/TLB.scala 131:84]
  wire  _hitVec_T_121 = _hitVec_T_118 == _hitVec_T_120; // @[src/main/scala/nutcore/mem/TLB.scala 131:48]
  wire  _hitVec_T_122 = io_md_2[52] & io_md_2[93:78] == satp_asid & _hitVec_T_121; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 209:132]
  wire [26:0] _hitVec_T_158 = {9'h1ff,io_md_3[77:60]}; // @[src/main/scala/nutcore/mem/TLB.scala 131:9]
  wire [26:0] _hitVec_T_159 = _hitVec_T_158 & io_md_3[120:94]; // @[src/main/scala/nutcore/mem/TLB.scala 131:37]
  wire [26:0] _hitVec_T_161 = _hitVec_T_158 & _hitVec_T_34; // @[src/main/scala/nutcore/mem/TLB.scala 131:84]
  wire  _hitVec_T_162 = _hitVec_T_159 == _hitVec_T_161; // @[src/main/scala/nutcore/mem/TLB.scala 131:48]
  wire  _hitVec_T_163 = io_md_3[52] & io_md_3[93:78] == satp_asid & _hitVec_T_162; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 209:132]
  wire [3:0] hitVec = {_hitVec_T_163,_hitVec_T_122,_hitVec_T_81,_hitVec_T_40}; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 209:211]
  wire  _hit_T = |hitVec; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 210:35]
  wire  hit = io_in_valid & |hitVec; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 210:25]
  wire  miss = io_in_valid & ~_hit_T; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 211:26]
  reg [63:0] victimWaymask_lfsr; // @[src/main/scala/utils/LFSR64.scala 25:23]
  wire  victimWaymask_xor = victimWaymask_lfsr[0] ^ victimWaymask_lfsr[1] ^ victimWaymask_lfsr[3] ^ victimWaymask_lfsr[4
    ]; // @[src/main/scala/utils/LFSR64.scala 26:43]
  wire [63:0] _victimWaymask_lfsr_T_2 = {victimWaymask_xor,victimWaymask_lfsr[63:1]}; // @[src/main/scala/utils/LFSR64.scala 28:41]
  wire [3:0] victimWaymask = 4'h1 << victimWaymask_lfsr[1:0]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 213:42]
  wire [3:0] waymask = hit ? hitVec : victimWaymask; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 214:20]
  wire [120:0] _hitMeta_T_4 = waymask[0] ? io_md_0 : 121'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [120:0] _hitMeta_T_5 = waymask[1] ? io_md_1 : 121'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [120:0] _hitMeta_T_6 = waymask[2] ? io_md_2 : 121'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [120:0] _hitMeta_T_7 = waymask[3] ? io_md_3 : 121'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [120:0] _hitMeta_T_8 = _hitMeta_T_4 | _hitMeta_T_5; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [120:0] _hitMeta_T_9 = _hitMeta_T_8 | _hitMeta_T_6; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [120:0] _hitMeta_T_10 = _hitMeta_T_9 | _hitMeta_T_7; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [7:0] hitMeta_flag = _hitMeta_T_10[59:52]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 220:70]
  wire [17:0] hitMeta_mask = _hitMeta_T_10[77:60]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 220:70]
  wire [15:0] hitMeta_asid = _hitMeta_T_10[93:78]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 220:70]
  wire [26:0] hitMeta_vpn = _hitMeta_T_10[120:94]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 220:70]
  wire [31:0] hitData_pteaddr = _hitMeta_T_10[31:0]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:70]
  wire [19:0] hitData_ppn = _hitMeta_T_10[51:32]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:70]
  wire  hitFlag_v = hitMeta_flag[0]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 222:38]
  wire  hitFlag_r = hitMeta_flag[1]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 222:38]
  wire  hitFlag_w = hitMeta_flag[2]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 222:38]
  wire  hitFlag_x = hitMeta_flag[3]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 222:38]
  wire  hitFlag_u = hitMeta_flag[4]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 222:38]
  wire  hitFlag_g = hitMeta_flag[5]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 222:38]
  wire  hitFlag_a = hitMeta_flag[6]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 222:38]
  wire  hitFlag_d = hitMeta_flag[7]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 222:38]
  wire  _hitWB_T = ~hitFlag_a; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 226:23]
  wire  _hitCheck_T = io_pf_priviledgeMode == 2'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 231:62]
  wire  _hitCheck_T_5 = io_pf_priviledgeMode == 2'h1; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 231:110]
  wire  hitCheck = hit & ~(io_pf_priviledgeMode == 2'h0 & ~hitFlag_u) & ~(io_pf_priviledgeMode == 2'h1 & hitFlag_u); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 231:87]
  wire  _hitExec_T_1 = hitCheck & ~_hitWB_T; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 233:26]
  wire  hitExec = hitCheck & ~_hitWB_T & hitFlag_x; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 233:41]
  wire  hitinstrPF = ~hitExec & hit; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 245:52]
  wire  _hitWB_T_9 = io_pf_loadPF | io_pf_storePF; // @[src/main/scala/nutcore/Bundle.scala 131:23]
  wire  _hitWB_T_11 = ~_hitWB_T_9; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 226:84]
  wire  hitWB = hit & ~hitFlag_a & ~hitinstrPF & ~_hitWB_T_9; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 226:81]
  wire [7:0] _hitRefillFlag_T_2 = {hitFlag_d,hitFlag_a,hitFlag_g,hitFlag_u,hitFlag_x,hitFlag_w,hitFlag_r,hitFlag_v}; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 227:79]
  wire [7:0] hitRefillFlag = 8'h40 | _hitRefillFlag_T_2; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 227:69]
  wire [39:0] _hitWBStore_T = {10'h0,hitData_ppn,2'h0,hitRefillFlag}; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 228:33]
  reg [39:0] hitWBStore; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 228:29]
  wire  hitLoad = _hitExec_T_1 & hitFlag_r; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 234:41]
  wire  hitStore = _hitExec_T_1 & hitFlag_w; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 235:42]
  reg [2:0] state; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 253:22]
  reg [1:0] level; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 254:22]
  reg [63:0] memRespStore; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 256:25]
  reg [17:0] missMaskStore; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 258:26]
  wire  memRdata_flag_v = io_mem_resp_bits_rdata[0]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 261:49]
  wire  memRdata_flag_r = io_mem_resp_bits_rdata[1]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 261:49]
  wire  memRdata_flag_w = io_mem_resp_bits_rdata[2]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 261:49]
  wire  memRdata_flag_x = io_mem_resp_bits_rdata[3]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 261:49]
  wire  memRdata_flag_u = io_mem_resp_bits_rdata[4]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 261:49]
  wire  memRdata_flag_g = io_mem_resp_bits_rdata[5]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 261:49]
  wire  memRdata_flag_a = io_mem_resp_bits_rdata[6]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 261:49]
  wire  memRdata_flag_d = io_mem_resp_bits_rdata[7]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 261:49]
  wire [1:0] memRdata_rsw = io_mem_resp_bits_rdata[9:8]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 261:49]
  wire [19:0] memRdata_ppn = io_mem_resp_bits_rdata[29:10]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 261:49]
  wire [33:0] memRdata_reserved = io_mem_resp_bits_rdata[63:30]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 261:49]
  reg [31:0] raddr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 262:18]
  wire  _alreadyOutFire_T = io_out_ready & io_out_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  reg  alreadyOutFire; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 263:33]
  wire  _GEN_2 = _alreadyOutFire_T | alreadyOutFire; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 263:{33,33,33}]
  reg  needFlush; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 266:26]
  wire  isFlush = needFlush | io_flush; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 268:27]
  wire  _GEN_3 = io_flush & state != 3'h0 | needFlush; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 266:26 269:{40,52}]
  wire  _GEN_4 = _alreadyOutFire_T & needFlush ? 1'h0 : _GEN_3; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 270:{35,47}]
  reg  missIPF; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 272:24]
  wire  _T_4 = 3'h0 == state; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 275:18]
  wire  _T_5 = ~io_flush; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 277:13]
  wire [31:0] _raddr_T_1 = {satp_ppn,vpn_vpn2,3'h0}; // @[src/main/scala/nutcore/mem/TLB.scala 89:8]
  wire  _T_9 = 3'h1 == state; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 275:18]
  wire  _T_10 = io_mem_req_ready & io_mem_req_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  wire [2:0] _GEN_15 = _T_10 ? 3'h2 : state; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 253:22 294:{36,44}]
  wire  _GEN_17 = isFlush ? 1'h0 : _GEN_4; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 291:22 293:19]
  wire  _T_11 = 3'h2 == state; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 275:18]
  wire [7:0] _missflag_T = {memRdata_flag_d,memRdata_flag_a,memRdata_flag_g,memRdata_flag_u,memRdata_flag_x,
    memRdata_flag_w,memRdata_flag_r,memRdata_flag_v}; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 298:44]
  wire  missflag_v = _missflag_T[0]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 298:44]
  wire  missflag_r = _missflag_T[1]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 298:44]
  wire  missflag_w = _missflag_T[2]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 298:44]
  wire  missflag_x = _missflag_T[3]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 298:44]
  wire  missflag_u = _missflag_T[4]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 298:44]
  wire  missflag_g = _missflag_T[5]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 298:44]
  wire  missflag_a = _missflag_T[6]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 298:44]
  wire  missflag_d = _missflag_T[7]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 298:44]
  wire  _T_12 = io_mem_resp_ready & io_mem_resp_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  wire  _T_15 = level == 2'h3; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 303:58]
  wire  _T_16 = level == 2'h2; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 303:73]
  wire  _T_18 = ~(missflag_r | missflag_x) & (level == 2'h3 | level == 2'h2); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 303:49]
  wire  _T_22 = ~missflag_v | ~missflag_r & missflag_w; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 304:28]
  reg [63:0] c; // @[src/main/scala/utils/GTimer.scala 24:20]
  wire [63:0] _c_T_1 = c + 64'h1; // @[src/main/scala/utils/GTimer.scala 25:12]
  wire  _T_25 = ~reset; // @[src/main/scala/utils/Debug.scala 56:24]
  wire [8:0] _raddr_T_3 = _T_15 ? vpn_vpn1 : vpn_vpn0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 317:50]
  wire [31:0] _raddr_T_5 = {memRdata_ppn,_raddr_T_3,3'h0}; // @[src/main/scala/nutcore/mem/TLB.scala 89:8]
  wire [2:0] _GEN_18 = ~missflag_v | ~missflag_r & missflag_w ? 3'h4 : 3'h1; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 304:60 305:43 316:19]
  wire  _GEN_19 = ~missflag_v | ~missflag_r & missflag_w | missIPF; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 272:24 304:60 306:45]
  wire [31:0] _GEN_20 = ~missflag_v | ~missflag_r & missflag_w ? raddr : _raddr_T_5; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 262:18 304:60 317:19]
  wire  permCheck = missflag_v & ~(_hitCheck_T & ~missflag_u) & ~(_hitCheck_T_5 & missflag_u); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 320:87]
  wire  permAD = ~missflag_a; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 321:71]
  wire  permExec = permCheck & ~permAD & missflag_x; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:47]
  wire [7:0] _missRefillFlag_T_2 = {missflag_d,missflag_a,missflag_g,missflag_u,missflag_x,missflag_w,missflag_r,
    missflag_v}; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 327:79]
  wire [7:0] _missRefillFlag_T_3 = 8'h40 | _missRefillFlag_T_2; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 327:68]
  wire [63:0] _memRespStore_T = io_mem_resp_bits_rdata | 64'h40; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 328:50]
  wire  _GEN_21 = ~permExec | missIPF; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 272:24 330:{30,40}]
  wire  _GEN_23 = ~permExec ? 1'h0 : 1'h1; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 330:30 259:32 333:30]
  wire [17:0] _missMask_T_2 = _T_16 ? 18'h3fe00 : 18'h3ffff; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 346:59]
  wire [17:0] _missMask_T_3 = _T_15 ? 18'h0 : _missMask_T_2; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 346:26]
  wire [7:0] _GEN_24 = level != 2'h0 ? _missRefillFlag_T_3 : 8'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 319:36 327:26 260:32]
  wire [63:0] _GEN_25 = level != 2'h0 ? _memRespStore_T : memRespStore; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 319:36 328:24 256:25]
  wire  _GEN_26 = level != 2'h0 ? _GEN_21 : missIPF; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 272:24 319:36]
  wire [2:0] _GEN_27 = level != 2'h0 ? 3'h4 : state; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 253:22 319:36]
  wire  _GEN_28 = level != 2'h0 & _GEN_23; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 259:32 319:36]
  wire [17:0] _GEN_29 = level != 2'h0 ? _missMask_T_3 : 18'h3ffff; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 319:36 346:20 257:26]
  wire [17:0] _GEN_37 = ~(missflag_r | missflag_x) & (level == 2'h3 | level == 2'h2) ? 18'h3ffff : _GEN_29; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 257:26 303:82]
  wire [17:0] _GEN_45 = isFlush ? 18'h3ffff : _GEN_37; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 300:24 257:26]
  wire [17:0] _GEN_54 = _T_12 ? _GEN_45 : 18'h3ffff; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 257:26 299:31]
  wire [17:0] _GEN_77 = 3'h2 == state ? _GEN_54 : 18'h3ffff; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 275:18 257:26]
  wire [17:0] _GEN_88 = 3'h1 == state ? 18'h3ffff : _GEN_77; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 275:18 257:26]
  wire [17:0] missMask = 3'h0 == state ? 18'h3ffff : _GEN_88; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 275:18 257:26]
  wire [17:0] _GEN_30 = level != 2'h0 ? missMask : missMaskStore; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 319:36 347:25 258:26]
  wire [2:0] _GEN_31 = ~(missflag_r | missflag_x) & (level == 2'h3 | level == 2'h2) ? _GEN_18 : _GEN_27; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 303:82]
  wire  _GEN_32 = ~(missflag_r | missflag_x) & (level == 2'h3 | level == 2'h2) ? _GEN_19 : _GEN_26; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 303:82]
  wire [31:0] _GEN_33 = ~(missflag_r | missflag_x) & (level == 2'h3 | level == 2'h2) ? _GEN_20 : raddr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 262:18 303:82]
  wire [7:0] _GEN_34 = ~(missflag_r | missflag_x) & (level == 2'h3 | level == 2'h2) ? 8'h0 : _GEN_24; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 260:32 303:82]
  wire [63:0] _GEN_35 = ~(missflag_r | missflag_x) & (level == 2'h3 | level == 2'h2) ? memRespStore : _GEN_25; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 256:25 303:82]
  wire  _GEN_36 = ~(missflag_r | missflag_x) & (level == 2'h3 | level == 2'h2) ? 1'h0 : _GEN_28; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 259:32 303:82]
  wire [17:0] _GEN_38 = ~(missflag_r | missflag_x) & (level == 2'h3 | level == 2'h2) ? missMaskStore : _GEN_30; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 258:26 303:82]
  wire [2:0] _GEN_39 = isFlush ? 3'h0 : _GEN_31; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 300:24 301:17]
  wire  _GEN_40 = isFlush ? missIPF : _GEN_32; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 272:24 300:24]
  wire [31:0] _GEN_41 = isFlush ? raddr : _GEN_33; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 262:18 300:24]
  wire [7:0] _GEN_42 = isFlush ? 8'h0 : _GEN_34; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 300:24 260:32]
  wire [63:0] _GEN_43 = isFlush ? memRespStore : _GEN_35; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 300:24 256:25]
  wire  _GEN_44 = isFlush ? 1'h0 : _GEN_36; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 300:24 259:32]
  wire [17:0] _GEN_46 = isFlush ? missMaskStore : _GEN_38; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 300:24 258:26]
  wire [1:0] _level_T_1 = level - 2'h1; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 349:24]
  wire [2:0] _GEN_47 = _T_12 ? _GEN_39 : state; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 253:22 299:31]
  wire  _GEN_48 = _T_12 ? _GEN_17 : _GEN_4; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 299:31]
  wire  _GEN_49 = _T_12 ? _GEN_40 : missIPF; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 272:24 299:31]
  wire [7:0] _GEN_51 = _T_12 ? _GEN_42 : 8'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 299:31 260:32]
  wire  _GEN_53 = _T_12 & _GEN_44; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 299:31 259:32]
  wire [1:0] _GEN_56 = _T_12 ? _level_T_1 : level; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 299:31 349:15 254:22]
  wire [2:0] _GEN_57 = _T_10 ? 3'h4 : state; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 253:22 357:{36,44}]
  wire [2:0] _GEN_58 = isFlush ? 3'h0 : _GEN_57; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 354:22 355:15]
  wire [2:0] _GEN_59 = _alreadyOutFire_T | io_flush | alreadyOutFire ? 3'h0 : state; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 360:71 361:13 253:22]
  wire  _GEN_60 = _alreadyOutFire_T | io_flush | alreadyOutFire ? 1'h0 : missIPF; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 360:71 362:15 272:24]
  wire  _GEN_61 = _alreadyOutFire_T | io_flush | alreadyOutFire ? 1'h0 : _GEN_2; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 360:71 363:22]
  wire [2:0] _GEN_62 = 3'h5 == state ? 3'h0 : state; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 275:18 367:13 253:22]
  wire [2:0] _GEN_63 = 3'h4 == state ? _GEN_59 : _GEN_62; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 275:18]
  wire  _GEN_64 = 3'h4 == state ? _GEN_60 : missIPF; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 275:18 272:24]
  wire  _GEN_65 = 3'h4 == state ? _GEN_61 : _GEN_2; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 275:18]
  wire [2:0] _GEN_66 = 3'h3 == state ? _GEN_58 : _GEN_63; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 275:18]
  wire  _GEN_67 = 3'h3 == state ? _GEN_17 : _GEN_4; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 275:18]
  wire  _GEN_68 = 3'h3 == state ? missIPF : _GEN_64; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 275:18 272:24]
  wire  _GEN_69 = 3'h3 == state ? _GEN_2 : _GEN_65; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 275:18]
  wire [7:0] _GEN_74 = 3'h2 == state ? _GEN_51 : 8'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 275:18 260:32]
  wire [7:0] _GEN_85 = 3'h1 == state ? 8'h0 : _GEN_74; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 275:18 260:32]
  wire  _GEN_87 = 3'h1 == state ? 1'h0 : 3'h2 == state & _GEN_53; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 275:18 259:32]
  wire [7:0] missRefillFlag = 3'h0 == state ? 8'h0 : _GEN_85; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 275:18 260:32]
  wire  missMetaRefill = 3'h0 == state ? 1'h0 : _GEN_87; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 275:18 259:32]
  wire  cmd = state == 3'h3; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 372:23]
  wire  _io_mem_req_valid_T_3 = ~isFlush; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 374:77]
  wire  _T_50 = state == 3'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 378:82]
  reg  REG; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 378:33]
  reg  REG_1; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 379:21]
  reg [3:0] REG_2; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 379:60]
  reg [26:0] REG_3; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 379:84]
  reg [15:0] REG_4; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 380:19]
  reg [17:0] REG_5; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 380:72]
  reg [7:0] REG_6; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 381:19]
  reg [19:0] REG_7; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 381:77]
  reg [31:0] REG_8; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 382:22]
  wire [59:0] io_mdWrite_wdata_lo = {REG_6,REG_7,REG_8}; // @[src/main/scala/nutcore/mem/TLB.scala 217:22]
  wire [60:0] io_mdWrite_wdata_hi = {REG_3,REG_4,REG_5}; // @[src/main/scala/nutcore/mem/TLB.scala 217:22]
  wire [31:0] _io_out_bits_addr_T_1 = {hitData_ppn,12'h0}; // @[src/main/scala/nutcore/mem/TLB.scala 127:24]
  wire [31:0] _io_out_bits_addr_T_3 = {2'h3,hitMeta_mask,12'h0}; // @[src/main/scala/nutcore/mem/TLB.scala 127:49]
  wire [31:0] _io_out_bits_addr_T_4 = _io_out_bits_addr_T_1 & _io_out_bits_addr_T_3; // @[src/main/scala/utils/BitUtils.scala 34:14]
  wire [31:0] _io_out_bits_addr_T_5 = ~_io_out_bits_addr_T_3; // @[src/main/scala/utils/BitUtils.scala 34:39]
  wire [31:0] _io_out_bits_addr_T_6 = io_in_bits_addr[31:0] & _io_out_bits_addr_T_5; // @[src/main/scala/utils/BitUtils.scala 34:37]
  wire [31:0] _io_out_bits_addr_T_7 = _io_out_bits_addr_T_4 | _io_out_bits_addr_T_6; // @[src/main/scala/utils/BitUtils.scala 34:26]
  wire [31:0] _io_out_bits_addr_T_20 = {memRespStore[29:10],12'h0}; // @[src/main/scala/nutcore/mem/TLB.scala 127:24]
  wire [31:0] _io_out_bits_addr_T_22 = {2'h3,missMaskStore,12'h0}; // @[src/main/scala/nutcore/mem/TLB.scala 127:49]
  wire [31:0] _io_out_bits_addr_T_23 = _io_out_bits_addr_T_20 & _io_out_bits_addr_T_22; // @[src/main/scala/utils/BitUtils.scala 34:14]
  wire [31:0] _io_out_bits_addr_T_24 = ~_io_out_bits_addr_T_22; // @[src/main/scala/utils/BitUtils.scala 34:39]
  wire [31:0] _io_out_bits_addr_T_25 = io_in_bits_addr[31:0] & _io_out_bits_addr_T_24; // @[src/main/scala/utils/BitUtils.scala 34:37]
  wire [31:0] _io_out_bits_addr_T_26 = _io_out_bits_addr_T_23 | _io_out_bits_addr_T_25; // @[src/main/scala/utils/BitUtils.scala 34:26]
  wire  _io_out_valid_T = ~hitWB; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 387:45]
  wire  _io_out_valid_T_7 = hit & ~hitWB ? _hitWB_T_11 : state == 3'h4; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 387:37]
  reg [63:0] c_4; // @[src/main/scala/utils/GTimer.scala 24:20]
  wire [63:0] _c_T_9 = c_4 + 64'h1; // @[src/main/scala/utils/GTimer.scala 25:12]
  reg [63:0] c_5; // @[src/main/scala/utils/GTimer.scala 24:20]
  wire [63:0] _c_T_11 = c_5 + 64'h1; // @[src/main/scala/utils/GTimer.scala 25:12]
  reg [63:0] c_6; // @[src/main/scala/utils/GTimer.scala 24:20]
  wire [63:0] _c_T_13 = c_6 + 64'h1; // @[src/main/scala/utils/GTimer.scala 25:12]
  wire [4:0] lo_1 = {memRdata_flag_u,memRdata_flag_x,memRdata_flag_w,memRdata_flag_r,memRdata_flag_v}; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 397:145]
  wire [63:0] _T_80 = {memRdata_reserved,memRdata_ppn,memRdata_rsw,memRdata_flag_d,memRdata_flag_a,memRdata_flag_g,lo_1}
    ; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 397:145]
  reg [63:0] c_7; // @[src/main/scala/utils/GTimer.scala 24:20]
  wire [63:0] _c_T_15 = c_7 + 64'h1; // @[src/main/scala/utils/GTimer.scala 25:12]
  reg [63:0] c_8; // @[src/main/scala/utils/GTimer.scala 24:20]
  wire [63:0] _c_T_17 = c_8 + 64'h1; // @[src/main/scala/utils/GTimer.scala 25:12]
  reg [63:0] c_9; // @[src/main/scala/utils/GTimer.scala 24:20]
  wire [63:0] _c_T_19 = c_9 + 64'h1; // @[src/main/scala/utils/GTimer.scala 25:12]
  reg [63:0] c_10; // @[src/main/scala/utils/GTimer.scala 24:20]
  wire [63:0] _c_T_21 = c_10 + 64'h1; // @[src/main/scala/utils/GTimer.scala 25:12]
  reg [63:0] c_11; // @[src/main/scala/utils/GTimer.scala 24:20]
  wire [63:0] _c_T_23 = c_11 + 64'h1; // @[src/main/scala/utils/GTimer.scala 25:12]
  wire  _GEN_112 = ~_T_4 & ~_T_9 & _T_11 & _T_12 & _io_mem_req_valid_T_3 & _T_18 & _T_22 & DISPLAY_ENABLE; // @[src/main/scala/utils/Debug.scala 56:24]
  assign io_in_ready = io_out_ready & _T_50 & ~miss & _io_out_valid_T & io_mdReady & _hitWB_T_11; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 389:86]
  assign io_out_valid = io_in_valid & _io_out_valid_T_7; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 387:31]
  assign io_out_bits_addr = hit ? _io_out_bits_addr_T_7 : _io_out_bits_addr_T_26; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 386:26]
  assign io_out_bits_user = io_in_bits_user; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 385:15]
  assign io_mdWrite_wen = REG; // @[src/main/scala/nutcore/mem/TLB.scala 214:14]
  assign io_mdWrite_windex = REG_1; // @[src/main/scala/nutcore/mem/TLB.scala 215:17]
  assign io_mdWrite_waymask = REG_2; // @[src/main/scala/nutcore/mem/TLB.scala 216:18]
  assign io_mdWrite_wdata = {io_mdWrite_wdata_hi,io_mdWrite_wdata_lo}; // @[src/main/scala/nutcore/mem/TLB.scala 217:22]
  assign io_mem_req_valid = (state == 3'h1 | cmd) & ~isFlush; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 374:74]
  assign io_mem_req_bits_addr = hitWB ? hitData_pteaddr : raddr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 373:35]
  assign io_mem_req_bits_size = 3'h3; // @[src/main/scala/bus/simplebus/SimpleBus.scala 66:15]
  assign io_mem_req_bits_cmd = {{3'd0}, cmd}; // @[src/main/scala/bus/simplebus/SimpleBus.scala 65:14]
  assign io_mem_req_bits_wmask = 8'hff; // @[src/main/scala/bus/simplebus/SimpleBus.scala 68:16]
  assign io_mem_req_bits_wdata = hitWB ? {{24'd0}, hitWBStore} : memRespStore; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 373:138]
  assign io_mem_resp_ready = 1'h1; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 375:21]
  assign io_pf_loadPF = 1'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 242:16]
  assign io_pf_storePF = 1'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 243:17]
  assign io_ipf = hit ? hitinstrPF : missIPF; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 391:16]
  assign io_isFinish = _alreadyOutFire_T | _hitWB_T_9; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 392:30]
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/utils/LFSR64.scala 25:23]
      victimWaymask_lfsr <= 64'h1234567887654321; // @[src/main/scala/utils/LFSR64.scala 25:23]
    end else if (victimWaymask_lfsr == 64'h0) begin // @[src/main/scala/utils/LFSR64.scala 28:18]
      victimWaymask_lfsr <= 64'h1;
    end else begin
      victimWaymask_lfsr <= _victimWaymask_lfsr_T_2;
    end
    if (hitWB) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 228:29]
      hitWBStore <= _hitWBStore_T; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 228:29]
    end
    if (reset) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 253:22]
      state <= 3'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 253:22]
    end else if (3'h0 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 275:18]
      if (~io_flush & hitWB) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 277:32]
        state <= 3'h3; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 278:15]
      end else if (miss & _T_5) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 281:37]
        state <= 3'h1; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 282:15]
      end
    end else if (3'h1 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 275:18]
      if (isFlush) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 291:22]
        state <= 3'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 292:15]
      end else begin
        state <= _GEN_15;
      end
    end else if (3'h2 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 275:18]
      state <= _GEN_47;
    end else begin
      state <= _GEN_66;
    end
    if (reset) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 254:22]
      level <= 2'h3; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 254:22]
    end else if (3'h0 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 275:18]
      if (!(~io_flush & hitWB)) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 277:32]
        if (miss & _T_5) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 281:37]
          level <= 2'h3; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 284:15]
        end
      end
    end else if (!(3'h1 == state)) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 275:18]
      if (3'h2 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 275:18]
        level <= _GEN_56;
      end
    end
    if (!(3'h0 == state)) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 275:18]
      if (!(3'h1 == state)) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 275:18]
        if (3'h2 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 275:18]
          if (_T_12) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 299:31]
            memRespStore <= _GEN_43;
          end
        end
      end
    end
    if (!(3'h0 == state)) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 275:18]
      if (!(3'h1 == state)) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 275:18]
        if (3'h2 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 275:18]
          if (_T_12) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 299:31]
            missMaskStore <= _GEN_46;
          end
        end
      end
    end
    if (3'h0 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 275:18]
      if (!(~io_flush & hitWB)) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 277:32]
        if (miss & _T_5) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 281:37]
          raddr <= _raddr_T_1; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 283:15]
        end
      end
    end else if (!(3'h1 == state)) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 275:18]
      if (3'h2 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 275:18]
        if (_T_12) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 299:31]
          raddr <= _GEN_41;
        end
      end
    end
    if (reset) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 263:33]
      alreadyOutFire <= 1'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 263:33]
    end else if (3'h0 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 275:18]
      if (~io_flush & hitWB) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 277:32]
        alreadyOutFire <= 1'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 280:24]
      end else if (miss & _T_5) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 281:37]
        alreadyOutFire <= 1'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 286:24]
      end else begin
        alreadyOutFire <= _GEN_2;
      end
    end else if (3'h1 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 275:18]
      alreadyOutFire <= _GEN_2;
    end else if (3'h2 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 275:18]
      alreadyOutFire <= _GEN_2;
    end else begin
      alreadyOutFire <= _GEN_69;
    end
    if (reset) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 266:26]
      needFlush <= 1'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 266:26]
    end else if (3'h0 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 275:18]
      if (~io_flush & hitWB) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 277:32]
        needFlush <= 1'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 279:19]
      end else if (miss & _T_5) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 281:37]
        needFlush <= 1'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 285:19]
      end else begin
        needFlush <= _GEN_4;
      end
    end else if (3'h1 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 275:18]
      if (isFlush) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 291:22]
        needFlush <= 1'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 293:19]
      end else begin
        needFlush <= _GEN_4;
      end
    end else if (3'h2 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 275:18]
      needFlush <= _GEN_48;
    end else begin
      needFlush <= _GEN_67;
    end
    if (reset) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 272:24]
      missIPF <= 1'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 272:24]
    end else if (!(3'h0 == state)) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 275:18]
      if (!(3'h1 == state)) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 275:18]
        if (3'h2 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 275:18]
          missIPF <= _GEN_49;
        end else begin
          missIPF <= _GEN_68;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/GTimer.scala 24:20]
      c <= 64'h0; // @[src/main/scala/utils/GTimer.scala 24:20]
    end else begin
      c <= _c_T_1; // @[src/main/scala/utils/GTimer.scala 25:7]
    end
    if (reset) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 378:33]
      REG <= 1'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 378:33]
    end else begin
      REG <= missMetaRefill & _io_mem_req_valid_T_3 | hitWB & state == 3'h0 & _io_mem_req_valid_T_3; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 378:33]
    end
    REG_1 <= io_in_bits_addr[12]; // @[src/main/scala/nutcore/mem/TLB.scala 200:19]
    if (hit) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 214:20]
      REG_2 <= hitVec;
    end else begin
      REG_2 <= victimWaymask;
    end
    REG_3 <= {hitVec_hi,vpn_vpn0}; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 379:89]
    if (hitWB) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 380:23]
      REG_4 <= hitMeta_asid;
    end else begin
      REG_4 <= satp_asid;
    end
    if (hitWB) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 380:76]
      REG_5 <= hitMeta_mask;
    end else if (3'h0 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 275:18]
      REG_5 <= 18'h3ffff; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 257:26]
    end else if (3'h1 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 275:18]
      REG_5 <= 18'h3ffff; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 257:26]
    end else if (3'h2 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 275:18]
      REG_5 <= _GEN_54;
    end else begin
      REG_5 <= 18'h3ffff; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 257:26]
    end
    if (hitWB) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 381:23]
      REG_6 <= hitRefillFlag;
    end else if (3'h0 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 275:18]
      REG_6 <= 8'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 260:32]
    end else if (3'h1 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 275:18]
      REG_6 <= 8'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 260:32]
    end else if (3'h2 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 275:18]
      REG_6 <= _GEN_51;
    end else begin
      REG_6 <= 8'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 260:32]
    end
    if (hitWB) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 381:81]
      REG_7 <= hitData_ppn;
    end else begin
      REG_7 <= memRdata_ppn;
    end
    if (hitWB) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 382:27]
      REG_8 <= hitData_pteaddr;
    end else begin
      REG_8 <= raddr;
    end
    if (reset) begin // @[src/main/scala/utils/GTimer.scala 24:20]
      c_4 <= 64'h0; // @[src/main/scala/utils/GTimer.scala 24:20]
    end else begin
      c_4 <= _c_T_9; // @[src/main/scala/utils/GTimer.scala 25:7]
    end
    if (reset) begin // @[src/main/scala/utils/GTimer.scala 24:20]
      c_5 <= 64'h0; // @[src/main/scala/utils/GTimer.scala 24:20]
    end else begin
      c_5 <= _c_T_11; // @[src/main/scala/utils/GTimer.scala 25:7]
    end
    if (reset) begin // @[src/main/scala/utils/GTimer.scala 24:20]
      c_6 <= 64'h0; // @[src/main/scala/utils/GTimer.scala 24:20]
    end else begin
      c_6 <= _c_T_13; // @[src/main/scala/utils/GTimer.scala 25:7]
    end
    if (reset) begin // @[src/main/scala/utils/GTimer.scala 24:20]
      c_7 <= 64'h0; // @[src/main/scala/utils/GTimer.scala 24:20]
    end else begin
      c_7 <= _c_T_15; // @[src/main/scala/utils/GTimer.scala 25:7]
    end
    if (reset) begin // @[src/main/scala/utils/GTimer.scala 24:20]
      c_8 <= 64'h0; // @[src/main/scala/utils/GTimer.scala 24:20]
    end else begin
      c_8 <= _c_T_17; // @[src/main/scala/utils/GTimer.scala 25:7]
    end
    if (reset) begin // @[src/main/scala/utils/GTimer.scala 24:20]
      c_9 <= 64'h0; // @[src/main/scala/utils/GTimer.scala 24:20]
    end else begin
      c_9 <= _c_T_19; // @[src/main/scala/utils/GTimer.scala 25:7]
    end
    if (reset) begin // @[src/main/scala/utils/GTimer.scala 24:20]
      c_10 <= 64'h0; // @[src/main/scala/utils/GTimer.scala 24:20]
    end else begin
      c_10 <= _c_T_21; // @[src/main/scala/utils/GTimer.scala 25:7]
    end
    if (reset) begin // @[src/main/scala/utils/GTimer.scala 24:20]
      c_11 <= 64'h0; // @[src/main/scala/utils/GTimer.scala 24:20]
    end else begin
      c_11 <= _c_T_23; // @[src/main/scala/utils/GTimer.scala 25:7]
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~_T_4 & ~_T_9 & _T_11 & _T_12 & _io_mem_req_valid_T_3 & _T_18 & _T_22 & DISPLAY_ENABLE & ~reset) begin
          $fwrite(32'h80000002,"[%d] EmbeddedTLBExec: ",c); // @[src/main/scala/utils/Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_112 & _T_25) begin
          $fwrite(32'h80000002,"tlbException!!! "); // @[src/main/scala/utils/Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_112 & _T_25) begin
          $fwrite(32'h80000002,
            " req:addr = 0x%x, cmd = %d, size = %d, wmask = 0x%x, wdata = 0x%x  Memreq:DecoupledIO(ready -> %d, valid -> %d, bits -> addr = 0x%x, cmd = %d, size = %d, wmask = 0x%x, wdata = 0x%x)  MemResp:DecoupledIO(ready -> %d, valid -> %d, bits -> rdata = %x, cmd = %d)"
            ,io_in_bits_addr,4'h0,3'h3,8'h0,64'h0,io_mem_req_ready,io_mem_req_valid,io_mem_req_bits_addr,
            io_mem_req_bits_cmd,io_mem_req_bits_size,io_mem_req_bits_wmask,io_mem_req_bits_wdata,io_mem_resp_ready,
            io_mem_resp_valid,io_mem_resp_bits_rdata,io_mem_resp_bits_cmd); // @[src/main/scala/utils/Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_112 & _T_25) begin
          $fwrite(32'h80000002," level:%d",level); // @[src/main/scala/utils/Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_112 & _T_25) begin
          $fwrite(32'h80000002,"\n"); // @[src/main/scala/utils/Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & ~reset) begin
          $fwrite(32'h80000002,"[%d] EmbeddedTLBExec: ",c_4); // @[src/main/scala/utils/Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_25) begin
          $fwrite(32'h80000002,"In(%d, %d) Out(%d, %d) InAddr:%x OutAddr:%x cmd:%d \n",io_in_valid,io_in_ready,
            io_out_valid,io_out_ready,io_in_bits_addr,io_out_bits_addr,4'h0); // @[src/main/scala/utils/Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & ~reset) begin
          $fwrite(32'h80000002,"[%d] EmbeddedTLBExec: ",c_5); // @[src/main/scala/utils/Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_25) begin
          $fwrite(32'h80000002,"isAMO:%d io.Flush:%d needFlush:%d alreadyOutFire:%d isFinish:%d\n",1'h0,io_flush,
            needFlush,alreadyOutFire,io_isFinish); // @[src/main/scala/utils/Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & ~reset) begin
          $fwrite(32'h80000002,"[%d] EmbeddedTLBExec: ",c_6); // @[src/main/scala/utils/Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_25) begin
          $fwrite(32'h80000002,
            "hit:%d hitWB:%d hitVPN:%x hitFlag:%x hitPPN:%x hitRefillFlag:%x hitWBStore:%x hitCheck:%d hitExec:%d hitLoad:%d hitStore:%d\n"
            ,hit,hitWB,hitMeta_vpn,_hitRefillFlag_T_2,hitData_ppn,hitRefillFlag,hitWBStore,hitCheck,hitExec,hitLoad,
            hitStore); // @[src/main/scala/utils/Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & ~reset) begin
          $fwrite(32'h80000002,"[%d] EmbeddedTLBExec: ",c_7); // @[src/main/scala/utils/Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_25) begin
          $fwrite(32'h80000002,
            "miss:%d state:%d level:%d raddr:%x memRdata:%x missMask:%x missRefillFlag:%x missMetaRefill:%d\n",miss,
            state,level,raddr,_T_80,missMask,missRefillFlag,missMetaRefill); // @[src/main/scala/utils/Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & ~reset) begin
          $fwrite(32'h80000002,"[%d] EmbeddedTLBExec: ",c_8); // @[src/main/scala/utils/Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_25) begin
          $fwrite(32'h80000002,"meta/data: (0)%x|%b|%x (1)%x|%b|%x (2)%x|%b|%x (3)%x|%b|%x rread:%d\n",io_md_0[120:94],
            io_md_0[59:52],io_md_0[51:32],io_md_1[120:94],io_md_1[59:52],io_md_1[51:32],io_md_2[120:94],io_md_2[59:52],
            io_md_2[51:32],io_md_3[120:94],io_md_3[59:52],io_md_3[51:32],io_mdReady); // @[src/main/scala/utils/Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & ~reset) begin
          $fwrite(32'h80000002,"[%d] EmbeddedTLBExec: ",c_9); // @[src/main/scala/utils/Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_25) begin
          $fwrite(32'h80000002,
            "md: wen:%d windex:%x waymask:%x vpn:%x asid:%x mask:%x flag:%x asid:%x ppn:%x pteaddr:%x\n",io_mdWrite_wen,
            io_mdWrite_windex,io_mdWrite_waymask,io_mdWrite_wdata[120:94],io_mdWrite_wdata[93:78],io_mdWrite_wdata[77:60
            ],io_mdWrite_wdata[59:52],io_mdWrite_wdata[93:78],io_mdWrite_wdata[51:32],io_mdWrite_wdata[31:0]); // @[src/main/scala/utils/Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & ~reset) begin
          $fwrite(32'h80000002,"[%d] EmbeddedTLBExec: ",c_10); // @[src/main/scala/utils/Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_25) begin
          $fwrite(32'h80000002,"MemReq(%d, %d) MemResp(%d, %d) addr:%x cmd:%d rdata:%x cmd:%d\n",io_mem_req_valid,
            io_mem_req_ready,io_mem_resp_valid,io_mem_resp_ready,io_mem_req_bits_addr,io_mem_req_bits_cmd,
            io_mem_resp_bits_rdata,io_mem_resp_bits_cmd); // @[src/main/scala/utils/Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & ~reset) begin
          $fwrite(32'h80000002,"[%d] EmbeddedTLBExec: ",c_11); // @[src/main/scala/utils/Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_25) begin
          $fwrite(32'h80000002,"io.ipf:%d hitinstrPF:%d missIPF:%d pf.loadPF:%d pf.storePF:%d loadPF:%d storePF:%d\n",
            io_ipf,hitinstrPF,missIPF,io_pf_loadPF,io_pf_storePF,1'h0,1'h0); // @[src/main/scala/utils/Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  victimWaymask_lfsr = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  hitWBStore = _RAND_1[39:0];
  _RAND_2 = {1{`RANDOM}};
  state = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  level = _RAND_3[1:0];
  _RAND_4 = {2{`RANDOM}};
  memRespStore = _RAND_4[63:0];
  _RAND_5 = {1{`RANDOM}};
  missMaskStore = _RAND_5[17:0];
  _RAND_6 = {1{`RANDOM}};
  raddr = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  alreadyOutFire = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  needFlush = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  missIPF = _RAND_9[0:0];
  _RAND_10 = {2{`RANDOM}};
  c = _RAND_10[63:0];
  _RAND_11 = {1{`RANDOM}};
  REG = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  REG_1 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  REG_2 = _RAND_13[3:0];
  _RAND_14 = {1{`RANDOM}};
  REG_3 = _RAND_14[26:0];
  _RAND_15 = {1{`RANDOM}};
  REG_4 = _RAND_15[15:0];
  _RAND_16 = {1{`RANDOM}};
  REG_5 = _RAND_16[17:0];
  _RAND_17 = {1{`RANDOM}};
  REG_6 = _RAND_17[7:0];
  _RAND_18 = {1{`RANDOM}};
  REG_7 = _RAND_18[19:0];
  _RAND_19 = {1{`RANDOM}};
  REG_8 = _RAND_19[31:0];
  _RAND_20 = {2{`RANDOM}};
  c_4 = _RAND_20[63:0];
  _RAND_21 = {2{`RANDOM}};
  c_5 = _RAND_21[63:0];
  _RAND_22 = {2{`RANDOM}};
  c_6 = _RAND_22[63:0];
  _RAND_23 = {2{`RANDOM}};
  c_7 = _RAND_23[63:0];
  _RAND_24 = {2{`RANDOM}};
  c_8 = _RAND_24[63:0];
  _RAND_25 = {2{`RANDOM}};
  c_9 = _RAND_25[63:0];
  _RAND_26 = {2{`RANDOM}};
  c_10 = _RAND_26[63:0];
  _RAND_27 = {2{`RANDOM}};
  c_11 = _RAND_27[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module EmbeddedTLBMD(
  input          clock,
  input          reset,
  output [120:0] io_tlbmd_0, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 41:14]
  output [120:0] io_tlbmd_1, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 41:14]
  output [120:0] io_tlbmd_2, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 41:14]
  output [120:0] io_tlbmd_3, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 41:14]
  input          io_write_wen, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 41:14]
  input  [3:0]   io_write_waymask, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 41:14]
  input  [120:0] io_write_wdata, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 41:14]
  output         io_ready // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 41:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [127:0] _RAND_0;
  reg [127:0] _RAND_1;
  reg [127:0] _RAND_2;
  reg [127:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  reg [120:0] tlbmd_0_0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 49:18]
  reg [120:0] tlbmd_0_1; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 49:18]
  reg [120:0] tlbmd_0_2; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 49:18]
  reg [120:0] tlbmd_0_3; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 49:18]
  reg  resetState; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 53:27]
  wire  _GEN_1 = resetState ? 1'h0 : resetState; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 55:22 53:27 55:35]
  wire  wen = resetState | io_write_wen; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 62:16]
  wire [3:0] waymask = resetState ? 4'hf : io_write_waymask; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 64:20]
  assign io_tlbmd_0 = tlbmd_0_0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 50:12]
  assign io_tlbmd_1 = tlbmd_0_1; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 50:12]
  assign io_tlbmd_2 = tlbmd_0_2; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 50:12]
  assign io_tlbmd_3 = tlbmd_0_3; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 50:12]
  assign io_ready = ~resetState; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 74:15]
  always @(posedge clock) begin
    if (wen & waymask[0]) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 69:21]
      if (resetState) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 65:21]
        tlbmd_0_0 <= 121'h0;
      end else begin
        tlbmd_0_0 <= io_write_wdata;
      end
    end
    if (wen & waymask[1]) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 69:21]
      if (resetState) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 65:21]
        tlbmd_0_1 <= 121'h0;
      end else begin
        tlbmd_0_1 <= io_write_wdata;
      end
    end
    if (wen & waymask[2]) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 69:21]
      if (resetState) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 65:21]
        tlbmd_0_2 <= 121'h0;
      end else begin
        tlbmd_0_2 <= io_write_wdata;
      end
    end
    if (wen & waymask[3]) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 69:21]
      if (resetState) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 65:21]
        tlbmd_0_3 <= 121'h0;
      end else begin
        tlbmd_0_3 <= io_write_wdata;
      end
    end
    resetState <= reset | _GEN_1; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 53:{27,27}]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {4{`RANDOM}};
  tlbmd_0_0 = _RAND_0[120:0];
  _RAND_1 = {4{`RANDOM}};
  tlbmd_0_1 = _RAND_1[120:0];
  _RAND_2 = {4{`RANDOM}};
  tlbmd_0_2 = _RAND_2[120:0];
  _RAND_3 = {4{`RANDOM}};
  tlbmd_0_3 = _RAND_3[120:0];
  _RAND_4 = {1{`RANDOM}};
  resetState = _RAND_4[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module EmbeddedTLB(
  input         clock,
  input         reset,
  output        io_in_req_ready, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 37:14]
  input         io_in_req_valid, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 37:14]
  input  [38:0] io_in_req_bits_addr, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 37:14]
  input  [86:0] io_in_req_bits_user, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 37:14]
  input         io_in_resp_ready, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 37:14]
  output        io_in_resp_valid, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 37:14]
  output [3:0]  io_in_resp_bits_cmd, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 37:14]
  output [63:0] io_in_resp_bits_rdata, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 37:14]
  output [86:0] io_in_resp_bits_user, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 37:14]
  input         io_out_req_ready, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 37:14]
  output        io_out_req_valid, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 37:14]
  output [31:0] io_out_req_bits_addr, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 37:14]
  output [3:0]  io_out_req_bits_cmd, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 37:14]
  output [63:0] io_out_req_bits_wdata, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 37:14]
  output [86:0] io_out_req_bits_user, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 37:14]
  output        io_out_resp_ready, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 37:14]
  input         io_out_resp_valid, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 37:14]
  input  [63:0] io_out_resp_bits_rdata, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 37:14]
  input  [86:0] io_out_resp_bits_user, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 37:14]
  input         io_mem_req_ready, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 37:14]
  output        io_mem_req_valid, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 37:14]
  output [31:0] io_mem_req_bits_addr, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 37:14]
  output [3:0]  io_mem_req_bits_cmd, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 37:14]
  output [63:0] io_mem_req_bits_wdata, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 37:14]
  input         io_mem_resp_valid, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 37:14]
  input  [3:0]  io_mem_resp_bits_cmd, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 37:14]
  input  [63:0] io_mem_resp_bits_rdata, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 37:14]
  input         io_flush, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 37:14]
  input  [1:0]  io_csrMMU_priviledgeMode, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 37:14]
  output        io_csrMMU_loadPF, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 37:14]
  output        io_csrMMU_storePF, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 37:14]
  input         io_cacheEmpty, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 37:14]
  output        io_ipf, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 37:14]
  input  [63:0] CSRSATP,
  input         DISPLAY_ENABLE,
  input         MOUFlushTLB
);
`ifdef RANDOMIZE_REG_INIT
  reg [127:0] _RAND_0;
  reg [127:0] _RAND_1;
  reg [127:0] _RAND_2;
  reg [127:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [95:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [63:0] _RAND_10;
`endif // RANDOMIZE_REG_INIT
  wire  tlbExec_clock; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 85:23]
  wire  tlbExec_reset; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 85:23]
  wire  tlbExec_io_in_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 85:23]
  wire  tlbExec_io_in_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 85:23]
  wire [38:0] tlbExec_io_in_bits_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 85:23]
  wire [86:0] tlbExec_io_in_bits_user; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 85:23]
  wire  tlbExec_io_out_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 85:23]
  wire  tlbExec_io_out_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 85:23]
  wire [31:0] tlbExec_io_out_bits_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 85:23]
  wire [86:0] tlbExec_io_out_bits_user; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 85:23]
  wire [120:0] tlbExec_io_md_0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 85:23]
  wire [120:0] tlbExec_io_md_1; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 85:23]
  wire [120:0] tlbExec_io_md_2; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 85:23]
  wire [120:0] tlbExec_io_md_3; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 85:23]
  wire  tlbExec_io_mdWrite_wen; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 85:23]
  wire  tlbExec_io_mdWrite_windex; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 85:23]
  wire [3:0] tlbExec_io_mdWrite_waymask; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 85:23]
  wire [120:0] tlbExec_io_mdWrite_wdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 85:23]
  wire  tlbExec_io_mdReady; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 85:23]
  wire  tlbExec_io_mem_req_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 85:23]
  wire  tlbExec_io_mem_req_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 85:23]
  wire [31:0] tlbExec_io_mem_req_bits_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 85:23]
  wire [2:0] tlbExec_io_mem_req_bits_size; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 85:23]
  wire [3:0] tlbExec_io_mem_req_bits_cmd; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 85:23]
  wire [7:0] tlbExec_io_mem_req_bits_wmask; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 85:23]
  wire [63:0] tlbExec_io_mem_req_bits_wdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 85:23]
  wire  tlbExec_io_mem_resp_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 85:23]
  wire  tlbExec_io_mem_resp_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 85:23]
  wire [3:0] tlbExec_io_mem_resp_bits_cmd; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 85:23]
  wire [63:0] tlbExec_io_mem_resp_bits_rdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 85:23]
  wire  tlbExec_io_flush; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 85:23]
  wire [63:0] tlbExec_io_satp; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 85:23]
  wire [1:0] tlbExec_io_pf_priviledgeMode; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 85:23]
  wire  tlbExec_io_pf_loadPF; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 85:23]
  wire  tlbExec_io_pf_storePF; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 85:23]
  wire  tlbExec_io_ipf; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 85:23]
  wire  tlbExec_io_isFinish; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 85:23]
  wire  tlbExec_DISPLAY_ENABLE; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 85:23]
  wire  mdTLB_clock; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 87:21]
  wire  mdTLB_reset; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 87:21]
  wire [120:0] mdTLB_io_tlbmd_0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 87:21]
  wire [120:0] mdTLB_io_tlbmd_1; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 87:21]
  wire [120:0] mdTLB_io_tlbmd_2; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 87:21]
  wire [120:0] mdTLB_io_tlbmd_3; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 87:21]
  wire  mdTLB_io_write_wen; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 87:21]
  wire [3:0] mdTLB_io_write_waymask; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 87:21]
  wire [120:0] mdTLB_io_write_wdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 87:21]
  wire  mdTLB_io_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 87:21]
  reg [120:0] r_0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 94:29]
  reg [120:0] r_1; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 94:29]
  reg [120:0] r_2; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 94:29]
  reg [120:0] r_3; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 94:29]
  wire  mdUpdate = io_in_req_valid & tlbExec_io_in_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 119:26]
  wire  vmEnable = CSRSATP[63:60] == 4'h8 & io_csrMMU_priviledgeMode < 2'h3; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 107:57]
  reg  valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 110:24]
  wire  _GEN_4 = tlbExec_io_isFinish ? 1'h0 : valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 110:24 111:{25,33}]
  wire  _GEN_5 = mdUpdate & vmEnable | _GEN_4; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 112:{50,58}]
  reg [38:0] tlbExec_io_in_bits_r_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 116:28]
  reg [86:0] tlbExec_io_in_bits_r_user; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 116:28]
  wire  _GEN_13 = ~vmEnable | io_out_req_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 128:19 129:26 141:23]
  wire  _GEN_14 = ~vmEnable ? io_in_req_valid : tlbExec_io_out_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 128:19 131:22 141:23]
  wire  _T_3 = tlbExec_io_ipf & vmEnable; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 157:26]
  reg [63:0] c; // @[src/main/scala/utils/GTimer.scala 24:20]
  wire [63:0] _c_T_1 = c + 64'h1; // @[src/main/scala/utils/GTimer.scala 25:12]
  wire  _T_8 = ~reset; // @[src/main/scala/utils/Debug.scala 56:24]
  reg [63:0] c_1; // @[src/main/scala/utils/GTimer.scala 24:20]
  wire [63:0] _c_T_3 = c_1 + 64'h1; // @[src/main/scala/utils/GTimer.scala 25:12]
  reg [63:0] c_2; // @[src/main/scala/utils/GTimer.scala 24:20]
  wire [63:0] _c_T_5 = c_2 + 64'h1; // @[src/main/scala/utils/GTimer.scala 25:12]
  reg [63:0] c_3; // @[src/main/scala/utils/GTimer.scala 24:20]
  wire [63:0] _c_T_7 = c_3 + 64'h1; // @[src/main/scala/utils/GTimer.scala 25:12]
  EmbeddedTLBExec tlbExec ( // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 85:23]
    .clock(tlbExec_clock),
    .reset(tlbExec_reset),
    .io_in_ready(tlbExec_io_in_ready),
    .io_in_valid(tlbExec_io_in_valid),
    .io_in_bits_addr(tlbExec_io_in_bits_addr),
    .io_in_bits_user(tlbExec_io_in_bits_user),
    .io_out_ready(tlbExec_io_out_ready),
    .io_out_valid(tlbExec_io_out_valid),
    .io_out_bits_addr(tlbExec_io_out_bits_addr),
    .io_out_bits_user(tlbExec_io_out_bits_user),
    .io_md_0(tlbExec_io_md_0),
    .io_md_1(tlbExec_io_md_1),
    .io_md_2(tlbExec_io_md_2),
    .io_md_3(tlbExec_io_md_3),
    .io_mdWrite_wen(tlbExec_io_mdWrite_wen),
    .io_mdWrite_windex(tlbExec_io_mdWrite_windex),
    .io_mdWrite_waymask(tlbExec_io_mdWrite_waymask),
    .io_mdWrite_wdata(tlbExec_io_mdWrite_wdata),
    .io_mdReady(tlbExec_io_mdReady),
    .io_mem_req_ready(tlbExec_io_mem_req_ready),
    .io_mem_req_valid(tlbExec_io_mem_req_valid),
    .io_mem_req_bits_addr(tlbExec_io_mem_req_bits_addr),
    .io_mem_req_bits_size(tlbExec_io_mem_req_bits_size),
    .io_mem_req_bits_cmd(tlbExec_io_mem_req_bits_cmd),
    .io_mem_req_bits_wmask(tlbExec_io_mem_req_bits_wmask),
    .io_mem_req_bits_wdata(tlbExec_io_mem_req_bits_wdata),
    .io_mem_resp_ready(tlbExec_io_mem_resp_ready),
    .io_mem_resp_valid(tlbExec_io_mem_resp_valid),
    .io_mem_resp_bits_cmd(tlbExec_io_mem_resp_bits_cmd),
    .io_mem_resp_bits_rdata(tlbExec_io_mem_resp_bits_rdata),
    .io_flush(tlbExec_io_flush),
    .io_satp(tlbExec_io_satp),
    .io_pf_priviledgeMode(tlbExec_io_pf_priviledgeMode),
    .io_pf_loadPF(tlbExec_io_pf_loadPF),
    .io_pf_storePF(tlbExec_io_pf_storePF),
    .io_ipf(tlbExec_io_ipf),
    .io_isFinish(tlbExec_io_isFinish),
    .DISPLAY_ENABLE(tlbExec_DISPLAY_ENABLE)
  );
  EmbeddedTLBMD mdTLB ( // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 87:21]
    .clock(mdTLB_clock),
    .reset(mdTLB_reset),
    .io_tlbmd_0(mdTLB_io_tlbmd_0),
    .io_tlbmd_1(mdTLB_io_tlbmd_1),
    .io_tlbmd_2(mdTLB_io_tlbmd_2),
    .io_tlbmd_3(mdTLB_io_tlbmd_3),
    .io_write_wen(mdTLB_io_write_wen),
    .io_write_waymask(mdTLB_io_write_waymask),
    .io_write_wdata(mdTLB_io_write_wdata),
    .io_ready(mdTLB_io_ready)
  );
  assign io_in_req_ready = ~vmEnable ? io_out_req_ready : tlbExec_io_in_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 115:16 128:19 132:21]
  assign io_in_resp_valid = _T_3 & io_cacheEmpty | io_out_resp_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 143:15 162:56 163:24]
  assign io_in_resp_bits_cmd = 4'h6; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 143:15 162:56 165:27]
  assign io_in_resp_bits_rdata = _T_3 & io_cacheEmpty ? 64'h0 : io_out_resp_bits_rdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 143:15 162:56 164:29]
  assign io_in_resp_bits_user = _T_3 & io_cacheEmpty ? tlbExec_io_in_bits_user : io_out_resp_bits_user; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 143:15 162:56 166:34]
  assign io_out_req_valid = tlbExec_io_ipf & vmEnable ? 1'h0 : _GEN_14; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 157:39 159:24]
  assign io_out_req_bits_addr = ~vmEnable ? io_in_req_bits_addr[31:0] : tlbExec_io_out_bits_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 128:19 133:26 141:23]
  assign io_out_req_bits_cmd = 4'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 128:19 135:25 141:23]
  assign io_out_req_bits_wdata = 64'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 128:19 137:27 141:23]
  assign io_out_req_bits_user = ~vmEnable ? io_in_req_bits_user : tlbExec_io_out_bits_user; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 128:19 138:32 141:23]
  assign io_out_resp_ready = io_in_resp_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 143:15]
  assign io_mem_req_valid = tlbExec_io_mem_req_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 92:18]
  assign io_mem_req_bits_addr = tlbExec_io_mem_req_bits_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 92:18]
  assign io_mem_req_bits_cmd = tlbExec_io_mem_req_bits_cmd; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 92:18]
  assign io_mem_req_bits_wdata = tlbExec_io_mem_req_bits_wdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 92:18]
  assign io_csrMMU_loadPF = 1'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 93:17]
  assign io_csrMMU_storePF = 1'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 93:17]
  assign io_ipf = _T_3 & io_cacheEmpty & tlbExec_io_ipf; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 162:56 167:14 99:10]
  assign tlbExec_clock = clock;
  assign tlbExec_reset = reset;
  assign tlbExec_io_in_valid = valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 117:17]
  assign tlbExec_io_in_bits_addr = tlbExec_io_in_bits_r_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 116:16]
  assign tlbExec_io_in_bits_user = tlbExec_io_in_bits_r_user; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 116:16]
  assign tlbExec_io_out_ready = tlbExec_io_ipf & vmEnable ? io_cacheEmpty & io_in_resp_ready : _GEN_13; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 157:39 158:28]
  assign tlbExec_io_md_0 = r_0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 94:17]
  assign tlbExec_io_md_1 = r_1; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 94:17]
  assign tlbExec_io_md_2 = r_2; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 94:17]
  assign tlbExec_io_md_3 = r_3; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 94:17]
  assign tlbExec_io_mdReady = mdTLB_io_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 95:22]
  assign tlbExec_io_mem_req_ready = io_mem_req_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 92:18]
  assign tlbExec_io_mem_resp_valid = io_mem_resp_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 92:18]
  assign tlbExec_io_mem_resp_bits_cmd = io_mem_resp_bits_cmd; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 92:18]
  assign tlbExec_io_mem_resp_bits_rdata = io_mem_resp_bits_rdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 92:18]
  assign tlbExec_io_flush = io_flush; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 90:20]
  assign tlbExec_io_satp = CSRSATP; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 81:22]
  assign tlbExec_io_pf_priviledgeMode = io_csrMMU_priviledgeMode; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 93:17]
  assign tlbExec_DISPLAY_ENABLE = DISPLAY_ENABLE;
  assign mdTLB_clock = clock;
  assign mdTLB_reset = reset | MOUFlushTLB; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 104:31]
  assign mdTLB_io_write_wen = tlbExec_io_mdWrite_wen; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 97:18]
  assign mdTLB_io_write_waymask = tlbExec_io_mdWrite_waymask; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 97:18]
  assign mdTLB_io_write_wdata = tlbExec_io_mdWrite_wdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 97:18]
  always @(posedge clock) begin
    if (mdUpdate) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 94:29]
      r_0 <= mdTLB_io_tlbmd_0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 94:29]
    end
    if (mdUpdate) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 94:29]
      r_1 <= mdTLB_io_tlbmd_1; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 94:29]
    end
    if (mdUpdate) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 94:29]
      r_2 <= mdTLB_io_tlbmd_2; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 94:29]
    end
    if (mdUpdate) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 94:29]
      r_3 <= mdTLB_io_tlbmd_3; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 94:29]
    end
    if (reset) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 110:24]
      valid <= 1'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 110:24]
    end else if (io_flush) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:20]
      valid <= 1'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end else begin
      valid <= _GEN_5;
    end
    if (mdUpdate) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 116:28]
      tlbExec_io_in_bits_r_addr <= io_in_req_bits_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 116:28]
    end
    if (mdUpdate) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 116:28]
      tlbExec_io_in_bits_r_user <= io_in_req_bits_user; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 116:28]
    end
    if (reset) begin // @[src/main/scala/utils/GTimer.scala 24:20]
      c <= 64'h0; // @[src/main/scala/utils/GTimer.scala 24:20]
    end else begin
      c <= _c_T_1; // @[src/main/scala/utils/GTimer.scala 25:7]
    end
    if (reset) begin // @[src/main/scala/utils/GTimer.scala 24:20]
      c_1 <= 64'h0; // @[src/main/scala/utils/GTimer.scala 24:20]
    end else begin
      c_1 <= _c_T_3; // @[src/main/scala/utils/GTimer.scala 25:7]
    end
    if (reset) begin // @[src/main/scala/utils/GTimer.scala 24:20]
      c_2 <= 64'h0; // @[src/main/scala/utils/GTimer.scala 24:20]
    end else begin
      c_2 <= _c_T_5; // @[src/main/scala/utils/GTimer.scala 25:7]
    end
    if (reset) begin // @[src/main/scala/utils/GTimer.scala 24:20]
      c_3 <= 64'h0; // @[src/main/scala/utils/GTimer.scala 24:20]
    end else begin
      c_3 <= _c_T_7; // @[src/main/scala/utils/GTimer.scala 25:7]
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & ~reset) begin
          $fwrite(32'h80000002,"[%d] EmbeddedTLB: ",c); // @[src/main/scala/utils/Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_8) begin
          $fwrite(32'h80000002,"InReq(%d, %d) InResp(%d, %d) OutReq(%d, %d) OutResp(%d, %d) vmEnable:%d mode:%d\n",
            io_in_req_valid,io_in_req_ready,io_in_resp_valid,io_in_resp_ready,io_out_req_valid,io_out_req_ready,
            io_out_resp_valid,io_out_resp_ready,vmEnable,io_csrMMU_priviledgeMode); // @[src/main/scala/utils/Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & ~reset) begin
          $fwrite(32'h80000002,"[%d] EmbeddedTLB: ",c_1); // @[src/main/scala/utils/Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_8) begin
          $fwrite(32'h80000002,"InReq: addr:%x cmd:%d wdata:%x OutReq: addr:%x cmd:%x wdata:%x\n",io_in_req_bits_addr,4'h0
            ,64'h0,io_out_req_bits_addr,io_out_req_bits_cmd,io_out_req_bits_wdata); // @[src/main/scala/utils/Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & ~reset) begin
          $fwrite(32'h80000002,"[%d] EmbeddedTLB: ",c_2); // @[src/main/scala/utils/Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_8) begin
          $fwrite(32'h80000002,"OutResp: rdata:%x cmd:%x Inresp: rdata:%x cmd:%x\n",io_out_resp_bits_rdata,4'h6,
            io_in_resp_bits_rdata,io_in_resp_bits_cmd); // @[src/main/scala/utils/Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & ~reset) begin
          $fwrite(32'h80000002,"[%d] EmbeddedTLB: ",c_3); // @[src/main/scala/utils/Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_8) begin
          $fwrite(32'h80000002,"satp:%x flush:%d cacheEmpty:%d instrPF:%d loadPF:%d storePF:%d \n",CSRSATP,io_flush,
            io_cacheEmpty,io_ipf,io_csrMMU_loadPF,io_csrMMU_storePF); // @[src/main/scala/utils/Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {4{`RANDOM}};
  r_0 = _RAND_0[120:0];
  _RAND_1 = {4{`RANDOM}};
  r_1 = _RAND_1[120:0];
  _RAND_2 = {4{`RANDOM}};
  r_2 = _RAND_2[120:0];
  _RAND_3 = {4{`RANDOM}};
  r_3 = _RAND_3[120:0];
  _RAND_4 = {1{`RANDOM}};
  valid = _RAND_4[0:0];
  _RAND_5 = {2{`RANDOM}};
  tlbExec_io_in_bits_r_addr = _RAND_5[38:0];
  _RAND_6 = {3{`RANDOM}};
  tlbExec_io_in_bits_r_user = _RAND_6[86:0];
  _RAND_7 = {2{`RANDOM}};
  c = _RAND_7[63:0];
  _RAND_8 = {2{`RANDOM}};
  c_1 = _RAND_8[63:0];
  _RAND_9 = {2{`RANDOM}};
  c_2 = _RAND_9[63:0];
  _RAND_10 = {2{`RANDOM}};
  c_3 = _RAND_10[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module CacheStage1(
  input         clock,
  input         reset,
  output        io_in_ready, // @[src/main/scala/nutcore/mem/Cache.scala 133:14]
  input         io_in_valid, // @[src/main/scala/nutcore/mem/Cache.scala 133:14]
  input  [31:0] io_in_bits_addr, // @[src/main/scala/nutcore/mem/Cache.scala 133:14]
  input  [2:0]  io_in_bits_size, // @[src/main/scala/nutcore/mem/Cache.scala 133:14]
  input  [3:0]  io_in_bits_cmd, // @[src/main/scala/nutcore/mem/Cache.scala 133:14]
  input  [7:0]  io_in_bits_wmask, // @[src/main/scala/nutcore/mem/Cache.scala 133:14]
  input  [63:0] io_in_bits_wdata, // @[src/main/scala/nutcore/mem/Cache.scala 133:14]
  input  [86:0] io_in_bits_user, // @[src/main/scala/nutcore/mem/Cache.scala 133:14]
  input         io_out_ready, // @[src/main/scala/nutcore/mem/Cache.scala 133:14]
  output        io_out_valid, // @[src/main/scala/nutcore/mem/Cache.scala 133:14]
  output [31:0] io_out_bits_req_addr, // @[src/main/scala/nutcore/mem/Cache.scala 133:14]
  output [86:0] io_out_bits_req_user, // @[src/main/scala/nutcore/mem/Cache.scala 133:14]
  input         io_metaReadBus_req_ready, // @[src/main/scala/nutcore/mem/Cache.scala 133:14]
  output        io_metaReadBus_req_valid, // @[src/main/scala/nutcore/mem/Cache.scala 133:14]
  output [6:0]  io_metaReadBus_req_bits_setIdx, // @[src/main/scala/nutcore/mem/Cache.scala 133:14]
  input  [18:0] io_metaReadBus_resp_data_0_tag, // @[src/main/scala/nutcore/mem/Cache.scala 133:14]
  input         io_metaReadBus_resp_data_0_valid, // @[src/main/scala/nutcore/mem/Cache.scala 133:14]
  input         io_metaReadBus_resp_data_0_dirty, // @[src/main/scala/nutcore/mem/Cache.scala 133:14]
  input  [18:0] io_metaReadBus_resp_data_1_tag, // @[src/main/scala/nutcore/mem/Cache.scala 133:14]
  input         io_metaReadBus_resp_data_1_valid, // @[src/main/scala/nutcore/mem/Cache.scala 133:14]
  input         io_metaReadBus_resp_data_1_dirty, // @[src/main/scala/nutcore/mem/Cache.scala 133:14]
  input  [18:0] io_metaReadBus_resp_data_2_tag, // @[src/main/scala/nutcore/mem/Cache.scala 133:14]
  input         io_metaReadBus_resp_data_2_valid, // @[src/main/scala/nutcore/mem/Cache.scala 133:14]
  input         io_metaReadBus_resp_data_2_dirty, // @[src/main/scala/nutcore/mem/Cache.scala 133:14]
  input  [18:0] io_metaReadBus_resp_data_3_tag, // @[src/main/scala/nutcore/mem/Cache.scala 133:14]
  input         io_metaReadBus_resp_data_3_valid, // @[src/main/scala/nutcore/mem/Cache.scala 133:14]
  input         io_metaReadBus_resp_data_3_dirty, // @[src/main/scala/nutcore/mem/Cache.scala 133:14]
  input         io_dataReadBus_req_ready, // @[src/main/scala/nutcore/mem/Cache.scala 133:14]
  output        io_dataReadBus_req_valid, // @[src/main/scala/nutcore/mem/Cache.scala 133:14]
  output [9:0]  io_dataReadBus_req_bits_setIdx, // @[src/main/scala/nutcore/mem/Cache.scala 133:14]
  input  [63:0] io_dataReadBus_resp_data_0_data, // @[src/main/scala/nutcore/mem/Cache.scala 133:14]
  input  [63:0] io_dataReadBus_resp_data_1_data, // @[src/main/scala/nutcore/mem/Cache.scala 133:14]
  input  [63:0] io_dataReadBus_resp_data_2_data, // @[src/main/scala/nutcore/mem/Cache.scala 133:14]
  input  [63:0] io_dataReadBus_resp_data_3_data, // @[src/main/scala/nutcore/mem/Cache.scala 133:14]
  input         DISPLAY_ENABLE
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  wire  _T = io_in_ready & io_in_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  wire  _T_4 = ~reset; // @[src/main/scala/nutcore/mem/Cache.scala 135:37]
  reg [63:0] c; // @[src/main/scala/utils/GTimer.scala 24:20]
  wire [63:0] _c_T_1 = c + 64'h1; // @[src/main/scala/utils/GTimer.scala 25:12]
  wire  _T_7 = _T & DISPLAY_ENABLE; // @[src/main/scala/utils/Debug.scala 55:16]
  wire  _io_in_ready_T_1 = io_out_ready & io_out_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  reg [63:0] c_1; // @[src/main/scala/utils/GTimer.scala 24:20]
  wire [63:0] _c_T_3 = c_1 + 64'h1; // @[src/main/scala/utils/GTimer.scala 25:12]
  assign io_in_ready = (~io_in_valid | _io_in_ready_T_1) & io_metaReadBus_req_ready & io_dataReadBus_req_ready; // @[src/main/scala/nutcore/mem/Cache.scala 145:76]
  assign io_out_valid = io_in_valid & io_metaReadBus_req_ready & io_dataReadBus_req_ready; // @[src/main/scala/nutcore/mem/Cache.scala 144:59]
  assign io_out_bits_req_addr = io_in_bits_addr; // @[src/main/scala/nutcore/mem/Cache.scala 143:19]
  assign io_out_bits_req_user = io_in_bits_user; // @[src/main/scala/nutcore/mem/Cache.scala 143:19]
  assign io_metaReadBus_req_valid = io_in_valid & io_out_ready; // @[src/main/scala/nutcore/mem/Cache.scala 139:34]
  assign io_metaReadBus_req_bits_setIdx = io_in_bits_addr[12:6]; // @[src/main/scala/nutcore/mem/Cache.scala 77:45]
  assign io_dataReadBus_req_valid = io_in_valid & io_out_ready; // @[src/main/scala/nutcore/mem/Cache.scala 139:34]
  assign io_dataReadBus_req_bits_setIdx = {io_in_bits_addr[12:6],io_in_bits_addr[5:3]}; // @[src/main/scala/nutcore/mem/Cache.scala 78:35]
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/utils/GTimer.scala 24:20]
      c <= 64'h0; // @[src/main/scala/utils/GTimer.scala 24:20]
    end else begin
      c <= _c_T_1; // @[src/main/scala/utils/GTimer.scala 25:7]
    end
    if (reset) begin // @[src/main/scala/utils/GTimer.scala 24:20]
      c_1 <= 64'h0; // @[src/main/scala/utils/GTimer.scala 24:20]
    end else begin
      c_1 <= _c_T_3; // @[src/main/scala/utils/GTimer.scala 25:7]
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_7 & _T_4) begin
          $fwrite(32'h80000002,"[%d] CacheStage1: ",c); // @[src/main/scala/utils/Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_7 & _T_4) begin
          $fwrite(32'h80000002,"[L1$] cache stage1, addr in: %x, user: %x id: %x\n",io_in_bits_addr,io_in_bits_user,1'h0
            ); // @[src/main/scala/utils/Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_4) begin
          $fwrite(32'h80000002,"[%d] CacheStage1: ",c_1); // @[src/main/scala/utils/Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_4) begin
          $fwrite(32'h80000002,
            "in.ready = %d, in.valid = %d, out.valid = %d, out.ready = %d, addr = %x, cmd = %x, dataReadBus.req.valid = %d\n"
            ,io_in_ready,io_in_valid,io_out_valid,io_out_ready,io_in_bits_addr,4'h0,io_dataReadBus_req_valid); // @[src/main/scala/utils/Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  c = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  c_1 = _RAND_1[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module CacheStage2(
  input         clock,
  input         reset,
  output        io_in_ready, // @[src/main/scala/nutcore/mem/Cache.scala 171:14]
  input         io_in_valid, // @[src/main/scala/nutcore/mem/Cache.scala 171:14]
  input  [31:0] io_in_bits_req_addr, // @[src/main/scala/nutcore/mem/Cache.scala 171:14]
  input  [2:0]  io_in_bits_req_size, // @[src/main/scala/nutcore/mem/Cache.scala 171:14]
  input  [3:0]  io_in_bits_req_cmd, // @[src/main/scala/nutcore/mem/Cache.scala 171:14]
  input  [7:0]  io_in_bits_req_wmask, // @[src/main/scala/nutcore/mem/Cache.scala 171:14]
  input  [63:0] io_in_bits_req_wdata, // @[src/main/scala/nutcore/mem/Cache.scala 171:14]
  input  [86:0] io_in_bits_req_user, // @[src/main/scala/nutcore/mem/Cache.scala 171:14]
  input         io_out_ready, // @[src/main/scala/nutcore/mem/Cache.scala 171:14]
  output        io_out_valid, // @[src/main/scala/nutcore/mem/Cache.scala 171:14]
  output [31:0] io_out_bits_req_addr, // @[src/main/scala/nutcore/mem/Cache.scala 171:14]
  output [86:0] io_out_bits_req_user, // @[src/main/scala/nutcore/mem/Cache.scala 171:14]
  output [18:0] io_out_bits_metas_0_tag, // @[src/main/scala/nutcore/mem/Cache.scala 171:14]
  output        io_out_bits_metas_0_valid, // @[src/main/scala/nutcore/mem/Cache.scala 171:14]
  output        io_out_bits_metas_0_dirty, // @[src/main/scala/nutcore/mem/Cache.scala 171:14]
  output [18:0] io_out_bits_metas_1_tag, // @[src/main/scala/nutcore/mem/Cache.scala 171:14]
  output        io_out_bits_metas_1_valid, // @[src/main/scala/nutcore/mem/Cache.scala 171:14]
  output        io_out_bits_metas_1_dirty, // @[src/main/scala/nutcore/mem/Cache.scala 171:14]
  output [18:0] io_out_bits_metas_2_tag, // @[src/main/scala/nutcore/mem/Cache.scala 171:14]
  output        io_out_bits_metas_2_valid, // @[src/main/scala/nutcore/mem/Cache.scala 171:14]
  output        io_out_bits_metas_2_dirty, // @[src/main/scala/nutcore/mem/Cache.scala 171:14]
  output [18:0] io_out_bits_metas_3_tag, // @[src/main/scala/nutcore/mem/Cache.scala 171:14]
  output        io_out_bits_metas_3_valid, // @[src/main/scala/nutcore/mem/Cache.scala 171:14]
  output        io_out_bits_metas_3_dirty, // @[src/main/scala/nutcore/mem/Cache.scala 171:14]
  output [63:0] io_out_bits_datas_0_data, // @[src/main/scala/nutcore/mem/Cache.scala 171:14]
  output [63:0] io_out_bits_datas_1_data, // @[src/main/scala/nutcore/mem/Cache.scala 171:14]
  output [63:0] io_out_bits_datas_2_data, // @[src/main/scala/nutcore/mem/Cache.scala 171:14]
  output [63:0] io_out_bits_datas_3_data, // @[src/main/scala/nutcore/mem/Cache.scala 171:14]
  output        io_out_bits_hit, // @[src/main/scala/nutcore/mem/Cache.scala 171:14]
  output [3:0]  io_out_bits_waymask, // @[src/main/scala/nutcore/mem/Cache.scala 171:14]
  output        io_out_bits_mmio, // @[src/main/scala/nutcore/mem/Cache.scala 171:14]
  output        io_out_bits_isForwardData, // @[src/main/scala/nutcore/mem/Cache.scala 171:14]
  output [63:0] io_out_bits_forwardData_data_data, // @[src/main/scala/nutcore/mem/Cache.scala 171:14]
  output [3:0]  io_out_bits_forwardData_waymask, // @[src/main/scala/nutcore/mem/Cache.scala 171:14]
  input  [18:0] io_metaReadResp_0_tag, // @[src/main/scala/nutcore/mem/Cache.scala 171:14]
  input         io_metaReadResp_0_valid, // @[src/main/scala/nutcore/mem/Cache.scala 171:14]
  input         io_metaReadResp_0_dirty, // @[src/main/scala/nutcore/mem/Cache.scala 171:14]
  input  [18:0] io_metaReadResp_1_tag, // @[src/main/scala/nutcore/mem/Cache.scala 171:14]
  input         io_metaReadResp_1_valid, // @[src/main/scala/nutcore/mem/Cache.scala 171:14]
  input         io_metaReadResp_1_dirty, // @[src/main/scala/nutcore/mem/Cache.scala 171:14]
  input  [18:0] io_metaReadResp_2_tag, // @[src/main/scala/nutcore/mem/Cache.scala 171:14]
  input         io_metaReadResp_2_valid, // @[src/main/scala/nutcore/mem/Cache.scala 171:14]
  input         io_metaReadResp_2_dirty, // @[src/main/scala/nutcore/mem/Cache.scala 171:14]
  input  [18:0] io_metaReadResp_3_tag, // @[src/main/scala/nutcore/mem/Cache.scala 171:14]
  input         io_metaReadResp_3_valid, // @[src/main/scala/nutcore/mem/Cache.scala 171:14]
  input         io_metaReadResp_3_dirty, // @[src/main/scala/nutcore/mem/Cache.scala 171:14]
  input  [63:0] io_dataReadResp_0_data, // @[src/main/scala/nutcore/mem/Cache.scala 171:14]
  input  [63:0] io_dataReadResp_1_data, // @[src/main/scala/nutcore/mem/Cache.scala 171:14]
  input  [63:0] io_dataReadResp_2_data, // @[src/main/scala/nutcore/mem/Cache.scala 171:14]
  input  [63:0] io_dataReadResp_3_data, // @[src/main/scala/nutcore/mem/Cache.scala 171:14]
  input         io_metaWriteBus_req_valid, // @[src/main/scala/nutcore/mem/Cache.scala 171:14]
  input  [6:0]  io_metaWriteBus_req_bits_setIdx, // @[src/main/scala/nutcore/mem/Cache.scala 171:14]
  input  [18:0] io_metaWriteBus_req_bits_data_tag, // @[src/main/scala/nutcore/mem/Cache.scala 171:14]
  input         io_metaWriteBus_req_bits_data_dirty, // @[src/main/scala/nutcore/mem/Cache.scala 171:14]
  input  [3:0]  io_metaWriteBus_req_bits_waymask, // @[src/main/scala/nutcore/mem/Cache.scala 171:14]
  input         io_dataWriteBus_req_valid, // @[src/main/scala/nutcore/mem/Cache.scala 171:14]
  input  [9:0]  io_dataWriteBus_req_bits_setIdx, // @[src/main/scala/nutcore/mem/Cache.scala 171:14]
  input  [63:0] io_dataWriteBus_req_bits_data_data, // @[src/main/scala/nutcore/mem/Cache.scala 171:14]
  input  [3:0]  io_dataWriteBus_req_bits_waymask, // @[src/main/scala/nutcore/mem/Cache.scala 171:14]
  input         DISPLAY_ENABLE
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [63:0] _RAND_12;
  reg [63:0] _RAND_13;
  reg [63:0] _RAND_14;
  reg [63:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [63:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [63:0] _RAND_19;
  reg [63:0] _RAND_20;
`endif // RANDOMIZE_REG_INIT
  wire [2:0] addr_wordIndex = io_in_bits_req_addr[5:3]; // @[src/main/scala/nutcore/mem/Cache.scala 174:31]
  wire [6:0] addr_index = io_in_bits_req_addr[12:6]; // @[src/main/scala/nutcore/mem/Cache.scala 174:31]
  wire [18:0] addr_tag = io_in_bits_req_addr[31:13]; // @[src/main/scala/nutcore/mem/Cache.scala 174:31]
  wire  isForwardMeta = io_in_valid & io_metaWriteBus_req_valid & io_metaWriteBus_req_bits_setIdx == addr_index; // @[src/main/scala/nutcore/mem/Cache.scala 176:64]
  reg  isForwardMetaReg; // @[src/main/scala/nutcore/mem/Cache.scala 177:33]
  wire  _GEN_0 = isForwardMeta | isForwardMetaReg; // @[src/main/scala/nutcore/mem/Cache.scala 178:24 177:33 178:43]
  wire  _T = io_in_ready & io_in_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  wire  _T_1 = ~io_in_valid; // @[src/main/scala/nutcore/mem/Cache.scala 179:23]
  wire  _T_2 = _T | ~io_in_valid; // @[src/main/scala/nutcore/mem/Cache.scala 179:20]
  reg [18:0] forwardMetaReg_data_tag; // @[src/main/scala/nutcore/mem/Cache.scala 180:33]
  reg  forwardMetaReg_data_dirty; // @[src/main/scala/nutcore/mem/Cache.scala 180:33]
  reg [3:0] forwardMetaReg_waymask; // @[src/main/scala/nutcore/mem/Cache.scala 180:33]
  wire [18:0] _GEN_3 = isForwardMeta ? io_metaWriteBus_req_bits_data_tag : forwardMetaReg_data_tag; // @[src/main/scala/nutcore/mem/Cache.scala 180:{33,33,33}]
  wire  _GEN_5 = isForwardMeta ? io_metaWriteBus_req_bits_data_dirty : forwardMetaReg_data_dirty; // @[src/main/scala/nutcore/mem/Cache.scala 180:{33,33,33}]
  wire [3:0] _GEN_6 = isForwardMeta ? io_metaWriteBus_req_bits_waymask : forwardMetaReg_waymask; // @[src/main/scala/nutcore/mem/Cache.scala 180:{33,33,33}]
  wire  pickForwardMeta = isForwardMetaReg | isForwardMeta; // @[src/main/scala/nutcore/mem/Cache.scala 183:42]
  wire  forwardWaymask_0 = _GEN_6[0]; // @[src/main/scala/nutcore/mem/Cache.scala 185:61]
  wire  forwardWaymask_1 = _GEN_6[1]; // @[src/main/scala/nutcore/mem/Cache.scala 185:61]
  wire  forwardWaymask_2 = _GEN_6[2]; // @[src/main/scala/nutcore/mem/Cache.scala 185:61]
  wire  forwardWaymask_3 = _GEN_6[3]; // @[src/main/scala/nutcore/mem/Cache.scala 185:61]
  wire [18:0] metaWay_0_tag = pickForwardMeta & forwardWaymask_0 ? _GEN_3 : io_metaReadResp_0_tag; // @[src/main/scala/nutcore/mem/Cache.scala 187:22]
  wire  metaWay_0_valid = pickForwardMeta & forwardWaymask_0 | io_metaReadResp_0_valid; // @[src/main/scala/nutcore/mem/Cache.scala 187:22]
  wire [18:0] metaWay_1_tag = pickForwardMeta & forwardWaymask_1 ? _GEN_3 : io_metaReadResp_1_tag; // @[src/main/scala/nutcore/mem/Cache.scala 187:22]
  wire  metaWay_1_valid = pickForwardMeta & forwardWaymask_1 | io_metaReadResp_1_valid; // @[src/main/scala/nutcore/mem/Cache.scala 187:22]
  wire [18:0] metaWay_2_tag = pickForwardMeta & forwardWaymask_2 ? _GEN_3 : io_metaReadResp_2_tag; // @[src/main/scala/nutcore/mem/Cache.scala 187:22]
  wire  metaWay_2_valid = pickForwardMeta & forwardWaymask_2 | io_metaReadResp_2_valid; // @[src/main/scala/nutcore/mem/Cache.scala 187:22]
  wire [18:0] metaWay_3_tag = pickForwardMeta & forwardWaymask_3 ? _GEN_3 : io_metaReadResp_3_tag; // @[src/main/scala/nutcore/mem/Cache.scala 187:22]
  wire  metaWay_3_valid = pickForwardMeta & forwardWaymask_3 | io_metaReadResp_3_valid; // @[src/main/scala/nutcore/mem/Cache.scala 187:22]
  wire  _hitVec_T_2 = metaWay_0_valid & metaWay_0_tag == addr_tag & io_in_valid; // @[src/main/scala/nutcore/mem/Cache.scala 190:73]
  wire  _hitVec_T_5 = metaWay_1_valid & metaWay_1_tag == addr_tag & io_in_valid; // @[src/main/scala/nutcore/mem/Cache.scala 190:73]
  wire  _hitVec_T_8 = metaWay_2_valid & metaWay_2_tag == addr_tag & io_in_valid; // @[src/main/scala/nutcore/mem/Cache.scala 190:73]
  wire  _hitVec_T_11 = metaWay_3_valid & metaWay_3_tag == addr_tag & io_in_valid; // @[src/main/scala/nutcore/mem/Cache.scala 190:73]
  wire [3:0] hitVec = {_hitVec_T_11,_hitVec_T_8,_hitVec_T_5,_hitVec_T_2}; // @[src/main/scala/nutcore/mem/Cache.scala 190:90]
  reg [63:0] victimWaymask_lfsr; // @[src/main/scala/utils/LFSR64.scala 25:23]
  wire  victimWaymask_xor = victimWaymask_lfsr[0] ^ victimWaymask_lfsr[1] ^ victimWaymask_lfsr[3] ^ victimWaymask_lfsr[4
    ]; // @[src/main/scala/utils/LFSR64.scala 26:43]
  wire [63:0] _victimWaymask_lfsr_T_2 = {victimWaymask_xor,victimWaymask_lfsr[63:1]}; // @[src/main/scala/utils/LFSR64.scala 28:41]
  wire [3:0] victimWaymask = 4'h1 << victimWaymask_lfsr[1:0]; // @[src/main/scala/nutcore/mem/Cache.scala 191:42]
  wire  _invalidVec_T = ~metaWay_0_valid; // @[src/main/scala/nutcore/mem/Cache.scala 193:45]
  wire  _invalidVec_T_1 = ~metaWay_1_valid; // @[src/main/scala/nutcore/mem/Cache.scala 193:45]
  wire  _invalidVec_T_2 = ~metaWay_2_valid; // @[src/main/scala/nutcore/mem/Cache.scala 193:45]
  wire  _invalidVec_T_3 = ~metaWay_3_valid; // @[src/main/scala/nutcore/mem/Cache.scala 193:45]
  wire [3:0] invalidVec = {_invalidVec_T_3,_invalidVec_T_2,_invalidVec_T_1,_invalidVec_T}; // @[src/main/scala/nutcore/mem/Cache.scala 193:56]
  wire  hasInvalidWay = |invalidVec; // @[src/main/scala/nutcore/mem/Cache.scala 194:34]
  wire [1:0] _refillInvalidWaymask_T_3 = invalidVec >= 4'h2 ? 2'h2 : 2'h1; // @[src/main/scala/nutcore/mem/Cache.scala 197:8]
  wire [2:0] _refillInvalidWaymask_T_4 = invalidVec >= 4'h4 ? 3'h4 : {{1'd0}, _refillInvalidWaymask_T_3}; // @[src/main/scala/nutcore/mem/Cache.scala 196:8]
  wire [3:0] refillInvalidWaymask = invalidVec >= 4'h8 ? 4'h8 : {{1'd0}, _refillInvalidWaymask_T_4}; // @[src/main/scala/nutcore/mem/Cache.scala 195:33]
  wire [3:0] _waymask_T = hasInvalidWay ? refillInvalidWaymask : victimWaymask; // @[src/main/scala/nutcore/mem/Cache.scala 200:49]
  wire [3:0] waymask = io_out_bits_hit ? hitVec : _waymask_T; // @[src/main/scala/nutcore/mem/Cache.scala 200:20]
  wire [1:0] _T_7 = waymask[0] + waymask[1]; // @[src/main/scala/nutcore/mem/Cache.scala 201:16]
  wire [1:0] _T_9 = waymask[2] + waymask[3]; // @[src/main/scala/nutcore/mem/Cache.scala 201:16]
  wire [2:0] _T_11 = _T_7 + _T_9; // @[src/main/scala/nutcore/mem/Cache.scala 201:16]
  wire  _T_13 = _T_11 > 3'h1; // @[src/main/scala/nutcore/mem/Cache.scala 201:26]
  reg [63:0] c; // @[src/main/scala/utils/GTimer.scala 24:20]
  wire [63:0] _c_T_1 = c + 64'h1; // @[src/main/scala/utils/GTimer.scala 25:12]
  wire  _T_16 = ~reset; // @[src/main/scala/utils/Debug.scala 56:24]
  reg [63:0] c_1; // @[src/main/scala/utils/GTimer.scala 24:20]
  wire [63:0] _c_T_3 = c_1 + 64'h1; // @[src/main/scala/utils/GTimer.scala 25:12]
  reg [63:0] c_2; // @[src/main/scala/utils/GTimer.scala 24:20]
  wire [63:0] _c_T_5 = c_2 + 64'h1; // @[src/main/scala/utils/GTimer.scala 25:12]
  reg [63:0] c_3; // @[src/main/scala/utils/GTimer.scala 24:20]
  wire [63:0] _c_T_7 = c_3 + 64'h1; // @[src/main/scala/utils/GTimer.scala 25:12]
  reg [63:0] c_4; // @[src/main/scala/utils/GTimer.scala 24:20]
  wire [63:0] _c_T_9 = c_4 + 64'h1; // @[src/main/scala/utils/GTimer.scala 25:12]
  reg [63:0] c_5; // @[src/main/scala/utils/GTimer.scala 24:20]
  wire [63:0] _c_T_11 = c_5 + 64'h1; // @[src/main/scala/utils/GTimer.scala 25:12]
  reg [63:0] c_6; // @[src/main/scala/utils/GTimer.scala 24:20]
  wire [63:0] _c_T_13 = c_6 + 64'h1; // @[src/main/scala/utils/GTimer.scala 25:12]
  reg [63:0] c_7; // @[src/main/scala/utils/GTimer.scala 24:20]
  wire [63:0] _c_T_15 = c_7 + 64'h1; // @[src/main/scala/utils/GTimer.scala 25:12]
  reg [63:0] c_8; // @[src/main/scala/utils/GTimer.scala 24:20]
  wire [63:0] _c_T_17 = c_8 + 64'h1; // @[src/main/scala/utils/GTimer.scala 25:12]
  reg [63:0] c_9; // @[src/main/scala/utils/GTimer.scala 24:20]
  wire [63:0] _c_T_19 = c_9 + 64'h1; // @[src/main/scala/utils/GTimer.scala 25:12]
  reg [63:0] c_10; // @[src/main/scala/utils/GTimer.scala 24:20]
  wire [63:0] _c_T_21 = c_10 + 64'h1; // @[src/main/scala/utils/GTimer.scala 25:12]
  wire [31:0] _io_out_bits_mmio_T = io_in_bits_req_addr ^ 32'h30000000; // @[src/main/scala/nutcore/NutCore.scala 87:11]
  wire  _io_out_bits_mmio_T_2 = _io_out_bits_mmio_T[31:28] == 4'h0; // @[src/main/scala/nutcore/NutCore.scala 87:44]
  wire [31:0] _io_out_bits_mmio_T_3 = io_in_bits_req_addr ^ 32'h40000000; // @[src/main/scala/nutcore/NutCore.scala 87:11]
  wire  _io_out_bits_mmio_T_5 = _io_out_bits_mmio_T_3[31:30] == 2'h0; // @[src/main/scala/nutcore/NutCore.scala 87:44]
  wire [9:0] _isForwardData_T_8 = {addr_index,addr_wordIndex}; // @[src/main/scala/nutcore/mem/Cache.scala 78:35]
  wire  _isForwardData_T_10 = io_dataWriteBus_req_valid & io_dataWriteBus_req_bits_setIdx == _isForwardData_T_8; // @[src/main/scala/nutcore/mem/Cache.scala 217:13]
  wire  isForwardData = io_in_valid & _isForwardData_T_10; // @[src/main/scala/nutcore/mem/Cache.scala 216:35]
  reg  isForwardDataReg; // @[src/main/scala/nutcore/mem/Cache.scala 219:33]
  wire  _GEN_8 = isForwardData | isForwardDataReg; // @[src/main/scala/nutcore/mem/Cache.scala 220:24 219:33 220:43]
  reg [63:0] forwardDataReg_data_data; // @[src/main/scala/nutcore/mem/Cache.scala 222:33]
  reg [3:0] forwardDataReg_waymask; // @[src/main/scala/nutcore/mem/Cache.scala 222:33]
  wire  _io_in_ready_T_1 = io_out_ready & io_out_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  reg [63:0] c_11; // @[src/main/scala/utils/GTimer.scala 24:20]
  wire [63:0] _c_T_23 = c_11 + 64'h1; // @[src/main/scala/utils/GTimer.scala 25:12]
  reg [63:0] c_12; // @[src/main/scala/utils/GTimer.scala 24:20]
  wire [63:0] _c_T_25 = c_12 + 64'h1; // @[src/main/scala/utils/GTimer.scala 25:12]
  wire  _GEN_13 = _T_13 & DISPLAY_ENABLE; // @[src/main/scala/utils/Debug.scala 56:24]
  assign io_in_ready = _T_1 | _io_in_ready_T_1; // @[src/main/scala/nutcore/mem/Cache.scala 228:31]
  assign io_out_valid = io_in_valid; // @[src/main/scala/nutcore/mem/Cache.scala 227:16]
  assign io_out_bits_req_addr = io_in_bits_req_addr; // @[src/main/scala/nutcore/mem/Cache.scala 226:19]
  assign io_out_bits_req_user = io_in_bits_req_user; // @[src/main/scala/nutcore/mem/Cache.scala 226:19]
  assign io_out_bits_metas_0_tag = pickForwardMeta & forwardWaymask_0 ? _GEN_3 : io_metaReadResp_0_tag; // @[src/main/scala/nutcore/mem/Cache.scala 187:22]
  assign io_out_bits_metas_0_valid = pickForwardMeta & forwardWaymask_0 | io_metaReadResp_0_valid; // @[src/main/scala/nutcore/mem/Cache.scala 187:22]
  assign io_out_bits_metas_0_dirty = pickForwardMeta & forwardWaymask_0 ? _GEN_5 : io_metaReadResp_0_dirty; // @[src/main/scala/nutcore/mem/Cache.scala 187:22]
  assign io_out_bits_metas_1_tag = pickForwardMeta & forwardWaymask_1 ? _GEN_3 : io_metaReadResp_1_tag; // @[src/main/scala/nutcore/mem/Cache.scala 187:22]
  assign io_out_bits_metas_1_valid = pickForwardMeta & forwardWaymask_1 | io_metaReadResp_1_valid; // @[src/main/scala/nutcore/mem/Cache.scala 187:22]
  assign io_out_bits_metas_1_dirty = pickForwardMeta & forwardWaymask_1 ? _GEN_5 : io_metaReadResp_1_dirty; // @[src/main/scala/nutcore/mem/Cache.scala 187:22]
  assign io_out_bits_metas_2_tag = pickForwardMeta & forwardWaymask_2 ? _GEN_3 : io_metaReadResp_2_tag; // @[src/main/scala/nutcore/mem/Cache.scala 187:22]
  assign io_out_bits_metas_2_valid = pickForwardMeta & forwardWaymask_2 | io_metaReadResp_2_valid; // @[src/main/scala/nutcore/mem/Cache.scala 187:22]
  assign io_out_bits_metas_2_dirty = pickForwardMeta & forwardWaymask_2 ? _GEN_5 : io_metaReadResp_2_dirty; // @[src/main/scala/nutcore/mem/Cache.scala 187:22]
  assign io_out_bits_metas_3_tag = pickForwardMeta & forwardWaymask_3 ? _GEN_3 : io_metaReadResp_3_tag; // @[src/main/scala/nutcore/mem/Cache.scala 187:22]
  assign io_out_bits_metas_3_valid = pickForwardMeta & forwardWaymask_3 | io_metaReadResp_3_valid; // @[src/main/scala/nutcore/mem/Cache.scala 187:22]
  assign io_out_bits_metas_3_dirty = pickForwardMeta & forwardWaymask_3 ? _GEN_5 : io_metaReadResp_3_dirty; // @[src/main/scala/nutcore/mem/Cache.scala 187:22]
  assign io_out_bits_datas_0_data = io_dataReadResp_0_data; // @[src/main/scala/nutcore/mem/Cache.scala 213:21]
  assign io_out_bits_datas_1_data = io_dataReadResp_1_data; // @[src/main/scala/nutcore/mem/Cache.scala 213:21]
  assign io_out_bits_datas_2_data = io_dataReadResp_2_data; // @[src/main/scala/nutcore/mem/Cache.scala 213:21]
  assign io_out_bits_datas_3_data = io_dataReadResp_3_data; // @[src/main/scala/nutcore/mem/Cache.scala 213:21]
  assign io_out_bits_hit = io_in_valid & |hitVec; // @[src/main/scala/nutcore/mem/Cache.scala 211:34]
  assign io_out_bits_waymask = io_out_bits_hit ? hitVec : _waymask_T; // @[src/main/scala/nutcore/mem/Cache.scala 200:20]
  assign io_out_bits_mmio = _io_out_bits_mmio_T_2 | _io_out_bits_mmio_T_5; // @[src/main/scala/nutcore/NutCore.scala 88:15]
  assign io_out_bits_isForwardData = isForwardDataReg | isForwardData; // @[src/main/scala/nutcore/mem/Cache.scala 223:49]
  assign io_out_bits_forwardData_data_data = isForwardData ? io_dataWriteBus_req_bits_data_data :
    forwardDataReg_data_data; // @[src/main/scala/nutcore/mem/Cache.scala 224:33]
  assign io_out_bits_forwardData_waymask = isForwardData ? io_dataWriteBus_req_bits_waymask : forwardDataReg_waymask; // @[src/main/scala/nutcore/mem/Cache.scala 224:33]
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/nutcore/mem/Cache.scala 177:33]
      isForwardMetaReg <= 1'h0; // @[src/main/scala/nutcore/mem/Cache.scala 177:33]
    end else if (_T | ~io_in_valid) begin // @[src/main/scala/nutcore/mem/Cache.scala 179:37]
      isForwardMetaReg <= 1'h0; // @[src/main/scala/nutcore/mem/Cache.scala 179:56]
    end else begin
      isForwardMetaReg <= _GEN_0;
    end
    if (isForwardMeta) begin // @[src/main/scala/nutcore/mem/Cache.scala 180:33]
      forwardMetaReg_data_tag <= io_metaWriteBus_req_bits_data_tag; // @[src/main/scala/nutcore/mem/Cache.scala 180:33]
    end
    if (isForwardMeta) begin // @[src/main/scala/nutcore/mem/Cache.scala 180:33]
      forwardMetaReg_data_dirty <= io_metaWriteBus_req_bits_data_dirty; // @[src/main/scala/nutcore/mem/Cache.scala 180:33]
    end
    if (isForwardMeta) begin // @[src/main/scala/nutcore/mem/Cache.scala 180:33]
      forwardMetaReg_waymask <= io_metaWriteBus_req_bits_waymask; // @[src/main/scala/nutcore/mem/Cache.scala 180:33]
    end
    if (reset) begin // @[src/main/scala/utils/LFSR64.scala 25:23]
      victimWaymask_lfsr <= 64'h1234567887654321; // @[src/main/scala/utils/LFSR64.scala 25:23]
    end else if (victimWaymask_lfsr == 64'h0) begin // @[src/main/scala/utils/LFSR64.scala 28:18]
      victimWaymask_lfsr <= 64'h1;
    end else begin
      victimWaymask_lfsr <= _victimWaymask_lfsr_T_2;
    end
    if (reset) begin // @[src/main/scala/utils/GTimer.scala 24:20]
      c <= 64'h0; // @[src/main/scala/utils/GTimer.scala 24:20]
    end else begin
      c <= _c_T_1; // @[src/main/scala/utils/GTimer.scala 25:7]
    end
    if (reset) begin // @[src/main/scala/utils/GTimer.scala 24:20]
      c_1 <= 64'h0; // @[src/main/scala/utils/GTimer.scala 24:20]
    end else begin
      c_1 <= _c_T_3; // @[src/main/scala/utils/GTimer.scala 25:7]
    end
    if (reset) begin // @[src/main/scala/utils/GTimer.scala 24:20]
      c_2 <= 64'h0; // @[src/main/scala/utils/GTimer.scala 24:20]
    end else begin
      c_2 <= _c_T_5; // @[src/main/scala/utils/GTimer.scala 25:7]
    end
    if (reset) begin // @[src/main/scala/utils/GTimer.scala 24:20]
      c_3 <= 64'h0; // @[src/main/scala/utils/GTimer.scala 24:20]
    end else begin
      c_3 <= _c_T_7; // @[src/main/scala/utils/GTimer.scala 25:7]
    end
    if (reset) begin // @[src/main/scala/utils/GTimer.scala 24:20]
      c_4 <= 64'h0; // @[src/main/scala/utils/GTimer.scala 24:20]
    end else begin
      c_4 <= _c_T_9; // @[src/main/scala/utils/GTimer.scala 25:7]
    end
    if (reset) begin // @[src/main/scala/utils/GTimer.scala 24:20]
      c_5 <= 64'h0; // @[src/main/scala/utils/GTimer.scala 24:20]
    end else begin
      c_5 <= _c_T_11; // @[src/main/scala/utils/GTimer.scala 25:7]
    end
    if (reset) begin // @[src/main/scala/utils/GTimer.scala 24:20]
      c_6 <= 64'h0; // @[src/main/scala/utils/GTimer.scala 24:20]
    end else begin
      c_6 <= _c_T_13; // @[src/main/scala/utils/GTimer.scala 25:7]
    end
    if (reset) begin // @[src/main/scala/utils/GTimer.scala 24:20]
      c_7 <= 64'h0; // @[src/main/scala/utils/GTimer.scala 24:20]
    end else begin
      c_7 <= _c_T_15; // @[src/main/scala/utils/GTimer.scala 25:7]
    end
    if (reset) begin // @[src/main/scala/utils/GTimer.scala 24:20]
      c_8 <= 64'h0; // @[src/main/scala/utils/GTimer.scala 24:20]
    end else begin
      c_8 <= _c_T_17; // @[src/main/scala/utils/GTimer.scala 25:7]
    end
    if (reset) begin // @[src/main/scala/utils/GTimer.scala 24:20]
      c_9 <= 64'h0; // @[src/main/scala/utils/GTimer.scala 24:20]
    end else begin
      c_9 <= _c_T_19; // @[src/main/scala/utils/GTimer.scala 25:7]
    end
    if (reset) begin // @[src/main/scala/utils/GTimer.scala 24:20]
      c_10 <= 64'h0; // @[src/main/scala/utils/GTimer.scala 24:20]
    end else begin
      c_10 <= _c_T_21; // @[src/main/scala/utils/GTimer.scala 25:7]
    end
    if (reset) begin // @[src/main/scala/nutcore/mem/Cache.scala 219:33]
      isForwardDataReg <= 1'h0; // @[src/main/scala/nutcore/mem/Cache.scala 219:33]
    end else if (_T_2) begin // @[src/main/scala/nutcore/mem/Cache.scala 221:37]
      isForwardDataReg <= 1'h0; // @[src/main/scala/nutcore/mem/Cache.scala 221:56]
    end else begin
      isForwardDataReg <= _GEN_8;
    end
    if (isForwardData) begin // @[src/main/scala/nutcore/mem/Cache.scala 222:33]
      forwardDataReg_data_data <= io_dataWriteBus_req_bits_data_data; // @[src/main/scala/nutcore/mem/Cache.scala 222:33]
    end
    if (isForwardData) begin // @[src/main/scala/nutcore/mem/Cache.scala 222:33]
      forwardDataReg_waymask <= io_dataWriteBus_req_bits_waymask; // @[src/main/scala/nutcore/mem/Cache.scala 222:33]
    end
    if (reset) begin // @[src/main/scala/utils/GTimer.scala 24:20]
      c_11 <= 64'h0; // @[src/main/scala/utils/GTimer.scala 24:20]
    end else begin
      c_11 <= _c_T_23; // @[src/main/scala/utils/GTimer.scala 25:7]
    end
    if (reset) begin // @[src/main/scala/utils/GTimer.scala 24:20]
      c_12 <= 64'h0; // @[src/main/scala/utils/GTimer.scala 24:20]
    end else begin
      c_12 <= _c_T_25; // @[src/main/scala/utils/GTimer.scala 25:7]
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_13 & DISPLAY_ENABLE & ~reset) begin
          $fwrite(32'h80000002,"[%d] CacheStage2: ",c); // @[src/main/scala/utils/Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_13 & _T_16) begin
          $fwrite(32'h80000002,"[ERROR] metaWay %x metat %x reqt %x\n",metaWay_0_valid,metaWay_0_tag,addr_tag); // @[src/main/scala/utils/Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_13 & DISPLAY_ENABLE & ~reset) begin
          $fwrite(32'h80000002,"[%d] CacheStage2: ",c_1); // @[src/main/scala/utils/Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_13 & _T_16) begin
          $fwrite(32'h80000002,"[ERROR] metaWay %x metat %x reqt %x\n",metaWay_1_valid,metaWay_1_tag,addr_tag); // @[src/main/scala/utils/Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_13 & DISPLAY_ENABLE & ~reset) begin
          $fwrite(32'h80000002,"[%d] CacheStage2: ",c_2); // @[src/main/scala/utils/Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_13 & _T_16) begin
          $fwrite(32'h80000002,"[ERROR] metaWay %x metat %x reqt %x\n",metaWay_2_valid,metaWay_2_tag,addr_tag); // @[src/main/scala/utils/Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_13 & DISPLAY_ENABLE & ~reset) begin
          $fwrite(32'h80000002,"[%d] CacheStage2: ",c_3); // @[src/main/scala/utils/Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_13 & _T_16) begin
          $fwrite(32'h80000002,"[ERROR] metaWay %x metat %x reqt %x\n",metaWay_3_valid,metaWay_3_tag,addr_tag); // @[src/main/scala/utils/Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_13 & DISPLAY_ENABLE & ~reset) begin
          $fwrite(32'h80000002,"[%d] CacheStage2: ",c_4); // @[src/main/scala/utils/Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_13 & _T_16) begin
          $fwrite(32'h80000002,"[ERROR] metaReadResp %x metat %x reqt %x\n",io_metaReadResp_0_valid,
            io_metaReadResp_0_tag,addr_tag); // @[src/main/scala/utils/Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_13 & DISPLAY_ENABLE & ~reset) begin
          $fwrite(32'h80000002,"[%d] CacheStage2: ",c_5); // @[src/main/scala/utils/Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_13 & _T_16) begin
          $fwrite(32'h80000002,"[ERROR] metaReadResp %x metat %x reqt %x\n",io_metaReadResp_1_valid,
            io_metaReadResp_1_tag,addr_tag); // @[src/main/scala/utils/Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_13 & DISPLAY_ENABLE & ~reset) begin
          $fwrite(32'h80000002,"[%d] CacheStage2: ",c_6); // @[src/main/scala/utils/Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_13 & _T_16) begin
          $fwrite(32'h80000002,"[ERROR] metaReadResp %x metat %x reqt %x\n",io_metaReadResp_2_valid,
            io_metaReadResp_2_tag,addr_tag); // @[src/main/scala/utils/Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_13 & DISPLAY_ENABLE & ~reset) begin
          $fwrite(32'h80000002,"[%d] CacheStage2: ",c_7); // @[src/main/scala/utils/Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_13 & _T_16) begin
          $fwrite(32'h80000002,"[ERROR] metaReadResp %x metat %x reqt %x\n",io_metaReadResp_3_valid,
            io_metaReadResp_3_tag,addr_tag); // @[src/main/scala/utils/Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_13 & DISPLAY_ENABLE & ~reset) begin
          $fwrite(32'h80000002,"[%d] CacheStage2: ",c_8); // @[src/main/scala/utils/Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_13 & _T_16) begin
          $fwrite(32'h80000002,"[ERROR] forwardMetaReg isForwardMetaReg %x %x metat %x wm %b\n",isForwardMetaReg,1'h1,
            forwardMetaReg_data_tag,forwardMetaReg_waymask); // @[src/main/scala/utils/Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_13 & DISPLAY_ENABLE & ~reset) begin
          $fwrite(32'h80000002,"[%d] CacheStage2: ",c_9); // @[src/main/scala/utils/Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_13 & _T_16) begin
          $fwrite(32'h80000002,"[ERROR] forwardMeta isForwardMeta %x %x metat %x wm %b\n",isForwardMeta,1'h1,
            io_metaWriteBus_req_bits_data_tag,io_metaWriteBus_req_bits_waymask); // @[src/main/scala/utils/Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_13 & DISPLAY_ENABLE & ~reset) begin
          $fwrite(32'h80000002,"[%d] CacheStage2: ",c_10); // @[src/main/scala/utils/Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_13 & _T_16) begin
          $fwrite(32'h80000002,"[ERROR] hit %b wmask %b hitvec %b\n",io_out_bits_hit,_GEN_6,hitVec); // @[src/main/scala/utils/Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_16 & ~(~(io_in_valid & _T_13))) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Cache.scala:208 assert(!(io.in.valid && PopCount(waymask) > 1.U))\n"); // @[src/main/scala/nutcore/mem/Cache.scala 208:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~(io_in_valid & _T_13)) & _T_16) begin
          $fatal; // @[src/main/scala/nutcore/mem/Cache.scala 208:9]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & ~reset) begin
          $fwrite(32'h80000002,"[%d] CacheStage2: ",c_11); // @[src/main/scala/utils/Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_16) begin
          $fwrite(32'h80000002,"[isFD:%d isFDreg:%d inFire:%d invalid:%d \n",isForwardData,isForwardDataReg,_T,
            io_in_valid); // @[src/main/scala/utils/Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & ~reset) begin
          $fwrite(32'h80000002,"[%d] CacheStage2: ",c_12); // @[src/main/scala/utils/Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_16) begin
          $fwrite(32'h80000002,"[isFM:%d isFMreg:%d metawreq:%x widx:%x ridx:%x \n",isForwardMeta,isForwardMetaReg,
            io_metaWriteBus_req_valid,io_metaWriteBus_req_bits_setIdx,addr_index); // @[src/main/scala/utils/Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  isForwardMetaReg = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  forwardMetaReg_data_tag = _RAND_1[18:0];
  _RAND_2 = {1{`RANDOM}};
  forwardMetaReg_data_dirty = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  forwardMetaReg_waymask = _RAND_3[3:0];
  _RAND_4 = {2{`RANDOM}};
  victimWaymask_lfsr = _RAND_4[63:0];
  _RAND_5 = {2{`RANDOM}};
  c = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  c_1 = _RAND_6[63:0];
  _RAND_7 = {2{`RANDOM}};
  c_2 = _RAND_7[63:0];
  _RAND_8 = {2{`RANDOM}};
  c_3 = _RAND_8[63:0];
  _RAND_9 = {2{`RANDOM}};
  c_4 = _RAND_9[63:0];
  _RAND_10 = {2{`RANDOM}};
  c_5 = _RAND_10[63:0];
  _RAND_11 = {2{`RANDOM}};
  c_6 = _RAND_11[63:0];
  _RAND_12 = {2{`RANDOM}};
  c_7 = _RAND_12[63:0];
  _RAND_13 = {2{`RANDOM}};
  c_8 = _RAND_13[63:0];
  _RAND_14 = {2{`RANDOM}};
  c_9 = _RAND_14[63:0];
  _RAND_15 = {2{`RANDOM}};
  c_10 = _RAND_15[63:0];
  _RAND_16 = {1{`RANDOM}};
  isForwardDataReg = _RAND_16[0:0];
  _RAND_17 = {2{`RANDOM}};
  forwardDataReg_data_data = _RAND_17[63:0];
  _RAND_18 = {1{`RANDOM}};
  forwardDataReg_waymask = _RAND_18[3:0];
  _RAND_19 = {2{`RANDOM}};
  c_11 = _RAND_19[63:0];
  _RAND_20 = {2{`RANDOM}};
  c_12 = _RAND_20[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Arbiter(
  input         io_in_0_valid, // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
  input  [6:0]  io_in_0_bits_setIdx, // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
  input  [18:0] io_in_0_bits_data_tag, // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
  input         io_in_0_bits_data_dirty, // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
  input  [3:0]  io_in_0_bits_waymask, // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
  input         io_in_1_valid, // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
  input  [6:0]  io_in_1_bits_setIdx, // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
  input  [18:0] io_in_1_bits_data_tag, // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
  input         io_in_1_bits_data_dirty, // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
  input  [3:0]  io_in_1_bits_waymask, // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
  output        io_out_valid, // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
  output [6:0]  io_out_bits_setIdx, // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
  output [18:0] io_out_bits_data_tag, // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
  output        io_out_bits_data_dirty, // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
  output [3:0]  io_out_bits_waymask // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
);
  wire  grant_1 = ~io_in_0_valid; // @[src/main/scala/chisel3/util/Arbiter.scala 45:78]
  assign io_out_valid = ~grant_1 | io_in_1_valid; // @[src/main/scala/chisel3/util/Arbiter.scala 148:31]
  assign io_out_bits_setIdx = io_in_0_valid ? io_in_0_bits_setIdx : io_in_1_bits_setIdx; // @[src/main/scala/chisel3/util/Arbiter.scala 137:15 139:26 141:19]
  assign io_out_bits_data_tag = io_in_0_valid ? io_in_0_bits_data_tag : io_in_1_bits_data_tag; // @[src/main/scala/chisel3/util/Arbiter.scala 137:15 139:26 141:19]
  assign io_out_bits_data_dirty = io_in_0_valid ? io_in_0_bits_data_dirty : io_in_1_bits_data_dirty; // @[src/main/scala/chisel3/util/Arbiter.scala 137:15 139:26 141:19]
  assign io_out_bits_waymask = io_in_0_valid ? io_in_0_bits_waymask : io_in_1_bits_waymask; // @[src/main/scala/chisel3/util/Arbiter.scala 137:15 139:26 141:19]
endmodule
module Arbiter_1(
  input         io_in_0_valid, // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
  input  [9:0]  io_in_0_bits_setIdx, // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
  input  [63:0] io_in_0_bits_data_data, // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
  input  [3:0]  io_in_0_bits_waymask, // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
  input         io_in_1_valid, // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
  input  [9:0]  io_in_1_bits_setIdx, // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
  input  [63:0] io_in_1_bits_data_data, // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
  input  [3:0]  io_in_1_bits_waymask, // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
  output        io_out_valid, // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
  output [9:0]  io_out_bits_setIdx, // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
  output [63:0] io_out_bits_data_data, // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
  output [3:0]  io_out_bits_waymask // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
);
  wire  grant_1 = ~io_in_0_valid; // @[src/main/scala/chisel3/util/Arbiter.scala 45:78]
  assign io_out_valid = ~grant_1 | io_in_1_valid; // @[src/main/scala/chisel3/util/Arbiter.scala 148:31]
  assign io_out_bits_setIdx = io_in_0_valid ? io_in_0_bits_setIdx : io_in_1_bits_setIdx; // @[src/main/scala/chisel3/util/Arbiter.scala 137:15 139:26 141:19]
  assign io_out_bits_data_data = io_in_0_valid ? io_in_0_bits_data_data : io_in_1_bits_data_data; // @[src/main/scala/chisel3/util/Arbiter.scala 137:15 139:26 141:19]
  assign io_out_bits_waymask = io_in_0_valid ? io_in_0_bits_waymask : io_in_1_bits_waymask; // @[src/main/scala/chisel3/util/Arbiter.scala 137:15 139:26 141:19]
endmodule
module CacheStage3(
  input         clock,
  input         reset,
  output        io_in_ready, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  input         io_in_valid, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  input  [31:0] io_in_bits_req_addr, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  input  [2:0]  io_in_bits_req_size, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  input  [3:0]  io_in_bits_req_cmd, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  input  [7:0]  io_in_bits_req_wmask, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  input  [63:0] io_in_bits_req_wdata, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  input  [86:0] io_in_bits_req_user, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  input  [18:0] io_in_bits_metas_0_tag, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  input         io_in_bits_metas_0_valid, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  input         io_in_bits_metas_0_dirty, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  input  [18:0] io_in_bits_metas_1_tag, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  input         io_in_bits_metas_1_valid, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  input         io_in_bits_metas_1_dirty, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  input  [18:0] io_in_bits_metas_2_tag, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  input         io_in_bits_metas_2_valid, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  input         io_in_bits_metas_2_dirty, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  input  [18:0] io_in_bits_metas_3_tag, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  input         io_in_bits_metas_3_valid, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  input         io_in_bits_metas_3_dirty, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  input  [63:0] io_in_bits_datas_0_data, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  input  [63:0] io_in_bits_datas_1_data, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  input  [63:0] io_in_bits_datas_2_data, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  input  [63:0] io_in_bits_datas_3_data, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  input         io_in_bits_hit, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  input  [3:0]  io_in_bits_waymask, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  input         io_in_bits_mmio, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  input         io_in_bits_isForwardData, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  input  [63:0] io_in_bits_forwardData_data_data, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  input  [3:0]  io_in_bits_forwardData_waymask, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  input         io_out_ready, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  output        io_out_valid, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  output [3:0]  io_out_bits_cmd, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  output [63:0] io_out_bits_rdata, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  output [86:0] io_out_bits_user, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  output        io_isFinish, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  input         io_flush, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  input         io_dataReadBus_req_ready, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  output        io_dataReadBus_req_valid, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  output [9:0]  io_dataReadBus_req_bits_setIdx, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  input  [63:0] io_dataReadBus_resp_data_0_data, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  input  [63:0] io_dataReadBus_resp_data_1_data, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  input  [63:0] io_dataReadBus_resp_data_2_data, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  input  [63:0] io_dataReadBus_resp_data_3_data, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  output        io_dataWriteBus_req_valid, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  output [9:0]  io_dataWriteBus_req_bits_setIdx, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  output [63:0] io_dataWriteBus_req_bits_data_data, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  output [3:0]  io_dataWriteBus_req_bits_waymask, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  output        io_metaWriteBus_req_valid, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  output [6:0]  io_metaWriteBus_req_bits_setIdx, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  output [18:0] io_metaWriteBus_req_bits_data_tag, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  output        io_metaWriteBus_req_bits_data_valid, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  output        io_metaWriteBus_req_bits_data_dirty, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  output [3:0]  io_metaWriteBus_req_bits_waymask, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  input         io_mem_req_ready, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  output        io_mem_req_valid, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  output [31:0] io_mem_req_bits_addr, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  output [2:0]  io_mem_req_bits_size, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  output [3:0]  io_mem_req_bits_cmd, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  output [7:0]  io_mem_req_bits_wmask, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  output [63:0] io_mem_req_bits_wdata, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  output        io_mem_resp_ready, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  input         io_mem_resp_valid, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  input  [3:0]  io_mem_resp_bits_cmd, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  input  [63:0] io_mem_resp_bits_rdata, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  input         io_mmio_req_ready, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  output        io_mmio_req_valid, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  output [31:0] io_mmio_req_bits_addr, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  output        io_mmio_resp_ready, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  input         io_mmio_resp_valid, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  input  [63:0] io_mmio_resp_bits_rdata, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  output        io_cohResp_valid, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  input         DISPLAY_ENABLE
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [63:0] _RAND_12;
  reg [63:0] _RAND_13;
  reg [63:0] _RAND_14;
  reg [63:0] _RAND_15;
  reg [63:0] _RAND_16;
  reg [63:0] _RAND_17;
  reg [63:0] _RAND_18;
  reg [63:0] _RAND_19;
  reg [63:0] _RAND_20;
  reg [63:0] _RAND_21;
  reg [63:0] _RAND_22;
  reg [63:0] _RAND_23;
`endif // RANDOMIZE_REG_INIT
  wire  metaWriteArb_io_in_0_valid; // @[src/main/scala/nutcore/mem/Cache.scala 254:28]
  wire [6:0] metaWriteArb_io_in_0_bits_setIdx; // @[src/main/scala/nutcore/mem/Cache.scala 254:28]
  wire [18:0] metaWriteArb_io_in_0_bits_data_tag; // @[src/main/scala/nutcore/mem/Cache.scala 254:28]
  wire  metaWriteArb_io_in_0_bits_data_dirty; // @[src/main/scala/nutcore/mem/Cache.scala 254:28]
  wire [3:0] metaWriteArb_io_in_0_bits_waymask; // @[src/main/scala/nutcore/mem/Cache.scala 254:28]
  wire  metaWriteArb_io_in_1_valid; // @[src/main/scala/nutcore/mem/Cache.scala 254:28]
  wire [6:0] metaWriteArb_io_in_1_bits_setIdx; // @[src/main/scala/nutcore/mem/Cache.scala 254:28]
  wire [18:0] metaWriteArb_io_in_1_bits_data_tag; // @[src/main/scala/nutcore/mem/Cache.scala 254:28]
  wire  metaWriteArb_io_in_1_bits_data_dirty; // @[src/main/scala/nutcore/mem/Cache.scala 254:28]
  wire [3:0] metaWriteArb_io_in_1_bits_waymask; // @[src/main/scala/nutcore/mem/Cache.scala 254:28]
  wire  metaWriteArb_io_out_valid; // @[src/main/scala/nutcore/mem/Cache.scala 254:28]
  wire [6:0] metaWriteArb_io_out_bits_setIdx; // @[src/main/scala/nutcore/mem/Cache.scala 254:28]
  wire [18:0] metaWriteArb_io_out_bits_data_tag; // @[src/main/scala/nutcore/mem/Cache.scala 254:28]
  wire  metaWriteArb_io_out_bits_data_dirty; // @[src/main/scala/nutcore/mem/Cache.scala 254:28]
  wire [3:0] metaWriteArb_io_out_bits_waymask; // @[src/main/scala/nutcore/mem/Cache.scala 254:28]
  wire  dataWriteArb_io_in_0_valid; // @[src/main/scala/nutcore/mem/Cache.scala 255:28]
  wire [9:0] dataWriteArb_io_in_0_bits_setIdx; // @[src/main/scala/nutcore/mem/Cache.scala 255:28]
  wire [63:0] dataWriteArb_io_in_0_bits_data_data; // @[src/main/scala/nutcore/mem/Cache.scala 255:28]
  wire [3:0] dataWriteArb_io_in_0_bits_waymask; // @[src/main/scala/nutcore/mem/Cache.scala 255:28]
  wire  dataWriteArb_io_in_1_valid; // @[src/main/scala/nutcore/mem/Cache.scala 255:28]
  wire [9:0] dataWriteArb_io_in_1_bits_setIdx; // @[src/main/scala/nutcore/mem/Cache.scala 255:28]
  wire [63:0] dataWriteArb_io_in_1_bits_data_data; // @[src/main/scala/nutcore/mem/Cache.scala 255:28]
  wire [3:0] dataWriteArb_io_in_1_bits_waymask; // @[src/main/scala/nutcore/mem/Cache.scala 255:28]
  wire  dataWriteArb_io_out_valid; // @[src/main/scala/nutcore/mem/Cache.scala 255:28]
  wire [9:0] dataWriteArb_io_out_bits_setIdx; // @[src/main/scala/nutcore/mem/Cache.scala 255:28]
  wire [63:0] dataWriteArb_io_out_bits_data_data; // @[src/main/scala/nutcore/mem/Cache.scala 255:28]
  wire [3:0] dataWriteArb_io_out_bits_waymask; // @[src/main/scala/nutcore/mem/Cache.scala 255:28]
  wire [2:0] addr_wordIndex = io_in_bits_req_addr[5:3]; // @[src/main/scala/nutcore/mem/Cache.scala 258:31]
  wire [6:0] addr_index = io_in_bits_req_addr[12:6]; // @[src/main/scala/nutcore/mem/Cache.scala 258:31]
  wire [18:0] addr_tag = io_in_bits_req_addr[31:13]; // @[src/main/scala/nutcore/mem/Cache.scala 258:31]
  wire  mmio = io_in_valid & io_in_bits_mmio; // @[src/main/scala/nutcore/mem/Cache.scala 259:26]
  wire  hit = io_in_valid & io_in_bits_hit; // @[src/main/scala/nutcore/mem/Cache.scala 260:25]
  wire  miss = io_in_valid & ~io_in_bits_hit; // @[src/main/scala/nutcore/mem/Cache.scala 261:26]
  wire [18:0] _meta_T_18 = io_in_bits_waymask[0] ? io_in_bits_metas_0_tag : 19'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [18:0] _meta_T_19 = io_in_bits_waymask[1] ? io_in_bits_metas_1_tag : 19'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [18:0] _meta_T_20 = io_in_bits_waymask[2] ? io_in_bits_metas_2_tag : 19'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [18:0] _meta_T_21 = io_in_bits_waymask[3] ? io_in_bits_metas_3_tag : 19'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [18:0] _meta_T_22 = _meta_T_18 | _meta_T_19; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [18:0] _meta_T_23 = _meta_T_22 | _meta_T_20; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [18:0] meta_tag = _meta_T_23 | _meta_T_21; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _T_3 = ~reset; // @[src/main/scala/nutcore/mem/Cache.scala 265:9]
  wire  useForwardData = io_in_bits_isForwardData & io_in_bits_waymask == io_in_bits_forwardData_waymask; // @[src/main/scala/nutcore/mem/Cache.scala 273:49]
  wire [63:0] _dataReadArray_T_4 = io_in_bits_waymask[0] ? io_in_bits_datas_0_data : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _dataReadArray_T_5 = io_in_bits_waymask[1] ? io_in_bits_datas_1_data : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _dataReadArray_T_6 = io_in_bits_waymask[2] ? io_in_bits_datas_2_data : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _dataReadArray_T_7 = io_in_bits_waymask[3] ? io_in_bits_datas_3_data : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _dataReadArray_T_8 = _dataReadArray_T_4 | _dataReadArray_T_5; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _dataReadArray_T_9 = _dataReadArray_T_8 | _dataReadArray_T_6; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _dataReadArray_T_10 = _dataReadArray_T_9 | _dataReadArray_T_7; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] dataRead = useForwardData ? io_in_bits_forwardData_data_data : _dataReadArray_T_10; // @[src/main/scala/nutcore/mem/Cache.scala 275:21]
  wire  _T_5 = io_out_ready & io_out_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  wire [9:0] dataHitWriteBus_x3 = {addr_index,addr_wordIndex}; // @[src/main/scala/nutcore/mem/Cache.scala 286:35]
  reg [3:0] state; // @[src/main/scala/nutcore/mem/Cache.scala 294:22]
  reg  needFlush; // @[src/main/scala/nutcore/mem/Cache.scala 295:26]
  wire  _GEN_1 = io_flush & state != 4'h0 | needFlush; // @[src/main/scala/nutcore/mem/Cache.scala 295:26 297:{41,53}]
  reg [2:0] readBeatCnt_value; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
  reg [2:0] writeBeatCnt_value; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
  reg [1:0] state2; // @[src/main/scala/nutcore/mem/Cache.scala 304:23]
  wire  _T_14 = state == 4'h3; // @[src/main/scala/nutcore/mem/Cache.scala 306:39]
  wire  _T_15 = state == 4'h8; // @[src/main/scala/nutcore/mem/Cache.scala 306:66]
  wire [2:0] _T_20 = _T_15 ? readBeatCnt_value : writeBeatCnt_value; // @[src/main/scala/nutcore/mem/Cache.scala 307:33]
  reg [63:0] dataWay_0_data; // @[src/main/scala/nutcore/mem/Cache.scala 308:26]
  reg [63:0] dataWay_1_data; // @[src/main/scala/nutcore/mem/Cache.scala 308:26]
  reg [63:0] dataWay_2_data; // @[src/main/scala/nutcore/mem/Cache.scala 308:26]
  reg [63:0] dataWay_3_data; // @[src/main/scala/nutcore/mem/Cache.scala 308:26]
  wire [63:0] _dataHitWay_T_4 = io_in_bits_waymask[0] ? dataWay_0_data : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _dataHitWay_T_5 = io_in_bits_waymask[1] ? dataWay_1_data : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _dataHitWay_T_6 = io_in_bits_waymask[2] ? dataWay_2_data : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _dataHitWay_T_7 = io_in_bits_waymask[3] ? dataWay_3_data : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _dataHitWay_T_8 = _dataHitWay_T_4 | _dataHitWay_T_5; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _dataHitWay_T_9 = _dataHitWay_T_8 | _dataHitWay_T_6; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _T_23 = io_dataReadBus_req_ready & io_dataReadBus_req_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  wire  _T_26 = io_mem_req_ready & io_mem_req_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  wire [1:0] _GEN_8 = _T_26 | io_cohResp_valid ? 2'h0 : state2; // @[src/main/scala/nutcore/mem/Cache.scala 314:105 304:23 314:96]
  wire [31:0] raddr = {io_in_bits_req_addr[31:3],3'h0}; // @[src/main/scala/nutcore/mem/Cache.scala 318:35]
  wire [31:0] waddr = {meta_tag,addr_index,6'h0}; // @[src/main/scala/nutcore/mem/Cache.scala 321:18]
  wire  _cmd_T = state == 4'h1; // @[src/main/scala/nutcore/mem/Cache.scala 322:23]
  wire [2:0] _cmd_T_2 = writeBeatCnt_value == 3'h7 ? 3'h7 : 3'h3; // @[src/main/scala/nutcore/mem/Cache.scala 323:8]
  wire [2:0] cmd = state == 4'h1 ? 3'h2 : _cmd_T_2; // @[src/main/scala/nutcore/mem/Cache.scala 322:16]
  wire  _io_mem_req_valid_T_2 = state2 == 2'h2; // @[src/main/scala/nutcore/mem/Cache.scala 329:89]
  reg  afterFirstRead; // @[src/main/scala/nutcore/mem/Cache.scala 336:31]
  reg  alreadyOutFire; // @[src/main/scala/nutcore/mem/Cache.scala 337:33]
  wire  _GEN_12 = _T_5 | alreadyOutFire; // @[src/main/scala/nutcore/mem/Cache.scala 337:{33,33,33}]
  wire  _readingFirst_T_1 = io_mem_resp_ready & io_mem_resp_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  wire  _readingFirst_T_3 = state == 4'h2; // @[src/main/scala/nutcore/mem/Cache.scala 338:68]
  wire  readingFirst = ~afterFirstRead & _readingFirst_T_1 & state == 4'h2; // @[src/main/scala/nutcore/mem/Cache.scala 338:58]
  wire  _inRdataRegDemand_T_2 = mmio ? state == 4'h6 : readingFirst; // @[src/main/scala/nutcore/mem/Cache.scala 340:39]
  reg [63:0] inRdataRegDemand; // @[src/main/scala/nutcore/mem/Cache.scala 339:35]
  wire  _io_cohResp_valid_T = state == 4'h0; // @[src/main/scala/nutcore/mem/Cache.scala 343:31]
  wire  _T_41 = io_mmio_req_ready & io_mmio_req_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  wire  _T_43 = io_mmio_resp_ready & io_mmio_resp_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  wire [3:0] _GEN_26 = _T_43 ? 4'h7 : state; // @[src/main/scala/nutcore/mem/Cache.scala 294:22 372:{48,56}]
  wire [2:0] _value_T_7 = readBeatCnt_value + 3'h1; // @[src/main/scala/chisel3/util/Counter.scala 77:24]
  wire [2:0] _GEN_27 = io_cohResp_valid ? _value_T_7 : readBeatCnt_value; // @[src/main/scala/nutcore/mem/Cache.scala 375:46 src/main/scala/chisel3/util/Counter.scala 77:15 61:40]
  wire [3:0] _GEN_29 = _T_26 ? 4'h2 : state; // @[src/main/scala/nutcore/mem/Cache.scala 379:48 380:13 294:22]
  wire [2:0] _GEN_30 = _T_26 ? addr_wordIndex : readBeatCnt_value; // @[src/main/scala/nutcore/mem/Cache.scala 379:48 381:25 src/main/scala/chisel3/util/Counter.scala 61:40]
  wire  _T_57 = io_mem_resp_bits_cmd == 4'h6; // @[src/main/scala/bus/simplebus/SimpleBus.scala 91:24]
  wire [3:0] _GEN_32 = _T_57 ? 4'h7 : state; // @[src/main/scala/nutcore/mem/Cache.scala 294:22 389:{44,52}]
  wire  _GEN_33 = _readingFirst_T_1 | afterFirstRead; // @[src/main/scala/nutcore/mem/Cache.scala 385:31 386:24 336:31]
  wire [2:0] _GEN_34 = _readingFirst_T_1 ? _value_T_7 : readBeatCnt_value; // @[src/main/scala/nutcore/mem/Cache.scala 385:31 src/main/scala/chisel3/util/Counter.scala 77:15 61:40]
  wire [3:0] _GEN_36 = _readingFirst_T_1 ? _GEN_32 : state; // @[src/main/scala/nutcore/mem/Cache.scala 294:22 385:31]
  wire [2:0] _value_T_11 = writeBeatCnt_value + 3'h1; // @[src/main/scala/chisel3/util/Counter.scala 77:24]
  wire [2:0] _GEN_37 = _T_26 ? _value_T_11 : writeBeatCnt_value; // @[src/main/scala/nutcore/mem/Cache.scala 394:30 src/main/scala/chisel3/util/Counter.scala 77:15 61:40]
  wire  _T_60 = io_mem_req_bits_cmd == 4'h7; // @[src/main/scala/bus/simplebus/SimpleBus.scala 78:27]
  wire [3:0] _GEN_38 = _T_60 & _T_26 ? 4'h4 : state; // @[src/main/scala/nutcore/mem/Cache.scala 294:22 395:{63,71}]
  wire [3:0] _GEN_39 = _readingFirst_T_1 ? 4'h1 : state; // @[src/main/scala/nutcore/mem/Cache.scala 294:22 398:{51,59}]
  wire [3:0] _GEN_40 = _T_5 | needFlush | alreadyOutFire ? 4'h0 : state; // @[src/main/scala/nutcore/mem/Cache.scala 294:22 399:{74,82}]
  wire [3:0] _GEN_41 = 4'h7 == state ? _GEN_40 : state; // @[src/main/scala/nutcore/mem/Cache.scala 353:18 294:22]
  wire [3:0] _GEN_42 = 4'h4 == state ? _GEN_39 : _GEN_41; // @[src/main/scala/nutcore/mem/Cache.scala 353:18]
  wire [2:0] _GEN_43 = 4'h3 == state ? _GEN_37 : writeBeatCnt_value; // @[src/main/scala/nutcore/mem/Cache.scala 353:18 src/main/scala/chisel3/util/Counter.scala 61:40]
  wire [3:0] _GEN_44 = 4'h3 == state ? _GEN_38 : _GEN_42; // @[src/main/scala/nutcore/mem/Cache.scala 353:18]
  wire  _GEN_45 = 4'h2 == state ? _GEN_33 : afterFirstRead; // @[src/main/scala/nutcore/mem/Cache.scala 353:18 336:31]
  wire [2:0] _GEN_46 = 4'h2 == state ? _GEN_34 : readBeatCnt_value; // @[src/main/scala/nutcore/mem/Cache.scala 353:18 src/main/scala/chisel3/util/Counter.scala 61:40]
  wire [3:0] _GEN_48 = 4'h2 == state ? _GEN_36 : _GEN_44; // @[src/main/scala/nutcore/mem/Cache.scala 353:18]
  wire [2:0] _GEN_49 = 4'h2 == state ? writeBeatCnt_value : _GEN_43; // @[src/main/scala/nutcore/mem/Cache.scala 353:18 src/main/scala/chisel3/util/Counter.scala 61:40]
  wire [3:0] _GEN_50 = 4'h1 == state ? _GEN_29 : _GEN_48; // @[src/main/scala/nutcore/mem/Cache.scala 353:18]
  wire [2:0] _GEN_51 = 4'h1 == state ? _GEN_30 : _GEN_46; // @[src/main/scala/nutcore/mem/Cache.scala 353:18]
  wire  _GEN_52 = 4'h1 == state ? afterFirstRead : _GEN_45; // @[src/main/scala/nutcore/mem/Cache.scala 353:18 336:31]
  wire [2:0] _GEN_54 = 4'h1 == state ? writeBeatCnt_value : _GEN_49; // @[src/main/scala/nutcore/mem/Cache.scala 353:18 src/main/scala/chisel3/util/Counter.scala 61:40]
  wire [2:0] _GEN_55 = 4'h8 == state ? _GEN_27 : _GEN_51; // @[src/main/scala/nutcore/mem/Cache.scala 353:18]
  wire [3:0] _GEN_56 = 4'h8 == state ? state : _GEN_50; // @[src/main/scala/nutcore/mem/Cache.scala 353:18]
  wire  _GEN_57 = 4'h8 == state ? afterFirstRead : _GEN_52; // @[src/main/scala/nutcore/mem/Cache.scala 353:18 336:31]
  wire [2:0] _GEN_59 = 4'h8 == state ? writeBeatCnt_value : _GEN_54; // @[src/main/scala/nutcore/mem/Cache.scala 353:18 src/main/scala/chisel3/util/Counter.scala 61:40]
  wire  dataRefillWriteBus_x9 = _readingFirst_T_3 & _readingFirst_T_1; // @[src/main/scala/nutcore/mem/Cache.scala 404:39]
  wire  _io_out_valid_T_4 = state == 4'h7; // @[src/main/scala/nutcore/mem/Cache.scala 446:48]
  wire  _io_out_valid_T_23 = mmio ? _io_out_valid_T_4 : afterFirstRead & ~alreadyOutFire; // @[src/main/scala/nutcore/mem/Cache.scala 447:45]
  wire  _io_out_valid_T_24 = hit | _io_out_valid_T_23; // @[src/main/scala/nutcore/mem/Cache.scala 447:28]
  wire [255:0] _T_89 = {io_in_bits_datas_3_data,io_in_bits_datas_2_data,io_in_bits_datas_1_data,io_in_bits_datas_0_data}
    ; // @[src/main/scala/nutcore/mem/Cache.scala 464:465]
  reg [63:0] c; // @[src/main/scala/utils/GTimer.scala 24:20]
  wire [63:0] _c_T_1 = c + 64'h1; // @[src/main/scala/utils/GTimer.scala 25:12]
  reg [63:0] c_1; // @[src/main/scala/utils/GTimer.scala 24:20]
  wire [63:0] _c_T_3 = c_1 + 64'h1; // @[src/main/scala/utils/GTimer.scala 25:12]
  reg [63:0] c_2; // @[src/main/scala/utils/GTimer.scala 24:20]
  wire [63:0] _c_T_5 = c_2 + 64'h1; // @[src/main/scala/utils/GTimer.scala 25:12]
  wire  _T_96 = io_metaWriteBus_req_valid & DISPLAY_ENABLE; // @[src/main/scala/utils/Debug.scala 55:16]
  reg [63:0] c_3; // @[src/main/scala/utils/GTimer.scala 24:20]
  wire [63:0] _c_T_7 = c_3 + 64'h1; // @[src/main/scala/utils/GTimer.scala 25:12]
  reg [63:0] c_4; // @[src/main/scala/utils/GTimer.scala 24:20]
  wire [63:0] _c_T_9 = c_4 + 64'h1; // @[src/main/scala/utils/GTimer.scala 25:12]
  reg [63:0] c_5; // @[src/main/scala/utils/GTimer.scala 24:20]
  wire [63:0] _c_T_11 = c_5 + 64'h1; // @[src/main/scala/utils/GTimer.scala 25:12]
  reg [63:0] c_6; // @[src/main/scala/utils/GTimer.scala 24:20]
  wire [63:0] _c_T_13 = c_6 + 64'h1; // @[src/main/scala/utils/GTimer.scala 25:12]
  reg [63:0] c_7; // @[src/main/scala/utils/GTimer.scala 24:20]
  wire [63:0] _c_T_15 = c_7 + 64'h1; // @[src/main/scala/utils/GTimer.scala 25:12]
  reg [63:0] c_8; // @[src/main/scala/utils/GTimer.scala 24:20]
  wire [63:0] _c_T_17 = c_8 + 64'h1; // @[src/main/scala/utils/GTimer.scala 25:12]
  wire  _T_128 = io_dataWriteBus_req_valid & DISPLAY_ENABLE; // @[src/main/scala/utils/Debug.scala 55:16]
  wire  _T_135 = _T_14 & _T_26; // @[src/main/scala/nutcore/mem/Cache.scala 473:35]
  reg [63:0] c_9; // @[src/main/scala/utils/GTimer.scala 24:20]
  wire [63:0] _c_T_19 = c_9 + 64'h1; // @[src/main/scala/utils/GTimer.scala 25:12]
  wire  _T_140 = _T_135 & DISPLAY_ENABLE; // @[src/main/scala/utils/Debug.scala 55:16]
  wire  _T_147 = _cmd_T & _T_26; // @[src/main/scala/nutcore/mem/Cache.scala 474:34]
  reg [63:0] c_10; // @[src/main/scala/utils/GTimer.scala 24:20]
  wire [63:0] _c_T_21 = c_10 + 64'h1; // @[src/main/scala/utils/GTimer.scala 25:12]
  wire  _T_152 = _T_147 & DISPLAY_ENABLE; // @[src/main/scala/utils/Debug.scala 55:16]
  reg [63:0] c_11; // @[src/main/scala/utils/GTimer.scala 24:20]
  wire [63:0] _c_T_23 = c_11 + 64'h1; // @[src/main/scala/utils/GTimer.scala 25:12]
  wire  _T_164 = dataRefillWriteBus_x9 & DISPLAY_ENABLE; // @[src/main/scala/utils/Debug.scala 55:16]
  Arbiter metaWriteArb ( // @[src/main/scala/nutcore/mem/Cache.scala 254:28]
    .io_in_0_valid(metaWriteArb_io_in_0_valid),
    .io_in_0_bits_setIdx(metaWriteArb_io_in_0_bits_setIdx),
    .io_in_0_bits_data_tag(metaWriteArb_io_in_0_bits_data_tag),
    .io_in_0_bits_data_dirty(metaWriteArb_io_in_0_bits_data_dirty),
    .io_in_0_bits_waymask(metaWriteArb_io_in_0_bits_waymask),
    .io_in_1_valid(metaWriteArb_io_in_1_valid),
    .io_in_1_bits_setIdx(metaWriteArb_io_in_1_bits_setIdx),
    .io_in_1_bits_data_tag(metaWriteArb_io_in_1_bits_data_tag),
    .io_in_1_bits_data_dirty(metaWriteArb_io_in_1_bits_data_dirty),
    .io_in_1_bits_waymask(metaWriteArb_io_in_1_bits_waymask),
    .io_out_valid(metaWriteArb_io_out_valid),
    .io_out_bits_setIdx(metaWriteArb_io_out_bits_setIdx),
    .io_out_bits_data_tag(metaWriteArb_io_out_bits_data_tag),
    .io_out_bits_data_dirty(metaWriteArb_io_out_bits_data_dirty),
    .io_out_bits_waymask(metaWriteArb_io_out_bits_waymask)
  );
  Arbiter_1 dataWriteArb ( // @[src/main/scala/nutcore/mem/Cache.scala 255:28]
    .io_in_0_valid(dataWriteArb_io_in_0_valid),
    .io_in_0_bits_setIdx(dataWriteArb_io_in_0_bits_setIdx),
    .io_in_0_bits_data_data(dataWriteArb_io_in_0_bits_data_data),
    .io_in_0_bits_waymask(dataWriteArb_io_in_0_bits_waymask),
    .io_in_1_valid(dataWriteArb_io_in_1_valid),
    .io_in_1_bits_setIdx(dataWriteArb_io_in_1_bits_setIdx),
    .io_in_1_bits_data_data(dataWriteArb_io_in_1_bits_data_data),
    .io_in_1_bits_waymask(dataWriteArb_io_in_1_bits_waymask),
    .io_out_valid(dataWriteArb_io_out_valid),
    .io_out_bits_setIdx(dataWriteArb_io_out_bits_setIdx),
    .io_out_bits_data_data(dataWriteArb_io_out_bits_data_data),
    .io_out_bits_waymask(dataWriteArb_io_out_bits_waymask)
  );
  assign io_in_ready = io_out_ready & _io_cohResp_valid_T & ~miss; // @[src/main/scala/nutcore/mem/Cache.scala 458:70]
  assign io_out_valid = io_in_valid & _io_out_valid_T_24; // @[src/main/scala/nutcore/mem/Cache.scala 445:31]
  assign io_out_bits_cmd = 4'h6; // @[src/main/scala/nutcore/mem/Cache.scala 440:21]
  assign io_out_bits_rdata = hit ? dataRead : inRdataRegDemand; // @[src/main/scala/nutcore/mem/Cache.scala 439:29]
  assign io_out_bits_user = io_in_bits_req_user; // @[src/main/scala/nutcore/mem/Cache.scala 442:56]
  assign io_isFinish = hit ? _T_5 : _io_out_valid_T_4 & _GEN_12; // @[src/main/scala/nutcore/mem/Cache.scala 455:8]
  assign io_dataReadBus_req_valid = (state == 4'h3 | state == 4'h8) & state2 == 2'h0; // @[src/main/scala/nutcore/mem/Cache.scala 306:81]
  assign io_dataReadBus_req_bits_setIdx = {addr_index,_T_20}; // @[src/main/scala/nutcore/mem/Cache.scala 307:17]
  assign io_dataWriteBus_req_valid = dataWriteArb_io_out_valid; // @[src/main/scala/nutcore/mem/Cache.scala 409:23]
  assign io_dataWriteBus_req_bits_setIdx = dataWriteArb_io_out_bits_setIdx; // @[src/main/scala/nutcore/mem/Cache.scala 409:23]
  assign io_dataWriteBus_req_bits_data_data = dataWriteArb_io_out_bits_data_data; // @[src/main/scala/nutcore/mem/Cache.scala 409:23]
  assign io_dataWriteBus_req_bits_waymask = dataWriteArb_io_out_bits_waymask; // @[src/main/scala/nutcore/mem/Cache.scala 409:23]
  assign io_metaWriteBus_req_valid = metaWriteArb_io_out_valid; // @[src/main/scala/nutcore/mem/Cache.scala 419:23]
  assign io_metaWriteBus_req_bits_setIdx = metaWriteArb_io_out_bits_setIdx; // @[src/main/scala/nutcore/mem/Cache.scala 419:23]
  assign io_metaWriteBus_req_bits_data_tag = metaWriteArb_io_out_bits_data_tag; // @[src/main/scala/nutcore/mem/Cache.scala 419:23]
  assign io_metaWriteBus_req_bits_data_valid = 1'h1; // @[src/main/scala/nutcore/mem/Cache.scala 419:23]
  assign io_metaWriteBus_req_bits_data_dirty = metaWriteArb_io_out_bits_data_dirty; // @[src/main/scala/nutcore/mem/Cache.scala 419:23]
  assign io_metaWriteBus_req_bits_waymask = metaWriteArb_io_out_bits_waymask; // @[src/main/scala/nutcore/mem/Cache.scala 419:23]
  assign io_mem_req_valid = _cmd_T | _T_14 & state2 == 2'h2; // @[src/main/scala/nutcore/mem/Cache.scala 329:48]
  assign io_mem_req_bits_addr = _cmd_T ? raddr : waddr; // @[src/main/scala/nutcore/mem/Cache.scala 324:35]
  assign io_mem_req_bits_size = 3'h3; // @[src/main/scala/bus/simplebus/SimpleBus.scala 66:15]
  assign io_mem_req_bits_cmd = {{1'd0}, cmd}; // @[src/main/scala/bus/simplebus/SimpleBus.scala 65:14]
  assign io_mem_req_bits_wmask = 8'hff; // @[src/main/scala/nutcore/mem/Cache.scala 326:37]
  assign io_mem_req_bits_wdata = _dataHitWay_T_9 | _dataHitWay_T_7; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign io_mem_resp_ready = 1'h1; // @[src/main/scala/nutcore/mem/Cache.scala 328:21]
  assign io_mmio_req_valid = state == 4'h5; // @[src/main/scala/nutcore/mem/Cache.scala 334:31]
  assign io_mmio_req_bits_addr = io_in_bits_req_addr; // @[src/main/scala/nutcore/mem/Cache.scala 332:20]
  assign io_mmio_resp_ready = 1'h1; // @[src/main/scala/nutcore/mem/Cache.scala 333:22]
  assign io_cohResp_valid = _T_15 & _io_mem_req_valid_T_2; // @[src/main/scala/nutcore/mem/Cache.scala 344:46]
  assign metaWriteArb_io_in_0_valid = 1'h0; // @[src/main/scala/nutcore/mem/Cache.scala 289:22]
  assign metaWriteArb_io_in_0_bits_setIdx = io_in_bits_req_addr[12:6]; // @[src/main/scala/nutcore/mem/Cache.scala 77:45]
  assign metaWriteArb_io_in_0_bits_data_tag = _meta_T_23 | _meta_T_21; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign metaWriteArb_io_in_0_bits_data_dirty = 1'h0; // @[src/main/scala/nutcore/mem/Cache.scala 290:16 95:16]
  assign metaWriteArb_io_in_0_bits_waymask = io_in_bits_waymask; // @[src/main/scala/nutcore/mem/Cache.scala 288:29 src/main/scala/utils/SRAMTemplate.scala 38:24]
  assign metaWriteArb_io_in_1_valid = dataRefillWriteBus_x9 & _T_57; // @[src/main/scala/nutcore/mem/Cache.scala 412:59]
  assign metaWriteArb_io_in_1_bits_setIdx = io_in_bits_req_addr[12:6]; // @[src/main/scala/nutcore/mem/Cache.scala 77:45]
  assign metaWriteArb_io_in_1_bits_data_tag = io_in_bits_req_addr[31:13]; // @[src/main/scala/nutcore/mem/Cache.scala 258:31]
  assign metaWriteArb_io_in_1_bits_data_dirty = 1'h0; // @[src/main/scala/nutcore/mem/Cache.scala 413:85]
  assign metaWriteArb_io_in_1_bits_waymask = io_in_bits_waymask; // @[src/main/scala/nutcore/mem/Cache.scala 411:32 src/main/scala/utils/SRAMTemplate.scala 38:24]
  assign dataWriteArb_io_in_0_valid = 1'h0; // @[src/main/scala/nutcore/mem/Cache.scala 283:22]
  assign dataWriteArb_io_in_0_bits_setIdx = {addr_index,addr_wordIndex}; // @[src/main/scala/nutcore/mem/Cache.scala 286:35]
  assign dataWriteArb_io_in_0_bits_data_data = useForwardData ? io_in_bits_forwardData_data_data : _dataReadArray_T_10; // @[src/main/scala/nutcore/mem/Cache.scala 275:21]
  assign dataWriteArb_io_in_0_bits_waymask = io_in_bits_waymask; // @[src/main/scala/nutcore/mem/Cache.scala 284:29 src/main/scala/utils/SRAMTemplate.scala 38:24]
  assign dataWriteArb_io_in_1_valid = _readingFirst_T_3 & _readingFirst_T_1; // @[src/main/scala/nutcore/mem/Cache.scala 404:39]
  assign dataWriteArb_io_in_1_bits_setIdx = {addr_index,readBeatCnt_value}; // @[src/main/scala/nutcore/mem/Cache.scala 404:72]
  assign dataWriteArb_io_in_1_bits_data_data = io_mem_resp_bits_rdata; // @[src/main/scala/utils/BitUtils.scala 34:26]
  assign dataWriteArb_io_in_1_bits_waymask = io_in_bits_waymask; // @[src/main/scala/nutcore/mem/Cache.scala 403:32 src/main/scala/utils/SRAMTemplate.scala 38:24]
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/nutcore/mem/Cache.scala 294:22]
      state <= 4'h0; // @[src/main/scala/nutcore/mem/Cache.scala 294:22]
    end else if (4'h0 == state) begin // @[src/main/scala/nutcore/mem/Cache.scala 353:18]
      if ((miss | mmio) & ~io_flush) begin // @[src/main/scala/nutcore/mem/Cache.scala 366:49]
        if (mmio) begin // @[src/main/scala/nutcore/mem/Cache.scala 367:21]
          state <= 4'h5;
        end else begin
          state <= 4'h1;
        end
      end
    end else if (4'h5 == state) begin // @[src/main/scala/nutcore/mem/Cache.scala 353:18]
      if (_T_41) begin // @[src/main/scala/nutcore/mem/Cache.scala 371:46]
        state <= 4'h6; // @[src/main/scala/nutcore/mem/Cache.scala 371:54]
      end
    end else if (4'h6 == state) begin // @[src/main/scala/nutcore/mem/Cache.scala 353:18]
      state <= _GEN_26;
    end else begin
      state <= _GEN_56;
    end
    if (reset) begin // @[src/main/scala/nutcore/mem/Cache.scala 295:26]
      needFlush <= 1'h0; // @[src/main/scala/nutcore/mem/Cache.scala 295:26]
    end else if (_T_5 & needFlush) begin // @[src/main/scala/nutcore/mem/Cache.scala 298:35]
      needFlush <= 1'h0; // @[src/main/scala/nutcore/mem/Cache.scala 298:47]
    end else begin
      needFlush <= _GEN_1;
    end
    if (reset) begin // @[src/main/scala/chisel3/util/Counter.scala 61:40]
      readBeatCnt_value <= 3'h0; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end else if (!(4'h0 == state)) begin // @[src/main/scala/nutcore/mem/Cache.scala 353:18]
      if (!(4'h5 == state)) begin // @[src/main/scala/nutcore/mem/Cache.scala 353:18]
        if (!(4'h6 == state)) begin // @[src/main/scala/nutcore/mem/Cache.scala 353:18]
          readBeatCnt_value <= _GEN_55;
        end
      end
    end
    if (reset) begin // @[src/main/scala/chisel3/util/Counter.scala 61:40]
      writeBeatCnt_value <= 3'h0; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end else if (!(4'h0 == state)) begin // @[src/main/scala/nutcore/mem/Cache.scala 353:18]
      if (!(4'h5 == state)) begin // @[src/main/scala/nutcore/mem/Cache.scala 353:18]
        if (!(4'h6 == state)) begin // @[src/main/scala/nutcore/mem/Cache.scala 353:18]
          writeBeatCnt_value <= _GEN_59;
        end
      end
    end
    if (reset) begin // @[src/main/scala/nutcore/mem/Cache.scala 304:23]
      state2 <= 2'h0; // @[src/main/scala/nutcore/mem/Cache.scala 304:23]
    end else if (2'h0 == state2) begin // @[src/main/scala/nutcore/mem/Cache.scala 311:19]
      if (_T_23) begin // @[src/main/scala/nutcore/mem/Cache.scala 312:51]
        state2 <= 2'h1; // @[src/main/scala/nutcore/mem/Cache.scala 312:60]
      end
    end else if (2'h1 == state2) begin // @[src/main/scala/nutcore/mem/Cache.scala 311:19]
      state2 <= 2'h2; // @[src/main/scala/nutcore/mem/Cache.scala 313:35]
    end else if (2'h2 == state2) begin // @[src/main/scala/nutcore/mem/Cache.scala 311:19]
      state2 <= _GEN_8;
    end
    if (state2 == 2'h1) begin // @[src/main/scala/nutcore/mem/Cache.scala 308:26]
      dataWay_0_data <= io_dataReadBus_resp_data_0_data; // @[src/main/scala/nutcore/mem/Cache.scala 308:26]
    end
    if (state2 == 2'h1) begin // @[src/main/scala/nutcore/mem/Cache.scala 308:26]
      dataWay_1_data <= io_dataReadBus_resp_data_1_data; // @[src/main/scala/nutcore/mem/Cache.scala 308:26]
    end
    if (state2 == 2'h1) begin // @[src/main/scala/nutcore/mem/Cache.scala 308:26]
      dataWay_2_data <= io_dataReadBus_resp_data_2_data; // @[src/main/scala/nutcore/mem/Cache.scala 308:26]
    end
    if (state2 == 2'h1) begin // @[src/main/scala/nutcore/mem/Cache.scala 308:26]
      dataWay_3_data <= io_dataReadBus_resp_data_3_data; // @[src/main/scala/nutcore/mem/Cache.scala 308:26]
    end
    if (reset) begin // @[src/main/scala/nutcore/mem/Cache.scala 336:31]
      afterFirstRead <= 1'h0; // @[src/main/scala/nutcore/mem/Cache.scala 336:31]
    end else if (4'h0 == state) begin // @[src/main/scala/nutcore/mem/Cache.scala 353:18]
      afterFirstRead <= 1'h0; // @[src/main/scala/nutcore/mem/Cache.scala 355:22]
    end else if (!(4'h5 == state)) begin // @[src/main/scala/nutcore/mem/Cache.scala 353:18]
      if (!(4'h6 == state)) begin // @[src/main/scala/nutcore/mem/Cache.scala 353:18]
        afterFirstRead <= _GEN_57;
      end
    end
    if (reset) begin // @[src/main/scala/nutcore/mem/Cache.scala 337:33]
      alreadyOutFire <= 1'h0; // @[src/main/scala/nutcore/mem/Cache.scala 337:33]
    end else if (4'h0 == state) begin // @[src/main/scala/nutcore/mem/Cache.scala 353:18]
      alreadyOutFire <= 1'h0; // @[src/main/scala/nutcore/mem/Cache.scala 356:22]
    end else begin
      alreadyOutFire <= _GEN_12;
    end
    if (_inRdataRegDemand_T_2) begin // @[src/main/scala/nutcore/mem/Cache.scala 339:35]
      if (mmio) begin // @[src/main/scala/nutcore/mem/Cache.scala 339:39]
        inRdataRegDemand <= io_mmio_resp_bits_rdata;
      end else begin
        inRdataRegDemand <= io_mem_resp_bits_rdata;
      end
    end
    if (reset) begin // @[src/main/scala/utils/GTimer.scala 24:20]
      c <= 64'h0; // @[src/main/scala/utils/GTimer.scala 24:20]
    end else begin
      c <= _c_T_1; // @[src/main/scala/utils/GTimer.scala 25:7]
    end
    if (reset) begin // @[src/main/scala/utils/GTimer.scala 24:20]
      c_1 <= 64'h0; // @[src/main/scala/utils/GTimer.scala 24:20]
    end else begin
      c_1 <= _c_T_3; // @[src/main/scala/utils/GTimer.scala 25:7]
    end
    if (reset) begin // @[src/main/scala/utils/GTimer.scala 24:20]
      c_2 <= 64'h0; // @[src/main/scala/utils/GTimer.scala 24:20]
    end else begin
      c_2 <= _c_T_5; // @[src/main/scala/utils/GTimer.scala 25:7]
    end
    if (reset) begin // @[src/main/scala/utils/GTimer.scala 24:20]
      c_3 <= 64'h0; // @[src/main/scala/utils/GTimer.scala 24:20]
    end else begin
      c_3 <= _c_T_7; // @[src/main/scala/utils/GTimer.scala 25:7]
    end
    if (reset) begin // @[src/main/scala/utils/GTimer.scala 24:20]
      c_4 <= 64'h0; // @[src/main/scala/utils/GTimer.scala 24:20]
    end else begin
      c_4 <= _c_T_9; // @[src/main/scala/utils/GTimer.scala 25:7]
    end
    if (reset) begin // @[src/main/scala/utils/GTimer.scala 24:20]
      c_5 <= 64'h0; // @[src/main/scala/utils/GTimer.scala 24:20]
    end else begin
      c_5 <= _c_T_11; // @[src/main/scala/utils/GTimer.scala 25:7]
    end
    if (reset) begin // @[src/main/scala/utils/GTimer.scala 24:20]
      c_6 <= 64'h0; // @[src/main/scala/utils/GTimer.scala 24:20]
    end else begin
      c_6 <= _c_T_13; // @[src/main/scala/utils/GTimer.scala 25:7]
    end
    if (reset) begin // @[src/main/scala/utils/GTimer.scala 24:20]
      c_7 <= 64'h0; // @[src/main/scala/utils/GTimer.scala 24:20]
    end else begin
      c_7 <= _c_T_15; // @[src/main/scala/utils/GTimer.scala 25:7]
    end
    if (reset) begin // @[src/main/scala/utils/GTimer.scala 24:20]
      c_8 <= 64'h0; // @[src/main/scala/utils/GTimer.scala 24:20]
    end else begin
      c_8 <= _c_T_17; // @[src/main/scala/utils/GTimer.scala 25:7]
    end
    if (reset) begin // @[src/main/scala/utils/GTimer.scala 24:20]
      c_9 <= 64'h0; // @[src/main/scala/utils/GTimer.scala 24:20]
    end else begin
      c_9 <= _c_T_19; // @[src/main/scala/utils/GTimer.scala 25:7]
    end
    if (reset) begin // @[src/main/scala/utils/GTimer.scala 24:20]
      c_10 <= 64'h0; // @[src/main/scala/utils/GTimer.scala 24:20]
    end else begin
      c_10 <= _c_T_21; // @[src/main/scala/utils/GTimer.scala 25:7]
    end
    if (reset) begin // @[src/main/scala/utils/GTimer.scala 24:20]
      c_11 <= 64'h0; // @[src/main/scala/utils/GTimer.scala 24:20]
    end else begin
      c_11 <= _c_T_23; // @[src/main/scala/utils/GTimer.scala 25:7]
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~(mmio & hit))) begin
          $fwrite(32'h80000002,
            "Assertion failed: MMIO request should not hit in cache\n    at Cache.scala:265 assert(!(mmio && hit), \"MMIO request should not hit in cache\")\n"
            ); // @[src/main/scala/nutcore/mem/Cache.scala 265:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~(mmio & hit)) & ~reset) begin
          $fatal; // @[src/main/scala/nutcore/mem/Cache.scala 265:9]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_3) begin
          $fwrite(32'h80000002,"[%d] CacheStage3: ",c); // @[src/main/scala/utils/Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_3) begin
          $fwrite(32'h80000002," metaread idx %x waymask %b metas %x%x:%x %x%x:%x %x%x:%x %x%x:%x %x\n",addr_index,
            io_in_bits_waymask,io_in_bits_metas_0_valid,io_in_bits_metas_0_dirty,io_in_bits_metas_0_tag,
            io_in_bits_metas_1_valid,io_in_bits_metas_1_dirty,io_in_bits_metas_1_tag,io_in_bits_metas_2_valid,
            io_in_bits_metas_2_dirty,io_in_bits_metas_2_tag,io_in_bits_metas_3_valid,io_in_bits_metas_3_dirty,
            io_in_bits_metas_3_tag,_T_89); // @[src/main/scala/utils/Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_96 & _T_3) begin
          $fwrite(32'h80000002,"[%d] CacheStage3: ",c_2); // @[src/main/scala/utils/Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_96 & _T_3) begin
          $fwrite(32'h80000002,"%d: [icache S3]: metawrite idx %x wmask %b meta %x%x:%x\n",c_1,
            io_metaWriteBus_req_bits_setIdx,io_metaWriteBus_req_bits_waymask,io_metaWriteBus_req_bits_data_valid,
            io_metaWriteBus_req_bits_data_dirty,io_metaWriteBus_req_bits_data_tag); // @[src/main/scala/utils/Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_3) begin
          $fwrite(32'h80000002,"[%d] CacheStage3: ",c_3); // @[src/main/scala/utils/Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_3) begin
          $fwrite(32'h80000002,
            " in.ready = %d, in.valid = %d, hit = %x, state = %d, addr = %x cmd:%d probe:%d isFinish:%d\n",io_in_ready,
            io_in_valid,hit,state,io_in_bits_req_addr,4'h0,1'h0,io_isFinish); // @[src/main/scala/utils/Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_3) begin
          $fwrite(32'h80000002,"[%d] CacheStage3: ",c_4); // @[src/main/scala/utils/Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_3) begin
          $fwrite(32'h80000002," out.valid:%d rdata:%x cmd:%d user:%x id:%x \n",io_out_valid,io_out_bits_rdata,
            io_out_bits_cmd,io_out_bits_user,1'h0); // @[src/main/scala/utils/Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_3) begin
          $fwrite(32'h80000002,"[%d] CacheStage3: ",c_5); // @[src/main/scala/utils/Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_3) begin
          $fwrite(32'h80000002," DHW: (%d, %d), data:%x setIdx:%x MHW:(%d, %d)\n",1'h0,1'h1,dataRead,dataHitWriteBus_x3,1'h0
            ,1'h1); // @[src/main/scala/utils/Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_3) begin
          $fwrite(32'h80000002,"[%d] CacheStage3: ",c_6); // @[src/main/scala/utils/Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_3) begin
          $fwrite(32'h80000002," DreadCache: %x \n",_T_89); // @[src/main/scala/utils/Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_3) begin
          $fwrite(32'h80000002,"[%d] CacheStage3: ",c_7); // @[src/main/scala/utils/Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_3) begin
          $fwrite(32'h80000002," useFD:%d isFD:%d FD:%x DreadArray:%x dataRead:%x inwaymask:%x FDwaymask:%x \n",
            useForwardData,io_in_bits_isForwardData,io_in_bits_forwardData_data_data,_dataReadArray_T_10,dataRead,
            io_in_bits_waymask,io_in_bits_forwardData_waymask); // @[src/main/scala/utils/Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_128 & _T_3) begin
          $fwrite(32'h80000002,"[%d] CacheStage3: ",c_8); // @[src/main/scala/utils/Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_128 & _T_3) begin
          $fwrite(32'h80000002,"[WB] waymask: %b data:%x setIdx:%x\n",io_dataWriteBus_req_bits_waymask,
            io_dataWriteBus_req_bits_data_data,io_dataWriteBus_req_bits_setIdx); // @[src/main/scala/utils/Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_140 & _T_3) begin
          $fwrite(32'h80000002,"[%d] CacheStage3: ",c_9); // @[src/main/scala/utils/Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_140 & _T_3) begin
          $fwrite(32'h80000002,"[COUTW] cnt %x addr %x data %x cmd %x size %x wmask %x tag %x idx %x waymask %b \n",
            writeBeatCnt_value,io_mem_req_bits_addr,io_mem_req_bits_wdata,io_mem_req_bits_cmd,io_mem_req_bits_size,
            io_mem_req_bits_wmask,addr_tag,addr_index,io_in_bits_waymask); // @[src/main/scala/utils/Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_152 & _T_3) begin
          $fwrite(32'h80000002,"[%d] CacheStage3: ",c_10); // @[src/main/scala/utils/Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_152 & _T_3) begin
          $fwrite(32'h80000002,"[COUTR] addr %x tag %x idx %x waymask %b \n",io_mem_req_bits_addr,addr_tag,addr_index,
            io_in_bits_waymask); // @[src/main/scala/utils/Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_164 & _T_3) begin
          $fwrite(32'h80000002,"[%d] CacheStage3: ",c_11); // @[src/main/scala/utils/Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_164 & _T_3) begin
          $fwrite(32'h80000002,"[COUTR] cnt %x data %x tag %x idx %x waymask %b \n",readBeatCnt_value,
            io_mem_resp_bits_rdata,addr_tag,addr_index,io_in_bits_waymask); // @[src/main/scala/utils/Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[3:0];
  _RAND_1 = {1{`RANDOM}};
  needFlush = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  readBeatCnt_value = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  writeBeatCnt_value = _RAND_3[2:0];
  _RAND_4 = {1{`RANDOM}};
  state2 = _RAND_4[1:0];
  _RAND_5 = {2{`RANDOM}};
  dataWay_0_data = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  dataWay_1_data = _RAND_6[63:0];
  _RAND_7 = {2{`RANDOM}};
  dataWay_2_data = _RAND_7[63:0];
  _RAND_8 = {2{`RANDOM}};
  dataWay_3_data = _RAND_8[63:0];
  _RAND_9 = {1{`RANDOM}};
  afterFirstRead = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  alreadyOutFire = _RAND_10[0:0];
  _RAND_11 = {2{`RANDOM}};
  inRdataRegDemand = _RAND_11[63:0];
  _RAND_12 = {2{`RANDOM}};
  c = _RAND_12[63:0];
  _RAND_13 = {2{`RANDOM}};
  c_1 = _RAND_13[63:0];
  _RAND_14 = {2{`RANDOM}};
  c_2 = _RAND_14[63:0];
  _RAND_15 = {2{`RANDOM}};
  c_3 = _RAND_15[63:0];
  _RAND_16 = {2{`RANDOM}};
  c_4 = _RAND_16[63:0];
  _RAND_17 = {2{`RANDOM}};
  c_5 = _RAND_17[63:0];
  _RAND_18 = {2{`RANDOM}};
  c_6 = _RAND_18[63:0];
  _RAND_19 = {2{`RANDOM}};
  c_7 = _RAND_19[63:0];
  _RAND_20 = {2{`RANDOM}};
  c_8 = _RAND_20[63:0];
  _RAND_21 = {2{`RANDOM}};
  c_9 = _RAND_21[63:0];
  _RAND_22 = {2{`RANDOM}};
  c_10 = _RAND_22[63:0];
  _RAND_23 = {2{`RANDOM}};
  c_11 = _RAND_23[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module SRAMTemplate_1(
  input         clock,
  input         reset,
  output        io_r_req_ready, // @[src/main/scala/utils/SRAMTemplate.scala 70:14]
  input         io_r_req_valid, // @[src/main/scala/utils/SRAMTemplate.scala 70:14]
  input  [6:0]  io_r_req_bits_setIdx, // @[src/main/scala/utils/SRAMTemplate.scala 70:14]
  output [18:0] io_r_resp_data_0_tag, // @[src/main/scala/utils/SRAMTemplate.scala 70:14]
  output        io_r_resp_data_0_valid, // @[src/main/scala/utils/SRAMTemplate.scala 70:14]
  output        io_r_resp_data_0_dirty, // @[src/main/scala/utils/SRAMTemplate.scala 70:14]
  output [18:0] io_r_resp_data_1_tag, // @[src/main/scala/utils/SRAMTemplate.scala 70:14]
  output        io_r_resp_data_1_valid, // @[src/main/scala/utils/SRAMTemplate.scala 70:14]
  output        io_r_resp_data_1_dirty, // @[src/main/scala/utils/SRAMTemplate.scala 70:14]
  output [18:0] io_r_resp_data_2_tag, // @[src/main/scala/utils/SRAMTemplate.scala 70:14]
  output        io_r_resp_data_2_valid, // @[src/main/scala/utils/SRAMTemplate.scala 70:14]
  output        io_r_resp_data_2_dirty, // @[src/main/scala/utils/SRAMTemplate.scala 70:14]
  output [18:0] io_r_resp_data_3_tag, // @[src/main/scala/utils/SRAMTemplate.scala 70:14]
  output        io_r_resp_data_3_valid, // @[src/main/scala/utils/SRAMTemplate.scala 70:14]
  output        io_r_resp_data_3_dirty, // @[src/main/scala/utils/SRAMTemplate.scala 70:14]
  input         io_w_req_valid, // @[src/main/scala/utils/SRAMTemplate.scala 70:14]
  input  [6:0]  io_w_req_bits_setIdx, // @[src/main/scala/utils/SRAMTemplate.scala 70:14]
  input  [18:0] io_w_req_bits_data_tag, // @[src/main/scala/utils/SRAMTemplate.scala 70:14]
  input         io_w_req_bits_data_dirty, // @[src/main/scala/utils/SRAMTemplate.scala 70:14]
  input  [3:0]  io_w_req_bits_waymask // @[src/main/scala/utils/SRAMTemplate.scala 70:14]
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_9;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
`endif // RANDOMIZE_REG_INIT
  reg [20:0] array_0 [0:127]; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
  wire  array_0_rdata_MPORT_en; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
  wire [6:0] array_0_rdata_MPORT_addr; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
  wire [20:0] array_0_rdata_MPORT_data; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
  wire [20:0] array_0_MPORT_data; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
  wire [6:0] array_0_MPORT_addr; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
  wire  array_0_MPORT_mask; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
  wire  array_0_MPORT_en; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
  reg  array_0_rdata_MPORT_en_pipe_0;
  reg [6:0] array_0_rdata_MPORT_addr_pipe_0;
  reg [20:0] array_1 [0:127]; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
  wire  array_1_rdata_MPORT_en; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
  wire [6:0] array_1_rdata_MPORT_addr; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
  wire [20:0] array_1_rdata_MPORT_data; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
  wire [20:0] array_1_MPORT_data; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
  wire [6:0] array_1_MPORT_addr; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
  wire  array_1_MPORT_mask; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
  wire  array_1_MPORT_en; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
  reg  array_1_rdata_MPORT_en_pipe_0;
  reg [6:0] array_1_rdata_MPORT_addr_pipe_0;
  reg [20:0] array_2 [0:127]; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
  wire  array_2_rdata_MPORT_en; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
  wire [6:0] array_2_rdata_MPORT_addr; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
  wire [20:0] array_2_rdata_MPORT_data; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
  wire [20:0] array_2_MPORT_data; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
  wire [6:0] array_2_MPORT_addr; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
  wire  array_2_MPORT_mask; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
  wire  array_2_MPORT_en; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
  reg  array_2_rdata_MPORT_en_pipe_0;
  reg [6:0] array_2_rdata_MPORT_addr_pipe_0;
  reg [20:0] array_3 [0:127]; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
  wire  array_3_rdata_MPORT_en; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
  wire [6:0] array_3_rdata_MPORT_addr; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
  wire [20:0] array_3_rdata_MPORT_data; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
  wire [20:0] array_3_MPORT_data; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
  wire [6:0] array_3_MPORT_addr; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
  wire  array_3_MPORT_mask; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
  wire  array_3_MPORT_en; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
  reg  array_3_rdata_MPORT_en_pipe_0;
  reg [6:0] array_3_rdata_MPORT_addr_pipe_0;
  reg  resetState; // @[src/main/scala/utils/SRAMTemplate.scala 80:30]
  reg [6:0] resetSet; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
  wire  wrap_wrap = resetSet == 7'h7f; // @[src/main/scala/chisel3/util/Counter.scala 73:24]
  wire [6:0] _wrap_value_T_1 = resetSet + 7'h1; // @[src/main/scala/chisel3/util/Counter.scala 77:24]
  wire  resetFinish = resetState & wrap_wrap; // @[src/main/scala/chisel3/util/Counter.scala 118:{16,23} 117:24]
  wire  _GEN_2 = resetFinish ? 1'h0 : resetState; // @[src/main/scala/utils/SRAMTemplate.scala 82:24 80:30 82:38]
  wire  wen = io_w_req_valid | resetState; // @[src/main/scala/utils/SRAMTemplate.scala 88:52]
  wire  _realRen_T = ~wen; // @[src/main/scala/utils/SRAMTemplate.scala 89:41]
  wire [20:0] _wdataword_T = {io_w_req_bits_data_tag,1'h1,io_w_req_bits_data_dirty}; // @[src/main/scala/utils/SRAMTemplate.scala 92:78]
  wire [3:0] waymask = resetState ? 4'hf : io_w_req_bits_waymask; // @[src/main/scala/utils/SRAMTemplate.scala 93:20]
  wire [20:0] _rdata_WIRE_1 = array_0_rdata_MPORT_data; // @[src/main/scala/utils/SRAMTemplate.scala 98:{78,78}]
  wire [20:0] _rdata_WIRE_2 = array_1_rdata_MPORT_data; // @[src/main/scala/utils/SRAMTemplate.scala 98:{78,78}]
  wire [20:0] _rdata_WIRE_3 = array_2_rdata_MPORT_data; // @[src/main/scala/utils/SRAMTemplate.scala 98:{78,78}]
  wire [20:0] _rdata_WIRE_4 = array_3_rdata_MPORT_data; // @[src/main/scala/utils/SRAMTemplate.scala 98:{78,78}]
  assign array_0_rdata_MPORT_en = array_0_rdata_MPORT_en_pipe_0;
  assign array_0_rdata_MPORT_addr = array_0_rdata_MPORT_addr_pipe_0;
  assign array_0_rdata_MPORT_data = array_0[array_0_rdata_MPORT_addr]; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
  assign array_0_MPORT_data = resetState ? 21'h0 : _wdataword_T;
  assign array_0_MPORT_addr = resetState ? resetSet : io_w_req_bits_setIdx;
  assign array_0_MPORT_mask = waymask[0];
  assign array_0_MPORT_en = io_w_req_valid | resetState;
  assign array_1_rdata_MPORT_en = array_1_rdata_MPORT_en_pipe_0;
  assign array_1_rdata_MPORT_addr = array_1_rdata_MPORT_addr_pipe_0;
  assign array_1_rdata_MPORT_data = array_1[array_1_rdata_MPORT_addr]; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
  assign array_1_MPORT_data = resetState ? 21'h0 : _wdataword_T;
  assign array_1_MPORT_addr = resetState ? resetSet : io_w_req_bits_setIdx;
  assign array_1_MPORT_mask = waymask[1];
  assign array_1_MPORT_en = io_w_req_valid | resetState;
  assign array_2_rdata_MPORT_en = array_2_rdata_MPORT_en_pipe_0;
  assign array_2_rdata_MPORT_addr = array_2_rdata_MPORT_addr_pipe_0;
  assign array_2_rdata_MPORT_data = array_2[array_2_rdata_MPORT_addr]; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
  assign array_2_MPORT_data = resetState ? 21'h0 : _wdataword_T;
  assign array_2_MPORT_addr = resetState ? resetSet : io_w_req_bits_setIdx;
  assign array_2_MPORT_mask = waymask[2];
  assign array_2_MPORT_en = io_w_req_valid | resetState;
  assign array_3_rdata_MPORT_en = array_3_rdata_MPORT_en_pipe_0;
  assign array_3_rdata_MPORT_addr = array_3_rdata_MPORT_addr_pipe_0;
  assign array_3_rdata_MPORT_data = array_3[array_3_rdata_MPORT_addr]; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
  assign array_3_MPORT_data = resetState ? 21'h0 : _wdataword_T;
  assign array_3_MPORT_addr = resetState ? resetSet : io_w_req_bits_setIdx;
  assign array_3_MPORT_mask = waymask[3];
  assign array_3_MPORT_en = io_w_req_valid | resetState;
  assign io_r_req_ready = ~resetState & _realRen_T; // @[src/main/scala/utils/SRAMTemplate.scala 101:33]
  assign io_r_resp_data_0_tag = _rdata_WIRE_1[20:2]; // @[src/main/scala/utils/SRAMTemplate.scala 98:78]
  assign io_r_resp_data_0_valid = _rdata_WIRE_1[1]; // @[src/main/scala/utils/SRAMTemplate.scala 98:78]
  assign io_r_resp_data_0_dirty = _rdata_WIRE_1[0]; // @[src/main/scala/utils/SRAMTemplate.scala 98:78]
  assign io_r_resp_data_1_tag = _rdata_WIRE_2[20:2]; // @[src/main/scala/utils/SRAMTemplate.scala 98:78]
  assign io_r_resp_data_1_valid = _rdata_WIRE_2[1]; // @[src/main/scala/utils/SRAMTemplate.scala 98:78]
  assign io_r_resp_data_1_dirty = _rdata_WIRE_2[0]; // @[src/main/scala/utils/SRAMTemplate.scala 98:78]
  assign io_r_resp_data_2_tag = _rdata_WIRE_3[20:2]; // @[src/main/scala/utils/SRAMTemplate.scala 98:78]
  assign io_r_resp_data_2_valid = _rdata_WIRE_3[1]; // @[src/main/scala/utils/SRAMTemplate.scala 98:78]
  assign io_r_resp_data_2_dirty = _rdata_WIRE_3[0]; // @[src/main/scala/utils/SRAMTemplate.scala 98:78]
  assign io_r_resp_data_3_tag = _rdata_WIRE_4[20:2]; // @[src/main/scala/utils/SRAMTemplate.scala 98:78]
  assign io_r_resp_data_3_valid = _rdata_WIRE_4[1]; // @[src/main/scala/utils/SRAMTemplate.scala 98:78]
  assign io_r_resp_data_3_dirty = _rdata_WIRE_4[0]; // @[src/main/scala/utils/SRAMTemplate.scala 98:78]
  always @(posedge clock) begin
    if (array_0_MPORT_en & array_0_MPORT_mask) begin
      array_0[array_0_MPORT_addr] <= array_0_MPORT_data; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
    end
    array_0_rdata_MPORT_en_pipe_0 <= io_r_req_valid & _realRen_T;
    if (io_r_req_valid & _realRen_T) begin
      array_0_rdata_MPORT_addr_pipe_0 <= io_r_req_bits_setIdx;
    end
    if (array_1_MPORT_en & array_1_MPORT_mask) begin
      array_1[array_1_MPORT_addr] <= array_1_MPORT_data; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
    end
    array_1_rdata_MPORT_en_pipe_0 <= io_r_req_valid & _realRen_T;
    if (io_r_req_valid & _realRen_T) begin
      array_1_rdata_MPORT_addr_pipe_0 <= io_r_req_bits_setIdx;
    end
    if (array_2_MPORT_en & array_2_MPORT_mask) begin
      array_2[array_2_MPORT_addr] <= array_2_MPORT_data; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
    end
    array_2_rdata_MPORT_en_pipe_0 <= io_r_req_valid & _realRen_T;
    if (io_r_req_valid & _realRen_T) begin
      array_2_rdata_MPORT_addr_pipe_0 <= io_r_req_bits_setIdx;
    end
    if (array_3_MPORT_en & array_3_MPORT_mask) begin
      array_3[array_3_MPORT_addr] <= array_3_MPORT_data; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
    end
    array_3_rdata_MPORT_en_pipe_0 <= io_r_req_valid & _realRen_T;
    if (io_r_req_valid & _realRen_T) begin
      array_3_rdata_MPORT_addr_pipe_0 <= io_r_req_bits_setIdx;
    end
    resetState <= reset | _GEN_2; // @[src/main/scala/utils/SRAMTemplate.scala 80:{30,30}]
    if (reset) begin // @[src/main/scala/chisel3/util/Counter.scala 61:40]
      resetSet <= 7'h0; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end else if (resetState) begin // @[src/main/scala/chisel3/util/Counter.scala 118:16]
      resetSet <= _wrap_value_T_1; // @[src/main/scala/chisel3/util/Counter.scala 77:15]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 128; initvar = initvar+1)
    array_0[initvar] = _RAND_0[20:0];
  _RAND_3 = {1{`RANDOM}};
  for (initvar = 0; initvar < 128; initvar = initvar+1)
    array_1[initvar] = _RAND_3[20:0];
  _RAND_6 = {1{`RANDOM}};
  for (initvar = 0; initvar < 128; initvar = initvar+1)
    array_2[initvar] = _RAND_6[20:0];
  _RAND_9 = {1{`RANDOM}};
  for (initvar = 0; initvar < 128; initvar = initvar+1)
    array_3[initvar] = _RAND_9[20:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  array_0_rdata_MPORT_en_pipe_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  array_0_rdata_MPORT_addr_pipe_0 = _RAND_2[6:0];
  _RAND_4 = {1{`RANDOM}};
  array_1_rdata_MPORT_en_pipe_0 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  array_1_rdata_MPORT_addr_pipe_0 = _RAND_5[6:0];
  _RAND_7 = {1{`RANDOM}};
  array_2_rdata_MPORT_en_pipe_0 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  array_2_rdata_MPORT_addr_pipe_0 = _RAND_8[6:0];
  _RAND_10 = {1{`RANDOM}};
  array_3_rdata_MPORT_en_pipe_0 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  array_3_rdata_MPORT_addr_pipe_0 = _RAND_11[6:0];
  _RAND_12 = {1{`RANDOM}};
  resetState = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  resetSet = _RAND_13[6:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Arbiter_2(
  output       io_in_0_ready, // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
  input        io_in_0_valid, // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
  input  [6:0] io_in_0_bits_setIdx, // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
  input        io_out_ready, // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
  output       io_out_valid, // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
  output [6:0] io_out_bits_setIdx // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
);
  assign io_in_0_ready = io_out_ready; // @[src/main/scala/chisel3/util/Arbiter.scala 147:19]
  assign io_out_valid = io_in_0_valid; // @[src/main/scala/chisel3/util/Arbiter.scala 148:31]
  assign io_out_bits_setIdx = io_in_0_bits_setIdx; // @[src/main/scala/chisel3/util/Arbiter.scala 137:15]
endmodule
module SRAMTemplateWithArbiter(
  input         clock,
  input         reset,
  output        io_r_0_req_ready, // @[src/main/scala/utils/SRAMTemplate.scala 116:14]
  input         io_r_0_req_valid, // @[src/main/scala/utils/SRAMTemplate.scala 116:14]
  input  [6:0]  io_r_0_req_bits_setIdx, // @[src/main/scala/utils/SRAMTemplate.scala 116:14]
  output [18:0] io_r_0_resp_data_0_tag, // @[src/main/scala/utils/SRAMTemplate.scala 116:14]
  output        io_r_0_resp_data_0_valid, // @[src/main/scala/utils/SRAMTemplate.scala 116:14]
  output        io_r_0_resp_data_0_dirty, // @[src/main/scala/utils/SRAMTemplate.scala 116:14]
  output [18:0] io_r_0_resp_data_1_tag, // @[src/main/scala/utils/SRAMTemplate.scala 116:14]
  output        io_r_0_resp_data_1_valid, // @[src/main/scala/utils/SRAMTemplate.scala 116:14]
  output        io_r_0_resp_data_1_dirty, // @[src/main/scala/utils/SRAMTemplate.scala 116:14]
  output [18:0] io_r_0_resp_data_2_tag, // @[src/main/scala/utils/SRAMTemplate.scala 116:14]
  output        io_r_0_resp_data_2_valid, // @[src/main/scala/utils/SRAMTemplate.scala 116:14]
  output        io_r_0_resp_data_2_dirty, // @[src/main/scala/utils/SRAMTemplate.scala 116:14]
  output [18:0] io_r_0_resp_data_3_tag, // @[src/main/scala/utils/SRAMTemplate.scala 116:14]
  output        io_r_0_resp_data_3_valid, // @[src/main/scala/utils/SRAMTemplate.scala 116:14]
  output        io_r_0_resp_data_3_dirty, // @[src/main/scala/utils/SRAMTemplate.scala 116:14]
  input         io_w_req_valid, // @[src/main/scala/utils/SRAMTemplate.scala 116:14]
  input  [6:0]  io_w_req_bits_setIdx, // @[src/main/scala/utils/SRAMTemplate.scala 116:14]
  input  [18:0] io_w_req_bits_data_tag, // @[src/main/scala/utils/SRAMTemplate.scala 116:14]
  input         io_w_req_bits_data_dirty, // @[src/main/scala/utils/SRAMTemplate.scala 116:14]
  input  [3:0]  io_w_req_bits_waymask // @[src/main/scala/utils/SRAMTemplate.scala 116:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
`endif // RANDOMIZE_REG_INIT
  wire  ram_clock; // @[src/main/scala/utils/SRAMTemplate.scala 121:19]
  wire  ram_reset; // @[src/main/scala/utils/SRAMTemplate.scala 121:19]
  wire  ram_io_r_req_ready; // @[src/main/scala/utils/SRAMTemplate.scala 121:19]
  wire  ram_io_r_req_valid; // @[src/main/scala/utils/SRAMTemplate.scala 121:19]
  wire [6:0] ram_io_r_req_bits_setIdx; // @[src/main/scala/utils/SRAMTemplate.scala 121:19]
  wire [18:0] ram_io_r_resp_data_0_tag; // @[src/main/scala/utils/SRAMTemplate.scala 121:19]
  wire  ram_io_r_resp_data_0_valid; // @[src/main/scala/utils/SRAMTemplate.scala 121:19]
  wire  ram_io_r_resp_data_0_dirty; // @[src/main/scala/utils/SRAMTemplate.scala 121:19]
  wire [18:0] ram_io_r_resp_data_1_tag; // @[src/main/scala/utils/SRAMTemplate.scala 121:19]
  wire  ram_io_r_resp_data_1_valid; // @[src/main/scala/utils/SRAMTemplate.scala 121:19]
  wire  ram_io_r_resp_data_1_dirty; // @[src/main/scala/utils/SRAMTemplate.scala 121:19]
  wire [18:0] ram_io_r_resp_data_2_tag; // @[src/main/scala/utils/SRAMTemplate.scala 121:19]
  wire  ram_io_r_resp_data_2_valid; // @[src/main/scala/utils/SRAMTemplate.scala 121:19]
  wire  ram_io_r_resp_data_2_dirty; // @[src/main/scala/utils/SRAMTemplate.scala 121:19]
  wire [18:0] ram_io_r_resp_data_3_tag; // @[src/main/scala/utils/SRAMTemplate.scala 121:19]
  wire  ram_io_r_resp_data_3_valid; // @[src/main/scala/utils/SRAMTemplate.scala 121:19]
  wire  ram_io_r_resp_data_3_dirty; // @[src/main/scala/utils/SRAMTemplate.scala 121:19]
  wire  ram_io_w_req_valid; // @[src/main/scala/utils/SRAMTemplate.scala 121:19]
  wire [6:0] ram_io_w_req_bits_setIdx; // @[src/main/scala/utils/SRAMTemplate.scala 121:19]
  wire [18:0] ram_io_w_req_bits_data_tag; // @[src/main/scala/utils/SRAMTemplate.scala 121:19]
  wire  ram_io_w_req_bits_data_dirty; // @[src/main/scala/utils/SRAMTemplate.scala 121:19]
  wire [3:0] ram_io_w_req_bits_waymask; // @[src/main/scala/utils/SRAMTemplate.scala 121:19]
  wire  readArb_io_in_0_ready; // @[src/main/scala/utils/SRAMTemplate.scala 124:23]
  wire  readArb_io_in_0_valid; // @[src/main/scala/utils/SRAMTemplate.scala 124:23]
  wire [6:0] readArb_io_in_0_bits_setIdx; // @[src/main/scala/utils/SRAMTemplate.scala 124:23]
  wire  readArb_io_out_ready; // @[src/main/scala/utils/SRAMTemplate.scala 124:23]
  wire  readArb_io_out_valid; // @[src/main/scala/utils/SRAMTemplate.scala 124:23]
  wire [6:0] readArb_io_out_bits_setIdx; // @[src/main/scala/utils/SRAMTemplate.scala 124:23]
  reg  REG; // @[src/main/scala/utils/SRAMTemplate.scala 130:58]
  reg [18:0] r_0_tag; // @[src/main/scala/utils/Hold.scala 23:65]
  reg  r_0_valid; // @[src/main/scala/utils/Hold.scala 23:65]
  reg  r_0_dirty; // @[src/main/scala/utils/Hold.scala 23:65]
  reg [18:0] r_1_tag; // @[src/main/scala/utils/Hold.scala 23:65]
  reg  r_1_valid; // @[src/main/scala/utils/Hold.scala 23:65]
  reg  r_1_dirty; // @[src/main/scala/utils/Hold.scala 23:65]
  reg [18:0] r_2_tag; // @[src/main/scala/utils/Hold.scala 23:65]
  reg  r_2_valid; // @[src/main/scala/utils/Hold.scala 23:65]
  reg  r_2_dirty; // @[src/main/scala/utils/Hold.scala 23:65]
  reg [18:0] r_3_tag; // @[src/main/scala/utils/Hold.scala 23:65]
  reg  r_3_valid; // @[src/main/scala/utils/Hold.scala 23:65]
  reg  r_3_dirty; // @[src/main/scala/utils/Hold.scala 23:65]
  SRAMTemplate_1 ram ( // @[src/main/scala/utils/SRAMTemplate.scala 121:19]
    .clock(ram_clock),
    .reset(ram_reset),
    .io_r_req_ready(ram_io_r_req_ready),
    .io_r_req_valid(ram_io_r_req_valid),
    .io_r_req_bits_setIdx(ram_io_r_req_bits_setIdx),
    .io_r_resp_data_0_tag(ram_io_r_resp_data_0_tag),
    .io_r_resp_data_0_valid(ram_io_r_resp_data_0_valid),
    .io_r_resp_data_0_dirty(ram_io_r_resp_data_0_dirty),
    .io_r_resp_data_1_tag(ram_io_r_resp_data_1_tag),
    .io_r_resp_data_1_valid(ram_io_r_resp_data_1_valid),
    .io_r_resp_data_1_dirty(ram_io_r_resp_data_1_dirty),
    .io_r_resp_data_2_tag(ram_io_r_resp_data_2_tag),
    .io_r_resp_data_2_valid(ram_io_r_resp_data_2_valid),
    .io_r_resp_data_2_dirty(ram_io_r_resp_data_2_dirty),
    .io_r_resp_data_3_tag(ram_io_r_resp_data_3_tag),
    .io_r_resp_data_3_valid(ram_io_r_resp_data_3_valid),
    .io_r_resp_data_3_dirty(ram_io_r_resp_data_3_dirty),
    .io_w_req_valid(ram_io_w_req_valid),
    .io_w_req_bits_setIdx(ram_io_w_req_bits_setIdx),
    .io_w_req_bits_data_tag(ram_io_w_req_bits_data_tag),
    .io_w_req_bits_data_dirty(ram_io_w_req_bits_data_dirty),
    .io_w_req_bits_waymask(ram_io_w_req_bits_waymask)
  );
  Arbiter_2 readArb ( // @[src/main/scala/utils/SRAMTemplate.scala 124:23]
    .io_in_0_ready(readArb_io_in_0_ready),
    .io_in_0_valid(readArb_io_in_0_valid),
    .io_in_0_bits_setIdx(readArb_io_in_0_bits_setIdx),
    .io_out_ready(readArb_io_out_ready),
    .io_out_valid(readArb_io_out_valid),
    .io_out_bits_setIdx(readArb_io_out_bits_setIdx)
  );
  assign io_r_0_req_ready = readArb_io_in_0_ready; // @[src/main/scala/utils/SRAMTemplate.scala 125:17]
  assign io_r_0_resp_data_0_tag = REG ? ram_io_r_resp_data_0_tag : r_0_tag; // @[src/main/scala/utils/Hold.scala 23:48]
  assign io_r_0_resp_data_0_valid = REG ? ram_io_r_resp_data_0_valid : r_0_valid; // @[src/main/scala/utils/Hold.scala 23:48]
  assign io_r_0_resp_data_0_dirty = REG ? ram_io_r_resp_data_0_dirty : r_0_dirty; // @[src/main/scala/utils/Hold.scala 23:48]
  assign io_r_0_resp_data_1_tag = REG ? ram_io_r_resp_data_1_tag : r_1_tag; // @[src/main/scala/utils/Hold.scala 23:48]
  assign io_r_0_resp_data_1_valid = REG ? ram_io_r_resp_data_1_valid : r_1_valid; // @[src/main/scala/utils/Hold.scala 23:48]
  assign io_r_0_resp_data_1_dirty = REG ? ram_io_r_resp_data_1_dirty : r_1_dirty; // @[src/main/scala/utils/Hold.scala 23:48]
  assign io_r_0_resp_data_2_tag = REG ? ram_io_r_resp_data_2_tag : r_2_tag; // @[src/main/scala/utils/Hold.scala 23:48]
  assign io_r_0_resp_data_2_valid = REG ? ram_io_r_resp_data_2_valid : r_2_valid; // @[src/main/scala/utils/Hold.scala 23:48]
  assign io_r_0_resp_data_2_dirty = REG ? ram_io_r_resp_data_2_dirty : r_2_dirty; // @[src/main/scala/utils/Hold.scala 23:48]
  assign io_r_0_resp_data_3_tag = REG ? ram_io_r_resp_data_3_tag : r_3_tag; // @[src/main/scala/utils/Hold.scala 23:48]
  assign io_r_0_resp_data_3_valid = REG ? ram_io_r_resp_data_3_valid : r_3_valid; // @[src/main/scala/utils/Hold.scala 23:48]
  assign io_r_0_resp_data_3_dirty = REG ? ram_io_r_resp_data_3_dirty : r_3_dirty; // @[src/main/scala/utils/Hold.scala 23:48]
  assign ram_clock = clock;
  assign ram_reset = reset;
  assign ram_io_r_req_valid = readArb_io_out_valid; // @[src/main/scala/utils/SRAMTemplate.scala 126:16]
  assign ram_io_r_req_bits_setIdx = readArb_io_out_bits_setIdx; // @[src/main/scala/utils/SRAMTemplate.scala 126:16]
  assign ram_io_w_req_valid = io_w_req_valid; // @[src/main/scala/utils/SRAMTemplate.scala 122:12]
  assign ram_io_w_req_bits_setIdx = io_w_req_bits_setIdx; // @[src/main/scala/utils/SRAMTemplate.scala 122:12]
  assign ram_io_w_req_bits_data_tag = io_w_req_bits_data_tag; // @[src/main/scala/utils/SRAMTemplate.scala 122:12]
  assign ram_io_w_req_bits_data_dirty = io_w_req_bits_data_dirty; // @[src/main/scala/utils/SRAMTemplate.scala 122:12]
  assign ram_io_w_req_bits_waymask = io_w_req_bits_waymask; // @[src/main/scala/utils/SRAMTemplate.scala 122:12]
  assign readArb_io_in_0_valid = io_r_0_req_valid; // @[src/main/scala/utils/SRAMTemplate.scala 125:17]
  assign readArb_io_in_0_bits_setIdx = io_r_0_req_bits_setIdx; // @[src/main/scala/utils/SRAMTemplate.scala 125:17]
  assign readArb_io_out_ready = ram_io_r_req_ready; // @[src/main/scala/utils/SRAMTemplate.scala 126:16]
  always @(posedge clock) begin
    REG <= io_r_0_req_ready & io_r_0_req_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
    if (reset) begin // @[src/main/scala/utils/Hold.scala 23:65]
      r_0_tag <= 19'h0; // @[src/main/scala/utils/Hold.scala 23:65]
    end else if (REG) begin // @[src/main/scala/utils/Hold.scala 23:65]
      r_0_tag <= ram_io_r_resp_data_0_tag; // @[src/main/scala/utils/Hold.scala 23:65]
    end
    if (reset) begin // @[src/main/scala/utils/Hold.scala 23:65]
      r_0_valid <= 1'h0; // @[src/main/scala/utils/Hold.scala 23:65]
    end else if (REG) begin // @[src/main/scala/utils/Hold.scala 23:65]
      r_0_valid <= ram_io_r_resp_data_0_valid; // @[src/main/scala/utils/Hold.scala 23:65]
    end
    if (reset) begin // @[src/main/scala/utils/Hold.scala 23:65]
      r_0_dirty <= 1'h0; // @[src/main/scala/utils/Hold.scala 23:65]
    end else if (REG) begin // @[src/main/scala/utils/Hold.scala 23:65]
      r_0_dirty <= ram_io_r_resp_data_0_dirty; // @[src/main/scala/utils/Hold.scala 23:65]
    end
    if (reset) begin // @[src/main/scala/utils/Hold.scala 23:65]
      r_1_tag <= 19'h0; // @[src/main/scala/utils/Hold.scala 23:65]
    end else if (REG) begin // @[src/main/scala/utils/Hold.scala 23:65]
      r_1_tag <= ram_io_r_resp_data_1_tag; // @[src/main/scala/utils/Hold.scala 23:65]
    end
    if (reset) begin // @[src/main/scala/utils/Hold.scala 23:65]
      r_1_valid <= 1'h0; // @[src/main/scala/utils/Hold.scala 23:65]
    end else if (REG) begin // @[src/main/scala/utils/Hold.scala 23:65]
      r_1_valid <= ram_io_r_resp_data_1_valid; // @[src/main/scala/utils/Hold.scala 23:65]
    end
    if (reset) begin // @[src/main/scala/utils/Hold.scala 23:65]
      r_1_dirty <= 1'h0; // @[src/main/scala/utils/Hold.scala 23:65]
    end else if (REG) begin // @[src/main/scala/utils/Hold.scala 23:65]
      r_1_dirty <= ram_io_r_resp_data_1_dirty; // @[src/main/scala/utils/Hold.scala 23:65]
    end
    if (reset) begin // @[src/main/scala/utils/Hold.scala 23:65]
      r_2_tag <= 19'h0; // @[src/main/scala/utils/Hold.scala 23:65]
    end else if (REG) begin // @[src/main/scala/utils/Hold.scala 23:65]
      r_2_tag <= ram_io_r_resp_data_2_tag; // @[src/main/scala/utils/Hold.scala 23:65]
    end
    if (reset) begin // @[src/main/scala/utils/Hold.scala 23:65]
      r_2_valid <= 1'h0; // @[src/main/scala/utils/Hold.scala 23:65]
    end else if (REG) begin // @[src/main/scala/utils/Hold.scala 23:65]
      r_2_valid <= ram_io_r_resp_data_2_valid; // @[src/main/scala/utils/Hold.scala 23:65]
    end
    if (reset) begin // @[src/main/scala/utils/Hold.scala 23:65]
      r_2_dirty <= 1'h0; // @[src/main/scala/utils/Hold.scala 23:65]
    end else if (REG) begin // @[src/main/scala/utils/Hold.scala 23:65]
      r_2_dirty <= ram_io_r_resp_data_2_dirty; // @[src/main/scala/utils/Hold.scala 23:65]
    end
    if (reset) begin // @[src/main/scala/utils/Hold.scala 23:65]
      r_3_tag <= 19'h0; // @[src/main/scala/utils/Hold.scala 23:65]
    end else if (REG) begin // @[src/main/scala/utils/Hold.scala 23:65]
      r_3_tag <= ram_io_r_resp_data_3_tag; // @[src/main/scala/utils/Hold.scala 23:65]
    end
    if (reset) begin // @[src/main/scala/utils/Hold.scala 23:65]
      r_3_valid <= 1'h0; // @[src/main/scala/utils/Hold.scala 23:65]
    end else if (REG) begin // @[src/main/scala/utils/Hold.scala 23:65]
      r_3_valid <= ram_io_r_resp_data_3_valid; // @[src/main/scala/utils/Hold.scala 23:65]
    end
    if (reset) begin // @[src/main/scala/utils/Hold.scala 23:65]
      r_3_dirty <= 1'h0; // @[src/main/scala/utils/Hold.scala 23:65]
    end else if (REG) begin // @[src/main/scala/utils/Hold.scala 23:65]
      r_3_dirty <= ram_io_r_resp_data_3_dirty; // @[src/main/scala/utils/Hold.scala 23:65]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  REG = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  r_0_tag = _RAND_1[18:0];
  _RAND_2 = {1{`RANDOM}};
  r_0_valid = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  r_0_dirty = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  r_1_tag = _RAND_4[18:0];
  _RAND_5 = {1{`RANDOM}};
  r_1_valid = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  r_1_dirty = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  r_2_tag = _RAND_7[18:0];
  _RAND_8 = {1{`RANDOM}};
  r_2_valid = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  r_2_dirty = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  r_3_tag = _RAND_10[18:0];
  _RAND_11 = {1{`RANDOM}};
  r_3_valid = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  r_3_dirty = _RAND_12[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module SRAMTemplate_2(
  input         clock,
  output        io_r_req_ready, // @[src/main/scala/utils/SRAMTemplate.scala 70:14]
  input         io_r_req_valid, // @[src/main/scala/utils/SRAMTemplate.scala 70:14]
  input  [9:0]  io_r_req_bits_setIdx, // @[src/main/scala/utils/SRAMTemplate.scala 70:14]
  output [63:0] io_r_resp_data_0_data, // @[src/main/scala/utils/SRAMTemplate.scala 70:14]
  output [63:0] io_r_resp_data_1_data, // @[src/main/scala/utils/SRAMTemplate.scala 70:14]
  output [63:0] io_r_resp_data_2_data, // @[src/main/scala/utils/SRAMTemplate.scala 70:14]
  output [63:0] io_r_resp_data_3_data, // @[src/main/scala/utils/SRAMTemplate.scala 70:14]
  input         io_w_req_valid, // @[src/main/scala/utils/SRAMTemplate.scala 70:14]
  input  [9:0]  io_w_req_bits_setIdx, // @[src/main/scala/utils/SRAMTemplate.scala 70:14]
  input  [63:0] io_w_req_bits_data_data, // @[src/main/scala/utils/SRAMTemplate.scala 70:14]
  input  [3:0]  io_w_req_bits_waymask // @[src/main/scala/utils/SRAMTemplate.scala 70:14]
);
`ifdef RANDOMIZE_MEM_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_9;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
`endif // RANDOMIZE_REG_INIT
  reg [63:0] array_0 [0:1023]; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
  wire  array_0_rdata_MPORT_en; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
  wire [9:0] array_0_rdata_MPORT_addr; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
  wire [63:0] array_0_rdata_MPORT_data; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
  wire [63:0] array_0_MPORT_data; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
  wire [9:0] array_0_MPORT_addr; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
  wire  array_0_MPORT_mask; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
  wire  array_0_MPORT_en; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
  reg  array_0_rdata_MPORT_en_pipe_0;
  reg [9:0] array_0_rdata_MPORT_addr_pipe_0;
  reg [63:0] array_1 [0:1023]; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
  wire  array_1_rdata_MPORT_en; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
  wire [9:0] array_1_rdata_MPORT_addr; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
  wire [63:0] array_1_rdata_MPORT_data; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
  wire [63:0] array_1_MPORT_data; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
  wire [9:0] array_1_MPORT_addr; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
  wire  array_1_MPORT_mask; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
  wire  array_1_MPORT_en; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
  reg  array_1_rdata_MPORT_en_pipe_0;
  reg [9:0] array_1_rdata_MPORT_addr_pipe_0;
  reg [63:0] array_2 [0:1023]; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
  wire  array_2_rdata_MPORT_en; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
  wire [9:0] array_2_rdata_MPORT_addr; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
  wire [63:0] array_2_rdata_MPORT_data; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
  wire [63:0] array_2_MPORT_data; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
  wire [9:0] array_2_MPORT_addr; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
  wire  array_2_MPORT_mask; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
  wire  array_2_MPORT_en; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
  reg  array_2_rdata_MPORT_en_pipe_0;
  reg [9:0] array_2_rdata_MPORT_addr_pipe_0;
  reg [63:0] array_3 [0:1023]; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
  wire  array_3_rdata_MPORT_en; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
  wire [9:0] array_3_rdata_MPORT_addr; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
  wire [63:0] array_3_rdata_MPORT_data; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
  wire [63:0] array_3_MPORT_data; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
  wire [9:0] array_3_MPORT_addr; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
  wire  array_3_MPORT_mask; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
  wire  array_3_MPORT_en; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
  reg  array_3_rdata_MPORT_en_pipe_0;
  reg [9:0] array_3_rdata_MPORT_addr_pipe_0;
  wire  _realRen_T = ~io_w_req_valid; // @[src/main/scala/utils/SRAMTemplate.scala 89:41]
  assign array_0_rdata_MPORT_en = array_0_rdata_MPORT_en_pipe_0;
  assign array_0_rdata_MPORT_addr = array_0_rdata_MPORT_addr_pipe_0;
  assign array_0_rdata_MPORT_data = array_0[array_0_rdata_MPORT_addr]; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
  assign array_0_MPORT_data = io_w_req_bits_data_data;
  assign array_0_MPORT_addr = io_w_req_bits_setIdx;
  assign array_0_MPORT_mask = io_w_req_bits_waymask[0];
  assign array_0_MPORT_en = io_w_req_valid;
  assign array_1_rdata_MPORT_en = array_1_rdata_MPORT_en_pipe_0;
  assign array_1_rdata_MPORT_addr = array_1_rdata_MPORT_addr_pipe_0;
  assign array_1_rdata_MPORT_data = array_1[array_1_rdata_MPORT_addr]; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
  assign array_1_MPORT_data = io_w_req_bits_data_data;
  assign array_1_MPORT_addr = io_w_req_bits_setIdx;
  assign array_1_MPORT_mask = io_w_req_bits_waymask[1];
  assign array_1_MPORT_en = io_w_req_valid;
  assign array_2_rdata_MPORT_en = array_2_rdata_MPORT_en_pipe_0;
  assign array_2_rdata_MPORT_addr = array_2_rdata_MPORT_addr_pipe_0;
  assign array_2_rdata_MPORT_data = array_2[array_2_rdata_MPORT_addr]; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
  assign array_2_MPORT_data = io_w_req_bits_data_data;
  assign array_2_MPORT_addr = io_w_req_bits_setIdx;
  assign array_2_MPORT_mask = io_w_req_bits_waymask[2];
  assign array_2_MPORT_en = io_w_req_valid;
  assign array_3_rdata_MPORT_en = array_3_rdata_MPORT_en_pipe_0;
  assign array_3_rdata_MPORT_addr = array_3_rdata_MPORT_addr_pipe_0;
  assign array_3_rdata_MPORT_data = array_3[array_3_rdata_MPORT_addr]; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
  assign array_3_MPORT_data = io_w_req_bits_data_data;
  assign array_3_MPORT_addr = io_w_req_bits_setIdx;
  assign array_3_MPORT_mask = io_w_req_bits_waymask[3];
  assign array_3_MPORT_en = io_w_req_valid;
  assign io_r_req_ready = ~io_w_req_valid; // @[src/main/scala/utils/SRAMTemplate.scala 101:53]
  assign io_r_resp_data_0_data = array_0_rdata_MPORT_data; // @[src/main/scala/utils/SRAMTemplate.scala 98:{78,78}]
  assign io_r_resp_data_1_data = array_1_rdata_MPORT_data; // @[src/main/scala/utils/SRAMTemplate.scala 98:{78,78}]
  assign io_r_resp_data_2_data = array_2_rdata_MPORT_data; // @[src/main/scala/utils/SRAMTemplate.scala 98:{78,78}]
  assign io_r_resp_data_3_data = array_3_rdata_MPORT_data; // @[src/main/scala/utils/SRAMTemplate.scala 98:{78,78}]
  always @(posedge clock) begin
    if (array_0_MPORT_en & array_0_MPORT_mask) begin
      array_0[array_0_MPORT_addr] <= array_0_MPORT_data; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
    end
    array_0_rdata_MPORT_en_pipe_0 <= io_r_req_valid & _realRen_T;
    if (io_r_req_valid & _realRen_T) begin
      array_0_rdata_MPORT_addr_pipe_0 <= io_r_req_bits_setIdx;
    end
    if (array_1_MPORT_en & array_1_MPORT_mask) begin
      array_1[array_1_MPORT_addr] <= array_1_MPORT_data; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
    end
    array_1_rdata_MPORT_en_pipe_0 <= io_r_req_valid & _realRen_T;
    if (io_r_req_valid & _realRen_T) begin
      array_1_rdata_MPORT_addr_pipe_0 <= io_r_req_bits_setIdx;
    end
    if (array_2_MPORT_en & array_2_MPORT_mask) begin
      array_2[array_2_MPORT_addr] <= array_2_MPORT_data; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
    end
    array_2_rdata_MPORT_en_pipe_0 <= io_r_req_valid & _realRen_T;
    if (io_r_req_valid & _realRen_T) begin
      array_2_rdata_MPORT_addr_pipe_0 <= io_r_req_bits_setIdx;
    end
    if (array_3_MPORT_en & array_3_MPORT_mask) begin
      array_3[array_3_MPORT_addr] <= array_3_MPORT_data; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
    end
    array_3_rdata_MPORT_en_pipe_0 <= io_r_req_valid & _realRen_T;
    if (io_r_req_valid & _realRen_T) begin
      array_3_rdata_MPORT_addr_pipe_0 <= io_r_req_bits_setIdx;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {2{`RANDOM}};
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    array_0[initvar] = _RAND_0[63:0];
  _RAND_3 = {2{`RANDOM}};
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    array_1[initvar] = _RAND_3[63:0];
  _RAND_6 = {2{`RANDOM}};
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    array_2[initvar] = _RAND_6[63:0];
  _RAND_9 = {2{`RANDOM}};
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    array_3[initvar] = _RAND_9[63:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  array_0_rdata_MPORT_en_pipe_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  array_0_rdata_MPORT_addr_pipe_0 = _RAND_2[9:0];
  _RAND_4 = {1{`RANDOM}};
  array_1_rdata_MPORT_en_pipe_0 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  array_1_rdata_MPORT_addr_pipe_0 = _RAND_5[9:0];
  _RAND_7 = {1{`RANDOM}};
  array_2_rdata_MPORT_en_pipe_0 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  array_2_rdata_MPORT_addr_pipe_0 = _RAND_8[9:0];
  _RAND_10 = {1{`RANDOM}};
  array_3_rdata_MPORT_en_pipe_0 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  array_3_rdata_MPORT_addr_pipe_0 = _RAND_11[9:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Arbiter_3(
  output       io_in_0_ready, // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
  input        io_in_0_valid, // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
  input  [9:0] io_in_0_bits_setIdx, // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
  output       io_in_1_ready, // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
  input        io_in_1_valid, // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
  input  [9:0] io_in_1_bits_setIdx, // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
  input        io_out_ready, // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
  output       io_out_valid, // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
  output [9:0] io_out_bits_setIdx // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
);
  wire  grant_1 = ~io_in_0_valid; // @[src/main/scala/chisel3/util/Arbiter.scala 45:78]
  assign io_in_0_ready = io_out_ready; // @[src/main/scala/chisel3/util/Arbiter.scala 147:19]
  assign io_in_1_ready = grant_1 & io_out_ready; // @[src/main/scala/chisel3/util/Arbiter.scala 147:19]
  assign io_out_valid = ~grant_1 | io_in_1_valid; // @[src/main/scala/chisel3/util/Arbiter.scala 148:31]
  assign io_out_bits_setIdx = io_in_0_valid ? io_in_0_bits_setIdx : io_in_1_bits_setIdx; // @[src/main/scala/chisel3/util/Arbiter.scala 137:15 139:26 141:19]
endmodule
module SRAMTemplateWithArbiter_1(
  input         clock,
  input         reset,
  output        io_r_0_req_ready, // @[src/main/scala/utils/SRAMTemplate.scala 116:14]
  input         io_r_0_req_valid, // @[src/main/scala/utils/SRAMTemplate.scala 116:14]
  input  [9:0]  io_r_0_req_bits_setIdx, // @[src/main/scala/utils/SRAMTemplate.scala 116:14]
  output [63:0] io_r_0_resp_data_0_data, // @[src/main/scala/utils/SRAMTemplate.scala 116:14]
  output [63:0] io_r_0_resp_data_1_data, // @[src/main/scala/utils/SRAMTemplate.scala 116:14]
  output [63:0] io_r_0_resp_data_2_data, // @[src/main/scala/utils/SRAMTemplate.scala 116:14]
  output [63:0] io_r_0_resp_data_3_data, // @[src/main/scala/utils/SRAMTemplate.scala 116:14]
  output        io_r_1_req_ready, // @[src/main/scala/utils/SRAMTemplate.scala 116:14]
  input         io_r_1_req_valid, // @[src/main/scala/utils/SRAMTemplate.scala 116:14]
  input  [9:0]  io_r_1_req_bits_setIdx, // @[src/main/scala/utils/SRAMTemplate.scala 116:14]
  output [63:0] io_r_1_resp_data_0_data, // @[src/main/scala/utils/SRAMTemplate.scala 116:14]
  output [63:0] io_r_1_resp_data_1_data, // @[src/main/scala/utils/SRAMTemplate.scala 116:14]
  output [63:0] io_r_1_resp_data_2_data, // @[src/main/scala/utils/SRAMTemplate.scala 116:14]
  output [63:0] io_r_1_resp_data_3_data, // @[src/main/scala/utils/SRAMTemplate.scala 116:14]
  input         io_w_req_valid, // @[src/main/scala/utils/SRAMTemplate.scala 116:14]
  input  [9:0]  io_w_req_bits_setIdx, // @[src/main/scala/utils/SRAMTemplate.scala 116:14]
  input  [63:0] io_w_req_bits_data_data, // @[src/main/scala/utils/SRAMTemplate.scala 116:14]
  input  [3:0]  io_w_req_bits_waymask // @[src/main/scala/utils/SRAMTemplate.scala 116:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [63:0] _RAND_9;
`endif // RANDOMIZE_REG_INIT
  wire  ram_clock; // @[src/main/scala/utils/SRAMTemplate.scala 121:19]
  wire  ram_io_r_req_ready; // @[src/main/scala/utils/SRAMTemplate.scala 121:19]
  wire  ram_io_r_req_valid; // @[src/main/scala/utils/SRAMTemplate.scala 121:19]
  wire [9:0] ram_io_r_req_bits_setIdx; // @[src/main/scala/utils/SRAMTemplate.scala 121:19]
  wire [63:0] ram_io_r_resp_data_0_data; // @[src/main/scala/utils/SRAMTemplate.scala 121:19]
  wire [63:0] ram_io_r_resp_data_1_data; // @[src/main/scala/utils/SRAMTemplate.scala 121:19]
  wire [63:0] ram_io_r_resp_data_2_data; // @[src/main/scala/utils/SRAMTemplate.scala 121:19]
  wire [63:0] ram_io_r_resp_data_3_data; // @[src/main/scala/utils/SRAMTemplate.scala 121:19]
  wire  ram_io_w_req_valid; // @[src/main/scala/utils/SRAMTemplate.scala 121:19]
  wire [9:0] ram_io_w_req_bits_setIdx; // @[src/main/scala/utils/SRAMTemplate.scala 121:19]
  wire [63:0] ram_io_w_req_bits_data_data; // @[src/main/scala/utils/SRAMTemplate.scala 121:19]
  wire [3:0] ram_io_w_req_bits_waymask; // @[src/main/scala/utils/SRAMTemplate.scala 121:19]
  wire  readArb_io_in_0_ready; // @[src/main/scala/utils/SRAMTemplate.scala 124:23]
  wire  readArb_io_in_0_valid; // @[src/main/scala/utils/SRAMTemplate.scala 124:23]
  wire [9:0] readArb_io_in_0_bits_setIdx; // @[src/main/scala/utils/SRAMTemplate.scala 124:23]
  wire  readArb_io_in_1_ready; // @[src/main/scala/utils/SRAMTemplate.scala 124:23]
  wire  readArb_io_in_1_valid; // @[src/main/scala/utils/SRAMTemplate.scala 124:23]
  wire [9:0] readArb_io_in_1_bits_setIdx; // @[src/main/scala/utils/SRAMTemplate.scala 124:23]
  wire  readArb_io_out_ready; // @[src/main/scala/utils/SRAMTemplate.scala 124:23]
  wire  readArb_io_out_valid; // @[src/main/scala/utils/SRAMTemplate.scala 124:23]
  wire [9:0] readArb_io_out_bits_setIdx; // @[src/main/scala/utils/SRAMTemplate.scala 124:23]
  reg  REG; // @[src/main/scala/utils/SRAMTemplate.scala 130:58]
  reg [63:0] r__0_data; // @[src/main/scala/utils/Hold.scala 23:65]
  reg [63:0] r__1_data; // @[src/main/scala/utils/Hold.scala 23:65]
  reg [63:0] r__2_data; // @[src/main/scala/utils/Hold.scala 23:65]
  reg [63:0] r__3_data; // @[src/main/scala/utils/Hold.scala 23:65]
  reg  REG_1; // @[src/main/scala/utils/SRAMTemplate.scala 130:58]
  reg [63:0] r_1_0_data; // @[src/main/scala/utils/Hold.scala 23:65]
  reg [63:0] r_1_1_data; // @[src/main/scala/utils/Hold.scala 23:65]
  reg [63:0] r_1_2_data; // @[src/main/scala/utils/Hold.scala 23:65]
  reg [63:0] r_1_3_data; // @[src/main/scala/utils/Hold.scala 23:65]
  SRAMTemplate_2 ram ( // @[src/main/scala/utils/SRAMTemplate.scala 121:19]
    .clock(ram_clock),
    .io_r_req_ready(ram_io_r_req_ready),
    .io_r_req_valid(ram_io_r_req_valid),
    .io_r_req_bits_setIdx(ram_io_r_req_bits_setIdx),
    .io_r_resp_data_0_data(ram_io_r_resp_data_0_data),
    .io_r_resp_data_1_data(ram_io_r_resp_data_1_data),
    .io_r_resp_data_2_data(ram_io_r_resp_data_2_data),
    .io_r_resp_data_3_data(ram_io_r_resp_data_3_data),
    .io_w_req_valid(ram_io_w_req_valid),
    .io_w_req_bits_setIdx(ram_io_w_req_bits_setIdx),
    .io_w_req_bits_data_data(ram_io_w_req_bits_data_data),
    .io_w_req_bits_waymask(ram_io_w_req_bits_waymask)
  );
  Arbiter_3 readArb ( // @[src/main/scala/utils/SRAMTemplate.scala 124:23]
    .io_in_0_ready(readArb_io_in_0_ready),
    .io_in_0_valid(readArb_io_in_0_valid),
    .io_in_0_bits_setIdx(readArb_io_in_0_bits_setIdx),
    .io_in_1_ready(readArb_io_in_1_ready),
    .io_in_1_valid(readArb_io_in_1_valid),
    .io_in_1_bits_setIdx(readArb_io_in_1_bits_setIdx),
    .io_out_ready(readArb_io_out_ready),
    .io_out_valid(readArb_io_out_valid),
    .io_out_bits_setIdx(readArb_io_out_bits_setIdx)
  );
  assign io_r_0_req_ready = readArb_io_in_0_ready; // @[src/main/scala/utils/SRAMTemplate.scala 125:17]
  assign io_r_0_resp_data_0_data = REG ? ram_io_r_resp_data_0_data : r__0_data; // @[src/main/scala/utils/Hold.scala 23:48]
  assign io_r_0_resp_data_1_data = REG ? ram_io_r_resp_data_1_data : r__1_data; // @[src/main/scala/utils/Hold.scala 23:48]
  assign io_r_0_resp_data_2_data = REG ? ram_io_r_resp_data_2_data : r__2_data; // @[src/main/scala/utils/Hold.scala 23:48]
  assign io_r_0_resp_data_3_data = REG ? ram_io_r_resp_data_3_data : r__3_data; // @[src/main/scala/utils/Hold.scala 23:48]
  assign io_r_1_req_ready = readArb_io_in_1_ready; // @[src/main/scala/utils/SRAMTemplate.scala 125:17]
  assign io_r_1_resp_data_0_data = REG_1 ? ram_io_r_resp_data_0_data : r_1_0_data; // @[src/main/scala/utils/Hold.scala 23:48]
  assign io_r_1_resp_data_1_data = REG_1 ? ram_io_r_resp_data_1_data : r_1_1_data; // @[src/main/scala/utils/Hold.scala 23:48]
  assign io_r_1_resp_data_2_data = REG_1 ? ram_io_r_resp_data_2_data : r_1_2_data; // @[src/main/scala/utils/Hold.scala 23:48]
  assign io_r_1_resp_data_3_data = REG_1 ? ram_io_r_resp_data_3_data : r_1_3_data; // @[src/main/scala/utils/Hold.scala 23:48]
  assign ram_clock = clock;
  assign ram_io_r_req_valid = readArb_io_out_valid; // @[src/main/scala/utils/SRAMTemplate.scala 126:16]
  assign ram_io_r_req_bits_setIdx = readArb_io_out_bits_setIdx; // @[src/main/scala/utils/SRAMTemplate.scala 126:16]
  assign ram_io_w_req_valid = io_w_req_valid; // @[src/main/scala/utils/SRAMTemplate.scala 122:12]
  assign ram_io_w_req_bits_setIdx = io_w_req_bits_setIdx; // @[src/main/scala/utils/SRAMTemplate.scala 122:12]
  assign ram_io_w_req_bits_data_data = io_w_req_bits_data_data; // @[src/main/scala/utils/SRAMTemplate.scala 122:12]
  assign ram_io_w_req_bits_waymask = io_w_req_bits_waymask; // @[src/main/scala/utils/SRAMTemplate.scala 122:12]
  assign readArb_io_in_0_valid = io_r_0_req_valid; // @[src/main/scala/utils/SRAMTemplate.scala 125:17]
  assign readArb_io_in_0_bits_setIdx = io_r_0_req_bits_setIdx; // @[src/main/scala/utils/SRAMTemplate.scala 125:17]
  assign readArb_io_in_1_valid = io_r_1_req_valid; // @[src/main/scala/utils/SRAMTemplate.scala 125:17]
  assign readArb_io_in_1_bits_setIdx = io_r_1_req_bits_setIdx; // @[src/main/scala/utils/SRAMTemplate.scala 125:17]
  assign readArb_io_out_ready = ram_io_r_req_ready; // @[src/main/scala/utils/SRAMTemplate.scala 126:16]
  always @(posedge clock) begin
    REG <= io_r_0_req_ready & io_r_0_req_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
    if (reset) begin // @[src/main/scala/utils/Hold.scala 23:65]
      r__0_data <= 64'h0; // @[src/main/scala/utils/Hold.scala 23:65]
    end else if (REG) begin // @[src/main/scala/utils/Hold.scala 23:65]
      r__0_data <= ram_io_r_resp_data_0_data; // @[src/main/scala/utils/Hold.scala 23:65]
    end
    if (reset) begin // @[src/main/scala/utils/Hold.scala 23:65]
      r__1_data <= 64'h0; // @[src/main/scala/utils/Hold.scala 23:65]
    end else if (REG) begin // @[src/main/scala/utils/Hold.scala 23:65]
      r__1_data <= ram_io_r_resp_data_1_data; // @[src/main/scala/utils/Hold.scala 23:65]
    end
    if (reset) begin // @[src/main/scala/utils/Hold.scala 23:65]
      r__2_data <= 64'h0; // @[src/main/scala/utils/Hold.scala 23:65]
    end else if (REG) begin // @[src/main/scala/utils/Hold.scala 23:65]
      r__2_data <= ram_io_r_resp_data_2_data; // @[src/main/scala/utils/Hold.scala 23:65]
    end
    if (reset) begin // @[src/main/scala/utils/Hold.scala 23:65]
      r__3_data <= 64'h0; // @[src/main/scala/utils/Hold.scala 23:65]
    end else if (REG) begin // @[src/main/scala/utils/Hold.scala 23:65]
      r__3_data <= ram_io_r_resp_data_3_data; // @[src/main/scala/utils/Hold.scala 23:65]
    end
    REG_1 <= io_r_1_req_ready & io_r_1_req_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
    if (reset) begin // @[src/main/scala/utils/Hold.scala 23:65]
      r_1_0_data <= 64'h0; // @[src/main/scala/utils/Hold.scala 23:65]
    end else if (REG_1) begin // @[src/main/scala/utils/Hold.scala 23:65]
      r_1_0_data <= ram_io_r_resp_data_0_data; // @[src/main/scala/utils/Hold.scala 23:65]
    end
    if (reset) begin // @[src/main/scala/utils/Hold.scala 23:65]
      r_1_1_data <= 64'h0; // @[src/main/scala/utils/Hold.scala 23:65]
    end else if (REG_1) begin // @[src/main/scala/utils/Hold.scala 23:65]
      r_1_1_data <= ram_io_r_resp_data_1_data; // @[src/main/scala/utils/Hold.scala 23:65]
    end
    if (reset) begin // @[src/main/scala/utils/Hold.scala 23:65]
      r_1_2_data <= 64'h0; // @[src/main/scala/utils/Hold.scala 23:65]
    end else if (REG_1) begin // @[src/main/scala/utils/Hold.scala 23:65]
      r_1_2_data <= ram_io_r_resp_data_2_data; // @[src/main/scala/utils/Hold.scala 23:65]
    end
    if (reset) begin // @[src/main/scala/utils/Hold.scala 23:65]
      r_1_3_data <= 64'h0; // @[src/main/scala/utils/Hold.scala 23:65]
    end else if (REG_1) begin // @[src/main/scala/utils/Hold.scala 23:65]
      r_1_3_data <= ram_io_r_resp_data_3_data; // @[src/main/scala/utils/Hold.scala 23:65]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  REG = _RAND_0[0:0];
  _RAND_1 = {2{`RANDOM}};
  r__0_data = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  r__1_data = _RAND_2[63:0];
  _RAND_3 = {2{`RANDOM}};
  r__2_data = _RAND_3[63:0];
  _RAND_4 = {2{`RANDOM}};
  r__3_data = _RAND_4[63:0];
  _RAND_5 = {1{`RANDOM}};
  REG_1 = _RAND_5[0:0];
  _RAND_6 = {2{`RANDOM}};
  r_1_0_data = _RAND_6[63:0];
  _RAND_7 = {2{`RANDOM}};
  r_1_1_data = _RAND_7[63:0];
  _RAND_8 = {2{`RANDOM}};
  r_1_2_data = _RAND_8[63:0];
  _RAND_9 = {2{`RANDOM}};
  r_1_3_data = _RAND_9[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Arbiter_4(
  output        io_in_0_ready, // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
  input         io_in_0_valid, // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
  input  [31:0] io_in_0_bits_addr, // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
  input  [86:0] io_in_0_bits_user, // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
  input         io_out_ready, // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
  output        io_out_valid, // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
  output [31:0] io_out_bits_addr, // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
  output [86:0] io_out_bits_user // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
);
  assign io_in_0_ready = io_out_ready; // @[src/main/scala/chisel3/util/Arbiter.scala 147:19]
  assign io_out_valid = io_in_0_valid; // @[src/main/scala/chisel3/util/Arbiter.scala 148:31]
  assign io_out_bits_addr = io_in_0_bits_addr; // @[src/main/scala/chisel3/util/Arbiter.scala 137:15]
  assign io_out_bits_user = io_in_0_bits_user; // @[src/main/scala/chisel3/util/Arbiter.scala 137:15]
endmodule
module Cache(
  input         clock,
  input         reset,
  output        io_in_req_ready, // @[src/main/scala/nutcore/mem/Cache.scala 122:14]
  input         io_in_req_valid, // @[src/main/scala/nutcore/mem/Cache.scala 122:14]
  input  [31:0] io_in_req_bits_addr, // @[src/main/scala/nutcore/mem/Cache.scala 122:14]
  input  [86:0] io_in_req_bits_user, // @[src/main/scala/nutcore/mem/Cache.scala 122:14]
  input         io_in_resp_ready, // @[src/main/scala/nutcore/mem/Cache.scala 122:14]
  output        io_in_resp_valid, // @[src/main/scala/nutcore/mem/Cache.scala 122:14]
  output [63:0] io_in_resp_bits_rdata, // @[src/main/scala/nutcore/mem/Cache.scala 122:14]
  output [86:0] io_in_resp_bits_user, // @[src/main/scala/nutcore/mem/Cache.scala 122:14]
  input  [1:0]  io_flush, // @[src/main/scala/nutcore/mem/Cache.scala 122:14]
  input         io_out_mem_req_ready, // @[src/main/scala/nutcore/mem/Cache.scala 122:14]
  output        io_out_mem_req_valid, // @[src/main/scala/nutcore/mem/Cache.scala 122:14]
  output [31:0] io_out_mem_req_bits_addr, // @[src/main/scala/nutcore/mem/Cache.scala 122:14]
  output [3:0]  io_out_mem_req_bits_cmd, // @[src/main/scala/nutcore/mem/Cache.scala 122:14]
  output [63:0] io_out_mem_req_bits_wdata, // @[src/main/scala/nutcore/mem/Cache.scala 122:14]
  input         io_out_mem_resp_valid, // @[src/main/scala/nutcore/mem/Cache.scala 122:14]
  input  [3:0]  io_out_mem_resp_bits_cmd, // @[src/main/scala/nutcore/mem/Cache.scala 122:14]
  input  [63:0] io_out_mem_resp_bits_rdata, // @[src/main/scala/nutcore/mem/Cache.scala 122:14]
  input         io_mmio_req_ready, // @[src/main/scala/nutcore/mem/Cache.scala 122:14]
  output        io_mmio_req_valid, // @[src/main/scala/nutcore/mem/Cache.scala 122:14]
  output [31:0] io_mmio_req_bits_addr, // @[src/main/scala/nutcore/mem/Cache.scala 122:14]
  input         io_mmio_resp_valid, // @[src/main/scala/nutcore/mem/Cache.scala 122:14]
  input  [63:0] io_mmio_resp_bits_rdata, // @[src/main/scala/nutcore/mem/Cache.scala 122:14]
  output        io_empty, // @[src/main/scala/nutcore/mem/Cache.scala 122:14]
  input         DISPLAY_ENABLE,
  input         MOUFlushICache
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [95:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [95:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [63:0] _RAND_18;
  reg [63:0] _RAND_19;
  reg [63:0] _RAND_20;
  reg [63:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [63:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [63:0] _RAND_28;
  reg [63:0] _RAND_29;
  reg [63:0] _RAND_30;
  reg [63:0] _RAND_31;
  reg [63:0] _RAND_32;
`endif // RANDOMIZE_REG_INIT
  wire  s1_clock; // @[src/main/scala/nutcore/mem/Cache.scala 480:18]
  wire  s1_reset; // @[src/main/scala/nutcore/mem/Cache.scala 480:18]
  wire  s1_io_in_ready; // @[src/main/scala/nutcore/mem/Cache.scala 480:18]
  wire  s1_io_in_valid; // @[src/main/scala/nutcore/mem/Cache.scala 480:18]
  wire [31:0] s1_io_in_bits_addr; // @[src/main/scala/nutcore/mem/Cache.scala 480:18]
  wire [2:0] s1_io_in_bits_size; // @[src/main/scala/nutcore/mem/Cache.scala 480:18]
  wire [3:0] s1_io_in_bits_cmd; // @[src/main/scala/nutcore/mem/Cache.scala 480:18]
  wire [7:0] s1_io_in_bits_wmask; // @[src/main/scala/nutcore/mem/Cache.scala 480:18]
  wire [63:0] s1_io_in_bits_wdata; // @[src/main/scala/nutcore/mem/Cache.scala 480:18]
  wire [86:0] s1_io_in_bits_user; // @[src/main/scala/nutcore/mem/Cache.scala 480:18]
  wire  s1_io_out_ready; // @[src/main/scala/nutcore/mem/Cache.scala 480:18]
  wire  s1_io_out_valid; // @[src/main/scala/nutcore/mem/Cache.scala 480:18]
  wire [31:0] s1_io_out_bits_req_addr; // @[src/main/scala/nutcore/mem/Cache.scala 480:18]
  wire [86:0] s1_io_out_bits_req_user; // @[src/main/scala/nutcore/mem/Cache.scala 480:18]
  wire  s1_io_metaReadBus_req_ready; // @[src/main/scala/nutcore/mem/Cache.scala 480:18]
  wire  s1_io_metaReadBus_req_valid; // @[src/main/scala/nutcore/mem/Cache.scala 480:18]
  wire [6:0] s1_io_metaReadBus_req_bits_setIdx; // @[src/main/scala/nutcore/mem/Cache.scala 480:18]
  wire [18:0] s1_io_metaReadBus_resp_data_0_tag; // @[src/main/scala/nutcore/mem/Cache.scala 480:18]
  wire  s1_io_metaReadBus_resp_data_0_valid; // @[src/main/scala/nutcore/mem/Cache.scala 480:18]
  wire  s1_io_metaReadBus_resp_data_0_dirty; // @[src/main/scala/nutcore/mem/Cache.scala 480:18]
  wire [18:0] s1_io_metaReadBus_resp_data_1_tag; // @[src/main/scala/nutcore/mem/Cache.scala 480:18]
  wire  s1_io_metaReadBus_resp_data_1_valid; // @[src/main/scala/nutcore/mem/Cache.scala 480:18]
  wire  s1_io_metaReadBus_resp_data_1_dirty; // @[src/main/scala/nutcore/mem/Cache.scala 480:18]
  wire [18:0] s1_io_metaReadBus_resp_data_2_tag; // @[src/main/scala/nutcore/mem/Cache.scala 480:18]
  wire  s1_io_metaReadBus_resp_data_2_valid; // @[src/main/scala/nutcore/mem/Cache.scala 480:18]
  wire  s1_io_metaReadBus_resp_data_2_dirty; // @[src/main/scala/nutcore/mem/Cache.scala 480:18]
  wire [18:0] s1_io_metaReadBus_resp_data_3_tag; // @[src/main/scala/nutcore/mem/Cache.scala 480:18]
  wire  s1_io_metaReadBus_resp_data_3_valid; // @[src/main/scala/nutcore/mem/Cache.scala 480:18]
  wire  s1_io_metaReadBus_resp_data_3_dirty; // @[src/main/scala/nutcore/mem/Cache.scala 480:18]
  wire  s1_io_dataReadBus_req_ready; // @[src/main/scala/nutcore/mem/Cache.scala 480:18]
  wire  s1_io_dataReadBus_req_valid; // @[src/main/scala/nutcore/mem/Cache.scala 480:18]
  wire [9:0] s1_io_dataReadBus_req_bits_setIdx; // @[src/main/scala/nutcore/mem/Cache.scala 480:18]
  wire [63:0] s1_io_dataReadBus_resp_data_0_data; // @[src/main/scala/nutcore/mem/Cache.scala 480:18]
  wire [63:0] s1_io_dataReadBus_resp_data_1_data; // @[src/main/scala/nutcore/mem/Cache.scala 480:18]
  wire [63:0] s1_io_dataReadBus_resp_data_2_data; // @[src/main/scala/nutcore/mem/Cache.scala 480:18]
  wire [63:0] s1_io_dataReadBus_resp_data_3_data; // @[src/main/scala/nutcore/mem/Cache.scala 480:18]
  wire  s1_DISPLAY_ENABLE; // @[src/main/scala/nutcore/mem/Cache.scala 480:18]
  wire  s2_clock; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire  s2_reset; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire  s2_io_in_ready; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire  s2_io_in_valid; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire [31:0] s2_io_in_bits_req_addr; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire [2:0] s2_io_in_bits_req_size; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire [3:0] s2_io_in_bits_req_cmd; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire [7:0] s2_io_in_bits_req_wmask; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire [63:0] s2_io_in_bits_req_wdata; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire [86:0] s2_io_in_bits_req_user; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire  s2_io_out_ready; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire  s2_io_out_valid; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire [31:0] s2_io_out_bits_req_addr; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire [86:0] s2_io_out_bits_req_user; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire [18:0] s2_io_out_bits_metas_0_tag; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire  s2_io_out_bits_metas_0_valid; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire  s2_io_out_bits_metas_0_dirty; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire [18:0] s2_io_out_bits_metas_1_tag; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire  s2_io_out_bits_metas_1_valid; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire  s2_io_out_bits_metas_1_dirty; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire [18:0] s2_io_out_bits_metas_2_tag; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire  s2_io_out_bits_metas_2_valid; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire  s2_io_out_bits_metas_2_dirty; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire [18:0] s2_io_out_bits_metas_3_tag; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire  s2_io_out_bits_metas_3_valid; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire  s2_io_out_bits_metas_3_dirty; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire [63:0] s2_io_out_bits_datas_0_data; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire [63:0] s2_io_out_bits_datas_1_data; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire [63:0] s2_io_out_bits_datas_2_data; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire [63:0] s2_io_out_bits_datas_3_data; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire  s2_io_out_bits_hit; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire [3:0] s2_io_out_bits_waymask; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire  s2_io_out_bits_mmio; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire  s2_io_out_bits_isForwardData; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire [63:0] s2_io_out_bits_forwardData_data_data; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire [3:0] s2_io_out_bits_forwardData_waymask; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire [18:0] s2_io_metaReadResp_0_tag; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire  s2_io_metaReadResp_0_valid; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire  s2_io_metaReadResp_0_dirty; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire [18:0] s2_io_metaReadResp_1_tag; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire  s2_io_metaReadResp_1_valid; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire  s2_io_metaReadResp_1_dirty; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire [18:0] s2_io_metaReadResp_2_tag; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire  s2_io_metaReadResp_2_valid; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire  s2_io_metaReadResp_2_dirty; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire [18:0] s2_io_metaReadResp_3_tag; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire  s2_io_metaReadResp_3_valid; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire  s2_io_metaReadResp_3_dirty; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire [63:0] s2_io_dataReadResp_0_data; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire [63:0] s2_io_dataReadResp_1_data; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire [63:0] s2_io_dataReadResp_2_data; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire [63:0] s2_io_dataReadResp_3_data; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire  s2_io_metaWriteBus_req_valid; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire [6:0] s2_io_metaWriteBus_req_bits_setIdx; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire [18:0] s2_io_metaWriteBus_req_bits_data_tag; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire  s2_io_metaWriteBus_req_bits_data_dirty; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire [3:0] s2_io_metaWriteBus_req_bits_waymask; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire  s2_io_dataWriteBus_req_valid; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire [9:0] s2_io_dataWriteBus_req_bits_setIdx; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire [63:0] s2_io_dataWriteBus_req_bits_data_data; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire [3:0] s2_io_dataWriteBus_req_bits_waymask; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire  s2_DISPLAY_ENABLE; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire  s3_clock; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire  s3_reset; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire  s3_io_in_ready; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire  s3_io_in_valid; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire [31:0] s3_io_in_bits_req_addr; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire [2:0] s3_io_in_bits_req_size; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire [3:0] s3_io_in_bits_req_cmd; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire [7:0] s3_io_in_bits_req_wmask; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire [63:0] s3_io_in_bits_req_wdata; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire [86:0] s3_io_in_bits_req_user; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire [18:0] s3_io_in_bits_metas_0_tag; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire  s3_io_in_bits_metas_0_valid; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire  s3_io_in_bits_metas_0_dirty; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire [18:0] s3_io_in_bits_metas_1_tag; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire  s3_io_in_bits_metas_1_valid; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire  s3_io_in_bits_metas_1_dirty; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire [18:0] s3_io_in_bits_metas_2_tag; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire  s3_io_in_bits_metas_2_valid; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire  s3_io_in_bits_metas_2_dirty; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire [18:0] s3_io_in_bits_metas_3_tag; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire  s3_io_in_bits_metas_3_valid; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire  s3_io_in_bits_metas_3_dirty; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire [63:0] s3_io_in_bits_datas_0_data; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire [63:0] s3_io_in_bits_datas_1_data; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire [63:0] s3_io_in_bits_datas_2_data; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire [63:0] s3_io_in_bits_datas_3_data; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire  s3_io_in_bits_hit; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire [3:0] s3_io_in_bits_waymask; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire  s3_io_in_bits_mmio; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire  s3_io_in_bits_isForwardData; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire [63:0] s3_io_in_bits_forwardData_data_data; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire [3:0] s3_io_in_bits_forwardData_waymask; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire  s3_io_out_ready; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire  s3_io_out_valid; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire [3:0] s3_io_out_bits_cmd; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire [63:0] s3_io_out_bits_rdata; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire [86:0] s3_io_out_bits_user; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire  s3_io_isFinish; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire  s3_io_flush; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire  s3_io_dataReadBus_req_ready; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire  s3_io_dataReadBus_req_valid; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire [9:0] s3_io_dataReadBus_req_bits_setIdx; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire [63:0] s3_io_dataReadBus_resp_data_0_data; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire [63:0] s3_io_dataReadBus_resp_data_1_data; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire [63:0] s3_io_dataReadBus_resp_data_2_data; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire [63:0] s3_io_dataReadBus_resp_data_3_data; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire  s3_io_dataWriteBus_req_valid; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire [9:0] s3_io_dataWriteBus_req_bits_setIdx; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire [63:0] s3_io_dataWriteBus_req_bits_data_data; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire [3:0] s3_io_dataWriteBus_req_bits_waymask; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire  s3_io_metaWriteBus_req_valid; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire [6:0] s3_io_metaWriteBus_req_bits_setIdx; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire [18:0] s3_io_metaWriteBus_req_bits_data_tag; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire  s3_io_metaWriteBus_req_bits_data_valid; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire  s3_io_metaWriteBus_req_bits_data_dirty; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire [3:0] s3_io_metaWriteBus_req_bits_waymask; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire  s3_io_mem_req_ready; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire  s3_io_mem_req_valid; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire [31:0] s3_io_mem_req_bits_addr; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire [2:0] s3_io_mem_req_bits_size; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire [3:0] s3_io_mem_req_bits_cmd; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire [7:0] s3_io_mem_req_bits_wmask; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire [63:0] s3_io_mem_req_bits_wdata; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire  s3_io_mem_resp_ready; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire  s3_io_mem_resp_valid; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire [3:0] s3_io_mem_resp_bits_cmd; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire [63:0] s3_io_mem_resp_bits_rdata; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire  s3_io_mmio_req_ready; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire  s3_io_mmio_req_valid; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire [31:0] s3_io_mmio_req_bits_addr; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire  s3_io_mmio_resp_ready; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire  s3_io_mmio_resp_valid; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire [63:0] s3_io_mmio_resp_bits_rdata; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire  s3_io_cohResp_valid; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire  s3_DISPLAY_ENABLE; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire  metaArray_clock; // @[src/main/scala/nutcore/mem/Cache.scala 483:25]
  wire  metaArray_reset; // @[src/main/scala/nutcore/mem/Cache.scala 483:25]
  wire  metaArray_io_r_0_req_ready; // @[src/main/scala/nutcore/mem/Cache.scala 483:25]
  wire  metaArray_io_r_0_req_valid; // @[src/main/scala/nutcore/mem/Cache.scala 483:25]
  wire [6:0] metaArray_io_r_0_req_bits_setIdx; // @[src/main/scala/nutcore/mem/Cache.scala 483:25]
  wire [18:0] metaArray_io_r_0_resp_data_0_tag; // @[src/main/scala/nutcore/mem/Cache.scala 483:25]
  wire  metaArray_io_r_0_resp_data_0_valid; // @[src/main/scala/nutcore/mem/Cache.scala 483:25]
  wire  metaArray_io_r_0_resp_data_0_dirty; // @[src/main/scala/nutcore/mem/Cache.scala 483:25]
  wire [18:0] metaArray_io_r_0_resp_data_1_tag; // @[src/main/scala/nutcore/mem/Cache.scala 483:25]
  wire  metaArray_io_r_0_resp_data_1_valid; // @[src/main/scala/nutcore/mem/Cache.scala 483:25]
  wire  metaArray_io_r_0_resp_data_1_dirty; // @[src/main/scala/nutcore/mem/Cache.scala 483:25]
  wire [18:0] metaArray_io_r_0_resp_data_2_tag; // @[src/main/scala/nutcore/mem/Cache.scala 483:25]
  wire  metaArray_io_r_0_resp_data_2_valid; // @[src/main/scala/nutcore/mem/Cache.scala 483:25]
  wire  metaArray_io_r_0_resp_data_2_dirty; // @[src/main/scala/nutcore/mem/Cache.scala 483:25]
  wire [18:0] metaArray_io_r_0_resp_data_3_tag; // @[src/main/scala/nutcore/mem/Cache.scala 483:25]
  wire  metaArray_io_r_0_resp_data_3_valid; // @[src/main/scala/nutcore/mem/Cache.scala 483:25]
  wire  metaArray_io_r_0_resp_data_3_dirty; // @[src/main/scala/nutcore/mem/Cache.scala 483:25]
  wire  metaArray_io_w_req_valid; // @[src/main/scala/nutcore/mem/Cache.scala 483:25]
  wire [6:0] metaArray_io_w_req_bits_setIdx; // @[src/main/scala/nutcore/mem/Cache.scala 483:25]
  wire [18:0] metaArray_io_w_req_bits_data_tag; // @[src/main/scala/nutcore/mem/Cache.scala 483:25]
  wire  metaArray_io_w_req_bits_data_dirty; // @[src/main/scala/nutcore/mem/Cache.scala 483:25]
  wire [3:0] metaArray_io_w_req_bits_waymask; // @[src/main/scala/nutcore/mem/Cache.scala 483:25]
  wire  dataArray_clock; // @[src/main/scala/nutcore/mem/Cache.scala 484:25]
  wire  dataArray_reset; // @[src/main/scala/nutcore/mem/Cache.scala 484:25]
  wire  dataArray_io_r_0_req_ready; // @[src/main/scala/nutcore/mem/Cache.scala 484:25]
  wire  dataArray_io_r_0_req_valid; // @[src/main/scala/nutcore/mem/Cache.scala 484:25]
  wire [9:0] dataArray_io_r_0_req_bits_setIdx; // @[src/main/scala/nutcore/mem/Cache.scala 484:25]
  wire [63:0] dataArray_io_r_0_resp_data_0_data; // @[src/main/scala/nutcore/mem/Cache.scala 484:25]
  wire [63:0] dataArray_io_r_0_resp_data_1_data; // @[src/main/scala/nutcore/mem/Cache.scala 484:25]
  wire [63:0] dataArray_io_r_0_resp_data_2_data; // @[src/main/scala/nutcore/mem/Cache.scala 484:25]
  wire [63:0] dataArray_io_r_0_resp_data_3_data; // @[src/main/scala/nutcore/mem/Cache.scala 484:25]
  wire  dataArray_io_r_1_req_ready; // @[src/main/scala/nutcore/mem/Cache.scala 484:25]
  wire  dataArray_io_r_1_req_valid; // @[src/main/scala/nutcore/mem/Cache.scala 484:25]
  wire [9:0] dataArray_io_r_1_req_bits_setIdx; // @[src/main/scala/nutcore/mem/Cache.scala 484:25]
  wire [63:0] dataArray_io_r_1_resp_data_0_data; // @[src/main/scala/nutcore/mem/Cache.scala 484:25]
  wire [63:0] dataArray_io_r_1_resp_data_1_data; // @[src/main/scala/nutcore/mem/Cache.scala 484:25]
  wire [63:0] dataArray_io_r_1_resp_data_2_data; // @[src/main/scala/nutcore/mem/Cache.scala 484:25]
  wire [63:0] dataArray_io_r_1_resp_data_3_data; // @[src/main/scala/nutcore/mem/Cache.scala 484:25]
  wire  dataArray_io_w_req_valid; // @[src/main/scala/nutcore/mem/Cache.scala 484:25]
  wire [9:0] dataArray_io_w_req_bits_setIdx; // @[src/main/scala/nutcore/mem/Cache.scala 484:25]
  wire [63:0] dataArray_io_w_req_bits_data_data; // @[src/main/scala/nutcore/mem/Cache.scala 484:25]
  wire [3:0] dataArray_io_w_req_bits_waymask; // @[src/main/scala/nutcore/mem/Cache.scala 484:25]
  wire  arb_io_in_0_ready; // @[src/main/scala/nutcore/mem/Cache.scala 493:19]
  wire  arb_io_in_0_valid; // @[src/main/scala/nutcore/mem/Cache.scala 493:19]
  wire [31:0] arb_io_in_0_bits_addr; // @[src/main/scala/nutcore/mem/Cache.scala 493:19]
  wire [86:0] arb_io_in_0_bits_user; // @[src/main/scala/nutcore/mem/Cache.scala 493:19]
  wire  arb_io_out_ready; // @[src/main/scala/nutcore/mem/Cache.scala 493:19]
  wire  arb_io_out_valid; // @[src/main/scala/nutcore/mem/Cache.scala 493:19]
  wire [31:0] arb_io_out_bits_addr; // @[src/main/scala/nutcore/mem/Cache.scala 493:19]
  wire [86:0] arb_io_out_bits_user; // @[src/main/scala/nutcore/mem/Cache.scala 493:19]
  wire  _T = s2_io_out_ready & s2_io_out_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  reg  valid; // @[src/main/scala/utils/Pipeline.scala 24:24]
  wire  _GEN_0 = _T ? 1'h0 : valid; // @[src/main/scala/utils/Pipeline.scala 24:24 25:{25,33}]
  wire  _T_2 = s1_io_out_valid & s2_io_in_ready; // @[src/main/scala/utils/Pipeline.scala 26:22]
  wire  _GEN_1 = s1_io_out_valid & s2_io_in_ready | _GEN_0; // @[src/main/scala/utils/Pipeline.scala 26:{38,46}]
  reg [31:0] s2_io_in_bits_r_req_addr; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg [86:0] s2_io_in_bits_r_req_user; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg  valid_1; // @[src/main/scala/utils/Pipeline.scala 24:24]
  wire  _GEN_9 = s3_io_isFinish ? 1'h0 : valid_1; // @[src/main/scala/utils/Pipeline.scala 24:24 25:{25,33}]
  wire  _T_4 = s2_io_out_valid & s3_io_in_ready; // @[src/main/scala/utils/Pipeline.scala 26:22]
  wire  _GEN_10 = s2_io_out_valid & s3_io_in_ready | _GEN_9; // @[src/main/scala/utils/Pipeline.scala 26:{38,46}]
  reg [31:0] s3_io_in_bits_r_req_addr; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg [86:0] s3_io_in_bits_r_req_user; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg [18:0] s3_io_in_bits_r_metas_0_tag; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg  s3_io_in_bits_r_metas_0_valid; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg  s3_io_in_bits_r_metas_0_dirty; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg [18:0] s3_io_in_bits_r_metas_1_tag; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg  s3_io_in_bits_r_metas_1_valid; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg  s3_io_in_bits_r_metas_1_dirty; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg [18:0] s3_io_in_bits_r_metas_2_tag; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg  s3_io_in_bits_r_metas_2_valid; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg  s3_io_in_bits_r_metas_2_dirty; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg [18:0] s3_io_in_bits_r_metas_3_tag; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg  s3_io_in_bits_r_metas_3_valid; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg  s3_io_in_bits_r_metas_3_dirty; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg [63:0] s3_io_in_bits_r_datas_0_data; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg [63:0] s3_io_in_bits_r_datas_1_data; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg [63:0] s3_io_in_bits_r_datas_2_data; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg [63:0] s3_io_in_bits_r_datas_3_data; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg  s3_io_in_bits_r_hit; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg [3:0] s3_io_in_bits_r_waymask; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg  s3_io_in_bits_r_mmio; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg  s3_io_in_bits_r_isForwardData; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg [63:0] s3_io_in_bits_r_forwardData_data_data; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg [3:0] s3_io_in_bits_r_forwardData_waymask; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg [63:0] c; // @[src/main/scala/utils/GTimer.scala 24:20]
  wire [63:0] _c_T_1 = c + 64'h1; // @[src/main/scala/utils/GTimer.scala 25:12]
  wire  _T_7 = ~reset; // @[src/main/scala/utils/Debug.scala 56:24]
  reg [63:0] c_1; // @[src/main/scala/utils/GTimer.scala 24:20]
  wire [63:0] _c_T_3 = c_1 + 64'h1; // @[src/main/scala/utils/GTimer.scala 25:12]
  reg [63:0] c_2; // @[src/main/scala/utils/GTimer.scala 24:20]
  wire [63:0] _c_T_5 = c_2 + 64'h1; // @[src/main/scala/utils/GTimer.scala 25:12]
  reg [63:0] c_3; // @[src/main/scala/utils/GTimer.scala 24:20]
  wire [63:0] _c_T_7 = c_3 + 64'h1; // @[src/main/scala/utils/GTimer.scala 25:12]
  reg [63:0] c_4; // @[src/main/scala/utils/GTimer.scala 24:20]
  wire [63:0] _c_T_9 = c_4 + 64'h1; // @[src/main/scala/utils/GTimer.scala 25:12]
  wire  _GEN_41 = s1_io_in_valid & DISPLAY_ENABLE; // @[src/main/scala/utils/Debug.scala 56:24]
  wire  _GEN_43 = s2_io_in_valid & DISPLAY_ENABLE; // @[src/main/scala/utils/Debug.scala 56:24]
  wire  _GEN_45 = s3_io_in_valid & DISPLAY_ENABLE; // @[src/main/scala/utils/Debug.scala 56:24]
  CacheStage1 s1 ( // @[src/main/scala/nutcore/mem/Cache.scala 480:18]
    .clock(s1_clock),
    .reset(s1_reset),
    .io_in_ready(s1_io_in_ready),
    .io_in_valid(s1_io_in_valid),
    .io_in_bits_addr(s1_io_in_bits_addr),
    .io_in_bits_size(s1_io_in_bits_size),
    .io_in_bits_cmd(s1_io_in_bits_cmd),
    .io_in_bits_wmask(s1_io_in_bits_wmask),
    .io_in_bits_wdata(s1_io_in_bits_wdata),
    .io_in_bits_user(s1_io_in_bits_user),
    .io_out_ready(s1_io_out_ready),
    .io_out_valid(s1_io_out_valid),
    .io_out_bits_req_addr(s1_io_out_bits_req_addr),
    .io_out_bits_req_user(s1_io_out_bits_req_user),
    .io_metaReadBus_req_ready(s1_io_metaReadBus_req_ready),
    .io_metaReadBus_req_valid(s1_io_metaReadBus_req_valid),
    .io_metaReadBus_req_bits_setIdx(s1_io_metaReadBus_req_bits_setIdx),
    .io_metaReadBus_resp_data_0_tag(s1_io_metaReadBus_resp_data_0_tag),
    .io_metaReadBus_resp_data_0_valid(s1_io_metaReadBus_resp_data_0_valid),
    .io_metaReadBus_resp_data_0_dirty(s1_io_metaReadBus_resp_data_0_dirty),
    .io_metaReadBus_resp_data_1_tag(s1_io_metaReadBus_resp_data_1_tag),
    .io_metaReadBus_resp_data_1_valid(s1_io_metaReadBus_resp_data_1_valid),
    .io_metaReadBus_resp_data_1_dirty(s1_io_metaReadBus_resp_data_1_dirty),
    .io_metaReadBus_resp_data_2_tag(s1_io_metaReadBus_resp_data_2_tag),
    .io_metaReadBus_resp_data_2_valid(s1_io_metaReadBus_resp_data_2_valid),
    .io_metaReadBus_resp_data_2_dirty(s1_io_metaReadBus_resp_data_2_dirty),
    .io_metaReadBus_resp_data_3_tag(s1_io_metaReadBus_resp_data_3_tag),
    .io_metaReadBus_resp_data_3_valid(s1_io_metaReadBus_resp_data_3_valid),
    .io_metaReadBus_resp_data_3_dirty(s1_io_metaReadBus_resp_data_3_dirty),
    .io_dataReadBus_req_ready(s1_io_dataReadBus_req_ready),
    .io_dataReadBus_req_valid(s1_io_dataReadBus_req_valid),
    .io_dataReadBus_req_bits_setIdx(s1_io_dataReadBus_req_bits_setIdx),
    .io_dataReadBus_resp_data_0_data(s1_io_dataReadBus_resp_data_0_data),
    .io_dataReadBus_resp_data_1_data(s1_io_dataReadBus_resp_data_1_data),
    .io_dataReadBus_resp_data_2_data(s1_io_dataReadBus_resp_data_2_data),
    .io_dataReadBus_resp_data_3_data(s1_io_dataReadBus_resp_data_3_data),
    .DISPLAY_ENABLE(s1_DISPLAY_ENABLE)
  );
  CacheStage2 s2 ( // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
    .clock(s2_clock),
    .reset(s2_reset),
    .io_in_ready(s2_io_in_ready),
    .io_in_valid(s2_io_in_valid),
    .io_in_bits_req_addr(s2_io_in_bits_req_addr),
    .io_in_bits_req_size(s2_io_in_bits_req_size),
    .io_in_bits_req_cmd(s2_io_in_bits_req_cmd),
    .io_in_bits_req_wmask(s2_io_in_bits_req_wmask),
    .io_in_bits_req_wdata(s2_io_in_bits_req_wdata),
    .io_in_bits_req_user(s2_io_in_bits_req_user),
    .io_out_ready(s2_io_out_ready),
    .io_out_valid(s2_io_out_valid),
    .io_out_bits_req_addr(s2_io_out_bits_req_addr),
    .io_out_bits_req_user(s2_io_out_bits_req_user),
    .io_out_bits_metas_0_tag(s2_io_out_bits_metas_0_tag),
    .io_out_bits_metas_0_valid(s2_io_out_bits_metas_0_valid),
    .io_out_bits_metas_0_dirty(s2_io_out_bits_metas_0_dirty),
    .io_out_bits_metas_1_tag(s2_io_out_bits_metas_1_tag),
    .io_out_bits_metas_1_valid(s2_io_out_bits_metas_1_valid),
    .io_out_bits_metas_1_dirty(s2_io_out_bits_metas_1_dirty),
    .io_out_bits_metas_2_tag(s2_io_out_bits_metas_2_tag),
    .io_out_bits_metas_2_valid(s2_io_out_bits_metas_2_valid),
    .io_out_bits_metas_2_dirty(s2_io_out_bits_metas_2_dirty),
    .io_out_bits_metas_3_tag(s2_io_out_bits_metas_3_tag),
    .io_out_bits_metas_3_valid(s2_io_out_bits_metas_3_valid),
    .io_out_bits_metas_3_dirty(s2_io_out_bits_metas_3_dirty),
    .io_out_bits_datas_0_data(s2_io_out_bits_datas_0_data),
    .io_out_bits_datas_1_data(s2_io_out_bits_datas_1_data),
    .io_out_bits_datas_2_data(s2_io_out_bits_datas_2_data),
    .io_out_bits_datas_3_data(s2_io_out_bits_datas_3_data),
    .io_out_bits_hit(s2_io_out_bits_hit),
    .io_out_bits_waymask(s2_io_out_bits_waymask),
    .io_out_bits_mmio(s2_io_out_bits_mmio),
    .io_out_bits_isForwardData(s2_io_out_bits_isForwardData),
    .io_out_bits_forwardData_data_data(s2_io_out_bits_forwardData_data_data),
    .io_out_bits_forwardData_waymask(s2_io_out_bits_forwardData_waymask),
    .io_metaReadResp_0_tag(s2_io_metaReadResp_0_tag),
    .io_metaReadResp_0_valid(s2_io_metaReadResp_0_valid),
    .io_metaReadResp_0_dirty(s2_io_metaReadResp_0_dirty),
    .io_metaReadResp_1_tag(s2_io_metaReadResp_1_tag),
    .io_metaReadResp_1_valid(s2_io_metaReadResp_1_valid),
    .io_metaReadResp_1_dirty(s2_io_metaReadResp_1_dirty),
    .io_metaReadResp_2_tag(s2_io_metaReadResp_2_tag),
    .io_metaReadResp_2_valid(s2_io_metaReadResp_2_valid),
    .io_metaReadResp_2_dirty(s2_io_metaReadResp_2_dirty),
    .io_metaReadResp_3_tag(s2_io_metaReadResp_3_tag),
    .io_metaReadResp_3_valid(s2_io_metaReadResp_3_valid),
    .io_metaReadResp_3_dirty(s2_io_metaReadResp_3_dirty),
    .io_dataReadResp_0_data(s2_io_dataReadResp_0_data),
    .io_dataReadResp_1_data(s2_io_dataReadResp_1_data),
    .io_dataReadResp_2_data(s2_io_dataReadResp_2_data),
    .io_dataReadResp_3_data(s2_io_dataReadResp_3_data),
    .io_metaWriteBus_req_valid(s2_io_metaWriteBus_req_valid),
    .io_metaWriteBus_req_bits_setIdx(s2_io_metaWriteBus_req_bits_setIdx),
    .io_metaWriteBus_req_bits_data_tag(s2_io_metaWriteBus_req_bits_data_tag),
    .io_metaWriteBus_req_bits_data_dirty(s2_io_metaWriteBus_req_bits_data_dirty),
    .io_metaWriteBus_req_bits_waymask(s2_io_metaWriteBus_req_bits_waymask),
    .io_dataWriteBus_req_valid(s2_io_dataWriteBus_req_valid),
    .io_dataWriteBus_req_bits_setIdx(s2_io_dataWriteBus_req_bits_setIdx),
    .io_dataWriteBus_req_bits_data_data(s2_io_dataWriteBus_req_bits_data_data),
    .io_dataWriteBus_req_bits_waymask(s2_io_dataWriteBus_req_bits_waymask),
    .DISPLAY_ENABLE(s2_DISPLAY_ENABLE)
  );
  CacheStage3 s3 ( // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
    .clock(s3_clock),
    .reset(s3_reset),
    .io_in_ready(s3_io_in_ready),
    .io_in_valid(s3_io_in_valid),
    .io_in_bits_req_addr(s3_io_in_bits_req_addr),
    .io_in_bits_req_size(s3_io_in_bits_req_size),
    .io_in_bits_req_cmd(s3_io_in_bits_req_cmd),
    .io_in_bits_req_wmask(s3_io_in_bits_req_wmask),
    .io_in_bits_req_wdata(s3_io_in_bits_req_wdata),
    .io_in_bits_req_user(s3_io_in_bits_req_user),
    .io_in_bits_metas_0_tag(s3_io_in_bits_metas_0_tag),
    .io_in_bits_metas_0_valid(s3_io_in_bits_metas_0_valid),
    .io_in_bits_metas_0_dirty(s3_io_in_bits_metas_0_dirty),
    .io_in_bits_metas_1_tag(s3_io_in_bits_metas_1_tag),
    .io_in_bits_metas_1_valid(s3_io_in_bits_metas_1_valid),
    .io_in_bits_metas_1_dirty(s3_io_in_bits_metas_1_dirty),
    .io_in_bits_metas_2_tag(s3_io_in_bits_metas_2_tag),
    .io_in_bits_metas_2_valid(s3_io_in_bits_metas_2_valid),
    .io_in_bits_metas_2_dirty(s3_io_in_bits_metas_2_dirty),
    .io_in_bits_metas_3_tag(s3_io_in_bits_metas_3_tag),
    .io_in_bits_metas_3_valid(s3_io_in_bits_metas_3_valid),
    .io_in_bits_metas_3_dirty(s3_io_in_bits_metas_3_dirty),
    .io_in_bits_datas_0_data(s3_io_in_bits_datas_0_data),
    .io_in_bits_datas_1_data(s3_io_in_bits_datas_1_data),
    .io_in_bits_datas_2_data(s3_io_in_bits_datas_2_data),
    .io_in_bits_datas_3_data(s3_io_in_bits_datas_3_data),
    .io_in_bits_hit(s3_io_in_bits_hit),
    .io_in_bits_waymask(s3_io_in_bits_waymask),
    .io_in_bits_mmio(s3_io_in_bits_mmio),
    .io_in_bits_isForwardData(s3_io_in_bits_isForwardData),
    .io_in_bits_forwardData_data_data(s3_io_in_bits_forwardData_data_data),
    .io_in_bits_forwardData_waymask(s3_io_in_bits_forwardData_waymask),
    .io_out_ready(s3_io_out_ready),
    .io_out_valid(s3_io_out_valid),
    .io_out_bits_cmd(s3_io_out_bits_cmd),
    .io_out_bits_rdata(s3_io_out_bits_rdata),
    .io_out_bits_user(s3_io_out_bits_user),
    .io_isFinish(s3_io_isFinish),
    .io_flush(s3_io_flush),
    .io_dataReadBus_req_ready(s3_io_dataReadBus_req_ready),
    .io_dataReadBus_req_valid(s3_io_dataReadBus_req_valid),
    .io_dataReadBus_req_bits_setIdx(s3_io_dataReadBus_req_bits_setIdx),
    .io_dataReadBus_resp_data_0_data(s3_io_dataReadBus_resp_data_0_data),
    .io_dataReadBus_resp_data_1_data(s3_io_dataReadBus_resp_data_1_data),
    .io_dataReadBus_resp_data_2_data(s3_io_dataReadBus_resp_data_2_data),
    .io_dataReadBus_resp_data_3_data(s3_io_dataReadBus_resp_data_3_data),
    .io_dataWriteBus_req_valid(s3_io_dataWriteBus_req_valid),
    .io_dataWriteBus_req_bits_setIdx(s3_io_dataWriteBus_req_bits_setIdx),
    .io_dataWriteBus_req_bits_data_data(s3_io_dataWriteBus_req_bits_data_data),
    .io_dataWriteBus_req_bits_waymask(s3_io_dataWriteBus_req_bits_waymask),
    .io_metaWriteBus_req_valid(s3_io_metaWriteBus_req_valid),
    .io_metaWriteBus_req_bits_setIdx(s3_io_metaWriteBus_req_bits_setIdx),
    .io_metaWriteBus_req_bits_data_tag(s3_io_metaWriteBus_req_bits_data_tag),
    .io_metaWriteBus_req_bits_data_valid(s3_io_metaWriteBus_req_bits_data_valid),
    .io_metaWriteBus_req_bits_data_dirty(s3_io_metaWriteBus_req_bits_data_dirty),
    .io_metaWriteBus_req_bits_waymask(s3_io_metaWriteBus_req_bits_waymask),
    .io_mem_req_ready(s3_io_mem_req_ready),
    .io_mem_req_valid(s3_io_mem_req_valid),
    .io_mem_req_bits_addr(s3_io_mem_req_bits_addr),
    .io_mem_req_bits_size(s3_io_mem_req_bits_size),
    .io_mem_req_bits_cmd(s3_io_mem_req_bits_cmd),
    .io_mem_req_bits_wmask(s3_io_mem_req_bits_wmask),
    .io_mem_req_bits_wdata(s3_io_mem_req_bits_wdata),
    .io_mem_resp_ready(s3_io_mem_resp_ready),
    .io_mem_resp_valid(s3_io_mem_resp_valid),
    .io_mem_resp_bits_cmd(s3_io_mem_resp_bits_cmd),
    .io_mem_resp_bits_rdata(s3_io_mem_resp_bits_rdata),
    .io_mmio_req_ready(s3_io_mmio_req_ready),
    .io_mmio_req_valid(s3_io_mmio_req_valid),
    .io_mmio_req_bits_addr(s3_io_mmio_req_bits_addr),
    .io_mmio_resp_ready(s3_io_mmio_resp_ready),
    .io_mmio_resp_valid(s3_io_mmio_resp_valid),
    .io_mmio_resp_bits_rdata(s3_io_mmio_resp_bits_rdata),
    .io_cohResp_valid(s3_io_cohResp_valid),
    .DISPLAY_ENABLE(s3_DISPLAY_ENABLE)
  );
  SRAMTemplateWithArbiter metaArray ( // @[src/main/scala/nutcore/mem/Cache.scala 483:25]
    .clock(metaArray_clock),
    .reset(metaArray_reset),
    .io_r_0_req_ready(metaArray_io_r_0_req_ready),
    .io_r_0_req_valid(metaArray_io_r_0_req_valid),
    .io_r_0_req_bits_setIdx(metaArray_io_r_0_req_bits_setIdx),
    .io_r_0_resp_data_0_tag(metaArray_io_r_0_resp_data_0_tag),
    .io_r_0_resp_data_0_valid(metaArray_io_r_0_resp_data_0_valid),
    .io_r_0_resp_data_0_dirty(metaArray_io_r_0_resp_data_0_dirty),
    .io_r_0_resp_data_1_tag(metaArray_io_r_0_resp_data_1_tag),
    .io_r_0_resp_data_1_valid(metaArray_io_r_0_resp_data_1_valid),
    .io_r_0_resp_data_1_dirty(metaArray_io_r_0_resp_data_1_dirty),
    .io_r_0_resp_data_2_tag(metaArray_io_r_0_resp_data_2_tag),
    .io_r_0_resp_data_2_valid(metaArray_io_r_0_resp_data_2_valid),
    .io_r_0_resp_data_2_dirty(metaArray_io_r_0_resp_data_2_dirty),
    .io_r_0_resp_data_3_tag(metaArray_io_r_0_resp_data_3_tag),
    .io_r_0_resp_data_3_valid(metaArray_io_r_0_resp_data_3_valid),
    .io_r_0_resp_data_3_dirty(metaArray_io_r_0_resp_data_3_dirty),
    .io_w_req_valid(metaArray_io_w_req_valid),
    .io_w_req_bits_setIdx(metaArray_io_w_req_bits_setIdx),
    .io_w_req_bits_data_tag(metaArray_io_w_req_bits_data_tag),
    .io_w_req_bits_data_dirty(metaArray_io_w_req_bits_data_dirty),
    .io_w_req_bits_waymask(metaArray_io_w_req_bits_waymask)
  );
  SRAMTemplateWithArbiter_1 dataArray ( // @[src/main/scala/nutcore/mem/Cache.scala 484:25]
    .clock(dataArray_clock),
    .reset(dataArray_reset),
    .io_r_0_req_ready(dataArray_io_r_0_req_ready),
    .io_r_0_req_valid(dataArray_io_r_0_req_valid),
    .io_r_0_req_bits_setIdx(dataArray_io_r_0_req_bits_setIdx),
    .io_r_0_resp_data_0_data(dataArray_io_r_0_resp_data_0_data),
    .io_r_0_resp_data_1_data(dataArray_io_r_0_resp_data_1_data),
    .io_r_0_resp_data_2_data(dataArray_io_r_0_resp_data_2_data),
    .io_r_0_resp_data_3_data(dataArray_io_r_0_resp_data_3_data),
    .io_r_1_req_ready(dataArray_io_r_1_req_ready),
    .io_r_1_req_valid(dataArray_io_r_1_req_valid),
    .io_r_1_req_bits_setIdx(dataArray_io_r_1_req_bits_setIdx),
    .io_r_1_resp_data_0_data(dataArray_io_r_1_resp_data_0_data),
    .io_r_1_resp_data_1_data(dataArray_io_r_1_resp_data_1_data),
    .io_r_1_resp_data_2_data(dataArray_io_r_1_resp_data_2_data),
    .io_r_1_resp_data_3_data(dataArray_io_r_1_resp_data_3_data),
    .io_w_req_valid(dataArray_io_w_req_valid),
    .io_w_req_bits_setIdx(dataArray_io_w_req_bits_setIdx),
    .io_w_req_bits_data_data(dataArray_io_w_req_bits_data_data),
    .io_w_req_bits_waymask(dataArray_io_w_req_bits_waymask)
  );
  Arbiter_4 arb ( // @[src/main/scala/nutcore/mem/Cache.scala 493:19]
    .io_in_0_ready(arb_io_in_0_ready),
    .io_in_0_valid(arb_io_in_0_valid),
    .io_in_0_bits_addr(arb_io_in_0_bits_addr),
    .io_in_0_bits_user(arb_io_in_0_bits_user),
    .io_out_ready(arb_io_out_ready),
    .io_out_valid(arb_io_out_valid),
    .io_out_bits_addr(arb_io_out_bits_addr),
    .io_out_bits_user(arb_io_out_bits_user)
  );
  assign io_in_req_ready = arb_io_in_0_ready; // @[src/main/scala/nutcore/mem/Cache.scala 494:28]
  assign io_in_resp_valid = s3_io_out_valid; // @[src/main/scala/nutcore/mem/Cache.scala 510:98]
  assign io_in_resp_bits_rdata = s3_io_out_bits_rdata; // @[src/main/scala/nutcore/mem/Cache.scala 504:14]
  assign io_in_resp_bits_user = s3_io_out_bits_user; // @[src/main/scala/nutcore/mem/Cache.scala 504:14]
  assign io_out_mem_req_valid = s3_io_mem_req_valid; // @[src/main/scala/nutcore/mem/Cache.scala 506:14]
  assign io_out_mem_req_bits_addr = s3_io_mem_req_bits_addr; // @[src/main/scala/nutcore/mem/Cache.scala 506:14]
  assign io_out_mem_req_bits_cmd = s3_io_mem_req_bits_cmd; // @[src/main/scala/nutcore/mem/Cache.scala 506:14]
  assign io_out_mem_req_bits_wdata = s3_io_mem_req_bits_wdata; // @[src/main/scala/nutcore/mem/Cache.scala 506:14]
  assign io_mmio_req_valid = s3_io_mmio_req_valid; // @[src/main/scala/nutcore/mem/Cache.scala 507:11]
  assign io_mmio_req_bits_addr = s3_io_mmio_req_bits_addr; // @[src/main/scala/nutcore/mem/Cache.scala 507:11]
  assign io_empty = ~s2_io_in_valid & ~s3_io_in_valid; // @[src/main/scala/nutcore/mem/Cache.scala 508:31]
  assign s1_clock = clock;
  assign s1_reset = reset;
  assign s1_io_in_valid = arb_io_out_valid; // @[src/main/scala/nutcore/mem/Cache.scala 496:12]
  assign s1_io_in_bits_addr = arb_io_out_bits_addr; // @[src/main/scala/nutcore/mem/Cache.scala 496:12]
  assign s1_io_in_bits_size = 3'h3; // @[src/main/scala/nutcore/mem/Cache.scala 496:12]
  assign s1_io_in_bits_cmd = 4'h0; // @[src/main/scala/nutcore/mem/Cache.scala 496:12]
  assign s1_io_in_bits_wmask = 8'h0; // @[src/main/scala/nutcore/mem/Cache.scala 496:12]
  assign s1_io_in_bits_wdata = 64'h0; // @[src/main/scala/nutcore/mem/Cache.scala 496:12]
  assign s1_io_in_bits_user = arb_io_out_bits_user; // @[src/main/scala/nutcore/mem/Cache.scala 496:12]
  assign s1_io_out_ready = s2_io_in_ready; // @[src/main/scala/utils/Pipeline.scala 29:16]
  assign s1_io_metaReadBus_req_ready = metaArray_io_r_0_req_ready; // @[src/main/scala/nutcore/mem/Cache.scala 528:21]
  assign s1_io_metaReadBus_resp_data_0_tag = metaArray_io_r_0_resp_data_0_tag; // @[src/main/scala/nutcore/mem/Cache.scala 528:21]
  assign s1_io_metaReadBus_resp_data_0_valid = metaArray_io_r_0_resp_data_0_valid; // @[src/main/scala/nutcore/mem/Cache.scala 528:21]
  assign s1_io_metaReadBus_resp_data_0_dirty = metaArray_io_r_0_resp_data_0_dirty; // @[src/main/scala/nutcore/mem/Cache.scala 528:21]
  assign s1_io_metaReadBus_resp_data_1_tag = metaArray_io_r_0_resp_data_1_tag; // @[src/main/scala/nutcore/mem/Cache.scala 528:21]
  assign s1_io_metaReadBus_resp_data_1_valid = metaArray_io_r_0_resp_data_1_valid; // @[src/main/scala/nutcore/mem/Cache.scala 528:21]
  assign s1_io_metaReadBus_resp_data_1_dirty = metaArray_io_r_0_resp_data_1_dirty; // @[src/main/scala/nutcore/mem/Cache.scala 528:21]
  assign s1_io_metaReadBus_resp_data_2_tag = metaArray_io_r_0_resp_data_2_tag; // @[src/main/scala/nutcore/mem/Cache.scala 528:21]
  assign s1_io_metaReadBus_resp_data_2_valid = metaArray_io_r_0_resp_data_2_valid; // @[src/main/scala/nutcore/mem/Cache.scala 528:21]
  assign s1_io_metaReadBus_resp_data_2_dirty = metaArray_io_r_0_resp_data_2_dirty; // @[src/main/scala/nutcore/mem/Cache.scala 528:21]
  assign s1_io_metaReadBus_resp_data_3_tag = metaArray_io_r_0_resp_data_3_tag; // @[src/main/scala/nutcore/mem/Cache.scala 528:21]
  assign s1_io_metaReadBus_resp_data_3_valid = metaArray_io_r_0_resp_data_3_valid; // @[src/main/scala/nutcore/mem/Cache.scala 528:21]
  assign s1_io_metaReadBus_resp_data_3_dirty = metaArray_io_r_0_resp_data_3_dirty; // @[src/main/scala/nutcore/mem/Cache.scala 528:21]
  assign s1_io_dataReadBus_req_ready = dataArray_io_r_0_req_ready; // @[src/main/scala/nutcore/mem/Cache.scala 529:21]
  assign s1_io_dataReadBus_resp_data_0_data = dataArray_io_r_0_resp_data_0_data; // @[src/main/scala/nutcore/mem/Cache.scala 529:21]
  assign s1_io_dataReadBus_resp_data_1_data = dataArray_io_r_0_resp_data_1_data; // @[src/main/scala/nutcore/mem/Cache.scala 529:21]
  assign s1_io_dataReadBus_resp_data_2_data = dataArray_io_r_0_resp_data_2_data; // @[src/main/scala/nutcore/mem/Cache.scala 529:21]
  assign s1_io_dataReadBus_resp_data_3_data = dataArray_io_r_0_resp_data_3_data; // @[src/main/scala/nutcore/mem/Cache.scala 529:21]
  assign s1_DISPLAY_ENABLE = DISPLAY_ENABLE;
  assign s2_clock = clock;
  assign s2_reset = reset;
  assign s2_io_in_valid = valid; // @[src/main/scala/utils/Pipeline.scala 31:17]
  assign s2_io_in_bits_req_addr = s2_io_in_bits_r_req_addr; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign s2_io_in_bits_req_size = 3'h3; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign s2_io_in_bits_req_cmd = 4'h0; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign s2_io_in_bits_req_wmask = 8'h0; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign s2_io_in_bits_req_wdata = 64'h0; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign s2_io_in_bits_req_user = s2_io_in_bits_r_req_user; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign s2_io_out_ready = s3_io_in_ready; // @[src/main/scala/utils/Pipeline.scala 29:16]
  assign s2_io_metaReadResp_0_tag = s1_io_metaReadBus_resp_data_0_tag; // @[src/main/scala/nutcore/mem/Cache.scala 535:22]
  assign s2_io_metaReadResp_0_valid = s1_io_metaReadBus_resp_data_0_valid; // @[src/main/scala/nutcore/mem/Cache.scala 535:22]
  assign s2_io_metaReadResp_0_dirty = s1_io_metaReadBus_resp_data_0_dirty; // @[src/main/scala/nutcore/mem/Cache.scala 535:22]
  assign s2_io_metaReadResp_1_tag = s1_io_metaReadBus_resp_data_1_tag; // @[src/main/scala/nutcore/mem/Cache.scala 535:22]
  assign s2_io_metaReadResp_1_valid = s1_io_metaReadBus_resp_data_1_valid; // @[src/main/scala/nutcore/mem/Cache.scala 535:22]
  assign s2_io_metaReadResp_1_dirty = s1_io_metaReadBus_resp_data_1_dirty; // @[src/main/scala/nutcore/mem/Cache.scala 535:22]
  assign s2_io_metaReadResp_2_tag = s1_io_metaReadBus_resp_data_2_tag; // @[src/main/scala/nutcore/mem/Cache.scala 535:22]
  assign s2_io_metaReadResp_2_valid = s1_io_metaReadBus_resp_data_2_valid; // @[src/main/scala/nutcore/mem/Cache.scala 535:22]
  assign s2_io_metaReadResp_2_dirty = s1_io_metaReadBus_resp_data_2_dirty; // @[src/main/scala/nutcore/mem/Cache.scala 535:22]
  assign s2_io_metaReadResp_3_tag = s1_io_metaReadBus_resp_data_3_tag; // @[src/main/scala/nutcore/mem/Cache.scala 535:22]
  assign s2_io_metaReadResp_3_valid = s1_io_metaReadBus_resp_data_3_valid; // @[src/main/scala/nutcore/mem/Cache.scala 535:22]
  assign s2_io_metaReadResp_3_dirty = s1_io_metaReadBus_resp_data_3_dirty; // @[src/main/scala/nutcore/mem/Cache.scala 535:22]
  assign s2_io_dataReadResp_0_data = s1_io_dataReadBus_resp_data_0_data; // @[src/main/scala/nutcore/mem/Cache.scala 536:22]
  assign s2_io_dataReadResp_1_data = s1_io_dataReadBus_resp_data_1_data; // @[src/main/scala/nutcore/mem/Cache.scala 536:22]
  assign s2_io_dataReadResp_2_data = s1_io_dataReadBus_resp_data_2_data; // @[src/main/scala/nutcore/mem/Cache.scala 536:22]
  assign s2_io_dataReadResp_3_data = s1_io_dataReadBus_resp_data_3_data; // @[src/main/scala/nutcore/mem/Cache.scala 536:22]
  assign s2_io_metaWriteBus_req_valid = s3_io_metaWriteBus_req_valid; // @[src/main/scala/nutcore/mem/Cache.scala 538:22]
  assign s2_io_metaWriteBus_req_bits_setIdx = s3_io_metaWriteBus_req_bits_setIdx; // @[src/main/scala/nutcore/mem/Cache.scala 538:22]
  assign s2_io_metaWriteBus_req_bits_data_tag = s3_io_metaWriteBus_req_bits_data_tag; // @[src/main/scala/nutcore/mem/Cache.scala 538:22]
  assign s2_io_metaWriteBus_req_bits_data_dirty = s3_io_metaWriteBus_req_bits_data_dirty; // @[src/main/scala/nutcore/mem/Cache.scala 538:22]
  assign s2_io_metaWriteBus_req_bits_waymask = s3_io_metaWriteBus_req_bits_waymask; // @[src/main/scala/nutcore/mem/Cache.scala 538:22]
  assign s2_io_dataWriteBus_req_valid = s3_io_dataWriteBus_req_valid; // @[src/main/scala/nutcore/mem/Cache.scala 537:22]
  assign s2_io_dataWriteBus_req_bits_setIdx = s3_io_dataWriteBus_req_bits_setIdx; // @[src/main/scala/nutcore/mem/Cache.scala 537:22]
  assign s2_io_dataWriteBus_req_bits_data_data = s3_io_dataWriteBus_req_bits_data_data; // @[src/main/scala/nutcore/mem/Cache.scala 537:22]
  assign s2_io_dataWriteBus_req_bits_waymask = s3_io_dataWriteBus_req_bits_waymask; // @[src/main/scala/nutcore/mem/Cache.scala 537:22]
  assign s2_DISPLAY_ENABLE = DISPLAY_ENABLE;
  assign s3_clock = clock;
  assign s3_reset = reset;
  assign s3_io_in_valid = valid_1; // @[src/main/scala/utils/Pipeline.scala 31:17]
  assign s3_io_in_bits_req_addr = s3_io_in_bits_r_req_addr; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign s3_io_in_bits_req_size = 3'h3; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign s3_io_in_bits_req_cmd = 4'h0; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign s3_io_in_bits_req_wmask = 8'h0; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign s3_io_in_bits_req_wdata = 64'h0; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign s3_io_in_bits_req_user = s3_io_in_bits_r_req_user; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign s3_io_in_bits_metas_0_tag = s3_io_in_bits_r_metas_0_tag; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign s3_io_in_bits_metas_0_valid = s3_io_in_bits_r_metas_0_valid; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign s3_io_in_bits_metas_0_dirty = s3_io_in_bits_r_metas_0_dirty; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign s3_io_in_bits_metas_1_tag = s3_io_in_bits_r_metas_1_tag; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign s3_io_in_bits_metas_1_valid = s3_io_in_bits_r_metas_1_valid; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign s3_io_in_bits_metas_1_dirty = s3_io_in_bits_r_metas_1_dirty; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign s3_io_in_bits_metas_2_tag = s3_io_in_bits_r_metas_2_tag; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign s3_io_in_bits_metas_2_valid = s3_io_in_bits_r_metas_2_valid; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign s3_io_in_bits_metas_2_dirty = s3_io_in_bits_r_metas_2_dirty; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign s3_io_in_bits_metas_3_tag = s3_io_in_bits_r_metas_3_tag; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign s3_io_in_bits_metas_3_valid = s3_io_in_bits_r_metas_3_valid; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign s3_io_in_bits_metas_3_dirty = s3_io_in_bits_r_metas_3_dirty; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign s3_io_in_bits_datas_0_data = s3_io_in_bits_r_datas_0_data; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign s3_io_in_bits_datas_1_data = s3_io_in_bits_r_datas_1_data; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign s3_io_in_bits_datas_2_data = s3_io_in_bits_r_datas_2_data; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign s3_io_in_bits_datas_3_data = s3_io_in_bits_r_datas_3_data; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign s3_io_in_bits_hit = s3_io_in_bits_r_hit; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign s3_io_in_bits_waymask = s3_io_in_bits_r_waymask; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign s3_io_in_bits_mmio = s3_io_in_bits_r_mmio; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign s3_io_in_bits_isForwardData = s3_io_in_bits_r_isForwardData; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign s3_io_in_bits_forwardData_data_data = s3_io_in_bits_r_forwardData_data_data; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign s3_io_in_bits_forwardData_waymask = s3_io_in_bits_r_forwardData_waymask; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign s3_io_out_ready = io_in_resp_ready; // @[src/main/scala/nutcore/mem/Cache.scala 504:14]
  assign s3_io_flush = io_flush[1]; // @[src/main/scala/nutcore/mem/Cache.scala 505:26]
  assign s3_io_dataReadBus_req_ready = dataArray_io_r_1_req_ready; // @[src/main/scala/nutcore/mem/Cache.scala 530:21]
  assign s3_io_dataReadBus_resp_data_0_data = dataArray_io_r_1_resp_data_0_data; // @[src/main/scala/nutcore/mem/Cache.scala 530:21]
  assign s3_io_dataReadBus_resp_data_1_data = dataArray_io_r_1_resp_data_1_data; // @[src/main/scala/nutcore/mem/Cache.scala 530:21]
  assign s3_io_dataReadBus_resp_data_2_data = dataArray_io_r_1_resp_data_2_data; // @[src/main/scala/nutcore/mem/Cache.scala 530:21]
  assign s3_io_dataReadBus_resp_data_3_data = dataArray_io_r_1_resp_data_3_data; // @[src/main/scala/nutcore/mem/Cache.scala 530:21]
  assign s3_io_mem_req_ready = io_out_mem_req_ready; // @[src/main/scala/nutcore/mem/Cache.scala 506:14]
  assign s3_io_mem_resp_valid = io_out_mem_resp_valid; // @[src/main/scala/nutcore/mem/Cache.scala 506:14]
  assign s3_io_mem_resp_bits_cmd = io_out_mem_resp_bits_cmd; // @[src/main/scala/nutcore/mem/Cache.scala 506:14]
  assign s3_io_mem_resp_bits_rdata = io_out_mem_resp_bits_rdata; // @[src/main/scala/nutcore/mem/Cache.scala 506:14]
  assign s3_io_mmio_req_ready = io_mmio_req_ready; // @[src/main/scala/nutcore/mem/Cache.scala 507:11]
  assign s3_io_mmio_resp_valid = io_mmio_resp_valid; // @[src/main/scala/nutcore/mem/Cache.scala 507:11]
  assign s3_io_mmio_resp_bits_rdata = io_mmio_resp_bits_rdata; // @[src/main/scala/nutcore/mem/Cache.scala 507:11]
  assign s3_DISPLAY_ENABLE = DISPLAY_ENABLE;
  assign metaArray_clock = clock;
  assign metaArray_reset = reset | MOUFlushICache; // @[src/main/scala/nutcore/mem/Cache.scala 490:37]
  assign metaArray_io_r_0_req_valid = s1_io_metaReadBus_req_valid; // @[src/main/scala/nutcore/mem/Cache.scala 528:21]
  assign metaArray_io_r_0_req_bits_setIdx = s1_io_metaReadBus_req_bits_setIdx; // @[src/main/scala/nutcore/mem/Cache.scala 528:21]
  assign metaArray_io_w_req_valid = s3_io_metaWriteBus_req_valid; // @[src/main/scala/nutcore/mem/Cache.scala 532:18]
  assign metaArray_io_w_req_bits_setIdx = s3_io_metaWriteBus_req_bits_setIdx; // @[src/main/scala/nutcore/mem/Cache.scala 532:18]
  assign metaArray_io_w_req_bits_data_tag = s3_io_metaWriteBus_req_bits_data_tag; // @[src/main/scala/nutcore/mem/Cache.scala 532:18]
  assign metaArray_io_w_req_bits_data_dirty = s3_io_metaWriteBus_req_bits_data_dirty; // @[src/main/scala/nutcore/mem/Cache.scala 532:18]
  assign metaArray_io_w_req_bits_waymask = s3_io_metaWriteBus_req_bits_waymask; // @[src/main/scala/nutcore/mem/Cache.scala 532:18]
  assign dataArray_clock = clock;
  assign dataArray_reset = reset;
  assign dataArray_io_r_0_req_valid = s1_io_dataReadBus_req_valid; // @[src/main/scala/nutcore/mem/Cache.scala 529:21]
  assign dataArray_io_r_0_req_bits_setIdx = s1_io_dataReadBus_req_bits_setIdx; // @[src/main/scala/nutcore/mem/Cache.scala 529:21]
  assign dataArray_io_r_1_req_valid = s3_io_dataReadBus_req_valid; // @[src/main/scala/nutcore/mem/Cache.scala 530:21]
  assign dataArray_io_r_1_req_bits_setIdx = s3_io_dataReadBus_req_bits_setIdx; // @[src/main/scala/nutcore/mem/Cache.scala 530:21]
  assign dataArray_io_w_req_valid = s3_io_dataWriteBus_req_valid; // @[src/main/scala/nutcore/mem/Cache.scala 533:18]
  assign dataArray_io_w_req_bits_setIdx = s3_io_dataWriteBus_req_bits_setIdx; // @[src/main/scala/nutcore/mem/Cache.scala 533:18]
  assign dataArray_io_w_req_bits_data_data = s3_io_dataWriteBus_req_bits_data_data; // @[src/main/scala/nutcore/mem/Cache.scala 533:18]
  assign dataArray_io_w_req_bits_waymask = s3_io_dataWriteBus_req_bits_waymask; // @[src/main/scala/nutcore/mem/Cache.scala 533:18]
  assign arb_io_in_0_valid = io_in_req_valid; // @[src/main/scala/nutcore/mem/Cache.scala 494:28]
  assign arb_io_in_0_bits_addr = io_in_req_bits_addr; // @[src/main/scala/nutcore/mem/Cache.scala 494:28]
  assign arb_io_in_0_bits_user = io_in_req_bits_user; // @[src/main/scala/nutcore/mem/Cache.scala 494:28]
  assign arb_io_out_ready = s1_io_in_ready; // @[src/main/scala/nutcore/mem/Cache.scala 496:12]
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/utils/Pipeline.scala 24:24]
      valid <= 1'h0; // @[src/main/scala/utils/Pipeline.scala 24:24]
    end else if (io_flush[0]) begin // @[src/main/scala/utils/Pipeline.scala 27:20]
      valid <= 1'h0; // @[src/main/scala/utils/Pipeline.scala 27:28]
    end else begin
      valid <= _GEN_1;
    end
    if (_T_2) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      s2_io_in_bits_r_req_addr <= s1_io_out_bits_req_addr; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_2) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      s2_io_in_bits_r_req_user <= s1_io_out_bits_req_user; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (reset) begin // @[src/main/scala/utils/Pipeline.scala 24:24]
      valid_1 <= 1'h0; // @[src/main/scala/utils/Pipeline.scala 24:24]
    end else if (io_flush[1]) begin // @[src/main/scala/utils/Pipeline.scala 27:20]
      valid_1 <= 1'h0; // @[src/main/scala/utils/Pipeline.scala 27:28]
    end else begin
      valid_1 <= _GEN_10;
    end
    if (_T_4) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      s3_io_in_bits_r_req_addr <= s2_io_out_bits_req_addr; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_4) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      s3_io_in_bits_r_req_user <= s2_io_out_bits_req_user; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_4) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      s3_io_in_bits_r_metas_0_tag <= s2_io_out_bits_metas_0_tag; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_4) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      s3_io_in_bits_r_metas_0_valid <= s2_io_out_bits_metas_0_valid; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_4) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      s3_io_in_bits_r_metas_0_dirty <= s2_io_out_bits_metas_0_dirty; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_4) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      s3_io_in_bits_r_metas_1_tag <= s2_io_out_bits_metas_1_tag; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_4) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      s3_io_in_bits_r_metas_1_valid <= s2_io_out_bits_metas_1_valid; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_4) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      s3_io_in_bits_r_metas_1_dirty <= s2_io_out_bits_metas_1_dirty; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_4) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      s3_io_in_bits_r_metas_2_tag <= s2_io_out_bits_metas_2_tag; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_4) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      s3_io_in_bits_r_metas_2_valid <= s2_io_out_bits_metas_2_valid; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_4) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      s3_io_in_bits_r_metas_2_dirty <= s2_io_out_bits_metas_2_dirty; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_4) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      s3_io_in_bits_r_metas_3_tag <= s2_io_out_bits_metas_3_tag; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_4) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      s3_io_in_bits_r_metas_3_valid <= s2_io_out_bits_metas_3_valid; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_4) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      s3_io_in_bits_r_metas_3_dirty <= s2_io_out_bits_metas_3_dirty; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_4) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      s3_io_in_bits_r_datas_0_data <= s2_io_out_bits_datas_0_data; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_4) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      s3_io_in_bits_r_datas_1_data <= s2_io_out_bits_datas_1_data; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_4) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      s3_io_in_bits_r_datas_2_data <= s2_io_out_bits_datas_2_data; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_4) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      s3_io_in_bits_r_datas_3_data <= s2_io_out_bits_datas_3_data; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_4) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      s3_io_in_bits_r_hit <= s2_io_out_bits_hit; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_4) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      s3_io_in_bits_r_waymask <= s2_io_out_bits_waymask; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_4) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      s3_io_in_bits_r_mmio <= s2_io_out_bits_mmio; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_4) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      s3_io_in_bits_r_isForwardData <= s2_io_out_bits_isForwardData; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_4) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      s3_io_in_bits_r_forwardData_data_data <= s2_io_out_bits_forwardData_data_data; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_4) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      s3_io_in_bits_r_forwardData_waymask <= s2_io_out_bits_forwardData_waymask; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (reset) begin // @[src/main/scala/utils/GTimer.scala 24:20]
      c <= 64'h0; // @[src/main/scala/utils/GTimer.scala 24:20]
    end else begin
      c <= _c_T_1; // @[src/main/scala/utils/GTimer.scala 25:7]
    end
    if (reset) begin // @[src/main/scala/utils/GTimer.scala 24:20]
      c_1 <= 64'h0; // @[src/main/scala/utils/GTimer.scala 24:20]
    end else begin
      c_1 <= _c_T_3; // @[src/main/scala/utils/GTimer.scala 25:7]
    end
    if (reset) begin // @[src/main/scala/utils/GTimer.scala 24:20]
      c_2 <= 64'h0; // @[src/main/scala/utils/GTimer.scala 24:20]
    end else begin
      c_2 <= _c_T_5; // @[src/main/scala/utils/GTimer.scala 25:7]
    end
    if (reset) begin // @[src/main/scala/utils/GTimer.scala 24:20]
      c_3 <= 64'h0; // @[src/main/scala/utils/GTimer.scala 24:20]
    end else begin
      c_3 <= _c_T_7; // @[src/main/scala/utils/GTimer.scala 25:7]
    end
    if (reset) begin // @[src/main/scala/utils/GTimer.scala 24:20]
      c_4 <= 64'h0; // @[src/main/scala/utils/GTimer.scala 24:20]
    end else begin
      c_4 <= _c_T_9; // @[src/main/scala/utils/GTimer.scala 25:7]
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & ~reset) begin
          $fwrite(32'h80000002,"[%d] Cache: ",c); // @[src/main/scala/utils/Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_7) begin
          $fwrite(32'h80000002,"InReq(%d, %d) InResp(%d, %d) \n",io_in_req_valid,io_in_req_ready,io_in_resp_valid,
            io_in_resp_ready); // @[src/main/scala/utils/Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & ~reset) begin
          $fwrite(32'h80000002,"[%d] Cache: ",c_1); // @[src/main/scala/utils/Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_7) begin
          $fwrite(32'h80000002,"{IN s1:(%d,%d), s2:(%d,%d), s3:(%d,%d)} {OUT s1:(%d,%d), s2:(%d,%d), s3:(%d,%d)}\n",
            s1_io_in_valid,s1_io_in_ready,s2_io_in_valid,s2_io_in_ready,s3_io_in_valid,s3_io_in_ready,s1_io_out_valid,
            s1_io_out_ready,s2_io_out_valid,s2_io_out_ready,s3_io_out_valid,s3_io_out_ready); // @[src/main/scala/utils/Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (s1_io_in_valid & DISPLAY_ENABLE & ~reset) begin
          $fwrite(32'h80000002,"[%d] Cache: ",c_2); // @[src/main/scala/utils/Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_41 & _T_7) begin
          $fwrite(32'h80000002,"[icache.S1]: addr = 0x%x, cmd = %d, size = %d, wmask = 0x%x, wdata = 0x%x\n",
            s1_io_in_bits_addr,s1_io_in_bits_cmd,s1_io_in_bits_size,s1_io_in_bits_wmask,s1_io_in_bits_wdata); // @[src/main/scala/utils/Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (s2_io_in_valid & DISPLAY_ENABLE & ~reset) begin
          $fwrite(32'h80000002,"[%d] Cache: ",c_3); // @[src/main/scala/utils/Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_43 & _T_7) begin
          $fwrite(32'h80000002,"[icache.S2]: addr = 0x%x, cmd = %d, size = %d, wmask = 0x%x, wdata = 0x%x\n",
            s2_io_in_bits_req_addr,s2_io_in_bits_req_cmd,s2_io_in_bits_req_size,s2_io_in_bits_req_wmask,
            s2_io_in_bits_req_wdata); // @[src/main/scala/utils/Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (s3_io_in_valid & DISPLAY_ENABLE & ~reset) begin
          $fwrite(32'h80000002,"[%d] Cache: ",c_4); // @[src/main/scala/utils/Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_45 & _T_7) begin
          $fwrite(32'h80000002,"[icache.S3]: addr = 0x%x, cmd = %d, size = %d, wmask = 0x%x, wdata = 0x%x\n",
            s3_io_in_bits_req_addr,s3_io_in_bits_req_cmd,s3_io_in_bits_req_size,s3_io_in_bits_req_wmask,
            s3_io_in_bits_req_wdata); // @[src/main/scala/utils/Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  valid = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  s2_io_in_bits_r_req_addr = _RAND_1[31:0];
  _RAND_2 = {3{`RANDOM}};
  s2_io_in_bits_r_req_user = _RAND_2[86:0];
  _RAND_3 = {1{`RANDOM}};
  valid_1 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  s3_io_in_bits_r_req_addr = _RAND_4[31:0];
  _RAND_5 = {3{`RANDOM}};
  s3_io_in_bits_r_req_user = _RAND_5[86:0];
  _RAND_6 = {1{`RANDOM}};
  s3_io_in_bits_r_metas_0_tag = _RAND_6[18:0];
  _RAND_7 = {1{`RANDOM}};
  s3_io_in_bits_r_metas_0_valid = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  s3_io_in_bits_r_metas_0_dirty = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  s3_io_in_bits_r_metas_1_tag = _RAND_9[18:0];
  _RAND_10 = {1{`RANDOM}};
  s3_io_in_bits_r_metas_1_valid = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  s3_io_in_bits_r_metas_1_dirty = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  s3_io_in_bits_r_metas_2_tag = _RAND_12[18:0];
  _RAND_13 = {1{`RANDOM}};
  s3_io_in_bits_r_metas_2_valid = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  s3_io_in_bits_r_metas_2_dirty = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  s3_io_in_bits_r_metas_3_tag = _RAND_15[18:0];
  _RAND_16 = {1{`RANDOM}};
  s3_io_in_bits_r_metas_3_valid = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  s3_io_in_bits_r_metas_3_dirty = _RAND_17[0:0];
  _RAND_18 = {2{`RANDOM}};
  s3_io_in_bits_r_datas_0_data = _RAND_18[63:0];
  _RAND_19 = {2{`RANDOM}};
  s3_io_in_bits_r_datas_1_data = _RAND_19[63:0];
  _RAND_20 = {2{`RANDOM}};
  s3_io_in_bits_r_datas_2_data = _RAND_20[63:0];
  _RAND_21 = {2{`RANDOM}};
  s3_io_in_bits_r_datas_3_data = _RAND_21[63:0];
  _RAND_22 = {1{`RANDOM}};
  s3_io_in_bits_r_hit = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  s3_io_in_bits_r_waymask = _RAND_23[3:0];
  _RAND_24 = {1{`RANDOM}};
  s3_io_in_bits_r_mmio = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  s3_io_in_bits_r_isForwardData = _RAND_25[0:0];
  _RAND_26 = {2{`RANDOM}};
  s3_io_in_bits_r_forwardData_data_data = _RAND_26[63:0];
  _RAND_27 = {1{`RANDOM}};
  s3_io_in_bits_r_forwardData_waymask = _RAND_27[3:0];
  _RAND_28 = {2{`RANDOM}};
  c = _RAND_28[63:0];
  _RAND_29 = {2{`RANDOM}};
  c_1 = _RAND_29[63:0];
  _RAND_30 = {2{`RANDOM}};
  c_2 = _RAND_30[63:0];
  _RAND_31 = {2{`RANDOM}};
  c_3 = _RAND_31[63:0];
  _RAND_32 = {2{`RANDOM}};
  c_4 = _RAND_32[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module EmbeddedTLBExec_1(
  input          clock,
  input          reset,
  output         io_in_ready, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 178:14]
  input          io_in_valid, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 178:14]
  input  [38:0]  io_in_bits_addr, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 178:14]
  input  [2:0]   io_in_bits_size, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 178:14]
  input  [3:0]   io_in_bits_cmd, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 178:14]
  input  [7:0]   io_in_bits_wmask, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 178:14]
  input  [63:0]  io_in_bits_wdata, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 178:14]
  input          io_out_ready, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 178:14]
  output         io_out_valid, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 178:14]
  output [31:0]  io_out_bits_addr, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 178:14]
  output [2:0]   io_out_bits_size, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 178:14]
  output [3:0]   io_out_bits_cmd, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 178:14]
  output [7:0]   io_out_bits_wmask, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 178:14]
  output [63:0]  io_out_bits_wdata, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 178:14]
  input  [120:0] io_md_0, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 178:14]
  input  [120:0] io_md_1, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 178:14]
  input  [120:0] io_md_2, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 178:14]
  input  [120:0] io_md_3, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 178:14]
  output         io_mdWrite_wen, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 178:14]
  output [3:0]   io_mdWrite_windex, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 178:14]
  output [3:0]   io_mdWrite_waymask, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 178:14]
  output [120:0] io_mdWrite_wdata, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 178:14]
  input          io_mdReady, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 178:14]
  input          io_mem_req_ready, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 178:14]
  output         io_mem_req_valid, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 178:14]
  output [31:0]  io_mem_req_bits_addr, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 178:14]
  output [2:0]   io_mem_req_bits_size, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 178:14]
  output [3:0]   io_mem_req_bits_cmd, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 178:14]
  output [7:0]   io_mem_req_bits_wmask, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 178:14]
  output [63:0]  io_mem_req_bits_wdata, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 178:14]
  output         io_mem_resp_ready, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 178:14]
  input          io_mem_resp_valid, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 178:14]
  input  [3:0]   io_mem_resp_bits_cmd, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 178:14]
  input  [63:0]  io_mem_resp_bits_rdata, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 178:14]
  input  [63:0]  io_satp, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 178:14]
  input  [1:0]   io_pf_priviledgeMode, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 178:14]
  input          io_pf_status_sum, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 178:14]
  input          io_pf_status_mxr, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 178:14]
  output         io_pf_loadPF, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 178:14]
  output         io_pf_storePF, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 178:14]
  output [38:0]  io_pf_addr, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 178:14]
  output         io_ipf, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 178:14]
  output         io_isFinish, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 178:14]
  input          ISAMO,
  input          DISPLAY_ENABLE
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [63:0] _RAND_20;
  reg [63:0] _RAND_21;
  reg [63:0] _RAND_22;
  reg [63:0] _RAND_23;
  reg [63:0] _RAND_24;
  reg [63:0] _RAND_25;
  reg [63:0] _RAND_26;
  reg [63:0] _RAND_27;
`endif // RANDOMIZE_REG_INIT
  wire [8:0] vpn_vpn0 = io_in_bits_addr[20:12]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 198:54]
  wire [8:0] vpn_vpn1 = io_in_bits_addr[29:21]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 198:54]
  wire [8:0] vpn_vpn2 = io_in_bits_addr[38:30]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 198:54]
  wire [19:0] satp_ppn = io_satp[19:0]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 200:30]
  wire [15:0] satp_asid = io_satp[59:44]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 200:30]
  wire [17:0] hitVec_hi = {vpn_vpn2,vpn_vpn1}; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 209:201]
  wire [26:0] _hitVec_T_34 = {vpn_vpn2,vpn_vpn1,vpn_vpn0}; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 209:201]
  wire [26:0] _hitVec_T_35 = {9'h1ff,io_md_0[77:60]}; // @[src/main/scala/nutcore/mem/TLB.scala 131:9]
  wire [26:0] _hitVec_T_36 = _hitVec_T_35 & io_md_0[120:94]; // @[src/main/scala/nutcore/mem/TLB.scala 131:37]
  wire [26:0] _hitVec_T_38 = _hitVec_T_35 & _hitVec_T_34; // @[src/main/scala/nutcore/mem/TLB.scala 131:84]
  wire  _hitVec_T_39 = _hitVec_T_36 == _hitVec_T_38; // @[src/main/scala/nutcore/mem/TLB.scala 131:48]
  wire  _hitVec_T_40 = io_md_0[52] & io_md_0[93:78] == satp_asid & _hitVec_T_39; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 209:132]
  wire [26:0] _hitVec_T_76 = {9'h1ff,io_md_1[77:60]}; // @[src/main/scala/nutcore/mem/TLB.scala 131:9]
  wire [26:0] _hitVec_T_77 = _hitVec_T_76 & io_md_1[120:94]; // @[src/main/scala/nutcore/mem/TLB.scala 131:37]
  wire [26:0] _hitVec_T_79 = _hitVec_T_76 & _hitVec_T_34; // @[src/main/scala/nutcore/mem/TLB.scala 131:84]
  wire  _hitVec_T_80 = _hitVec_T_77 == _hitVec_T_79; // @[src/main/scala/nutcore/mem/TLB.scala 131:48]
  wire  _hitVec_T_81 = io_md_1[52] & io_md_1[93:78] == satp_asid & _hitVec_T_80; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 209:132]
  wire [26:0] _hitVec_T_117 = {9'h1ff,io_md_2[77:60]}; // @[src/main/scala/nutcore/mem/TLB.scala 131:9]
  wire [26:0] _hitVec_T_118 = _hitVec_T_117 & io_md_2[120:94]; // @[src/main/scala/nutcore/mem/TLB.scala 131:37]
  wire [26:0] _hitVec_T_120 = _hitVec_T_117 & _hitVec_T_34; // @[src/main/scala/nutcore/mem/TLB.scala 131:84]
  wire  _hitVec_T_121 = _hitVec_T_118 == _hitVec_T_120; // @[src/main/scala/nutcore/mem/TLB.scala 131:48]
  wire  _hitVec_T_122 = io_md_2[52] & io_md_2[93:78] == satp_asid & _hitVec_T_121; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 209:132]
  wire [26:0] _hitVec_T_158 = {9'h1ff,io_md_3[77:60]}; // @[src/main/scala/nutcore/mem/TLB.scala 131:9]
  wire [26:0] _hitVec_T_159 = _hitVec_T_158 & io_md_3[120:94]; // @[src/main/scala/nutcore/mem/TLB.scala 131:37]
  wire [26:0] _hitVec_T_161 = _hitVec_T_158 & _hitVec_T_34; // @[src/main/scala/nutcore/mem/TLB.scala 131:84]
  wire  _hitVec_T_162 = _hitVec_T_159 == _hitVec_T_161; // @[src/main/scala/nutcore/mem/TLB.scala 131:48]
  wire  _hitVec_T_163 = io_md_3[52] & io_md_3[93:78] == satp_asid & _hitVec_T_162; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 209:132]
  wire [3:0] hitVec = {_hitVec_T_163,_hitVec_T_122,_hitVec_T_81,_hitVec_T_40}; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 209:211]
  wire  _hit_T = |hitVec; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 210:35]
  wire  hit = io_in_valid & |hitVec; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 210:25]
  wire  miss = io_in_valid & ~_hit_T; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 211:26]
  reg [63:0] victimWaymask_lfsr; // @[src/main/scala/utils/LFSR64.scala 25:23]
  wire  victimWaymask_xor = victimWaymask_lfsr[0] ^ victimWaymask_lfsr[1] ^ victimWaymask_lfsr[3] ^ victimWaymask_lfsr[4
    ]; // @[src/main/scala/utils/LFSR64.scala 26:43]
  wire [63:0] _victimWaymask_lfsr_T_2 = {victimWaymask_xor,victimWaymask_lfsr[63:1]}; // @[src/main/scala/utils/LFSR64.scala 28:41]
  wire [3:0] victimWaymask = 4'h1 << victimWaymask_lfsr[1:0]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 213:42]
  wire [3:0] waymask = hit ? hitVec : victimWaymask; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 214:20]
  wire [120:0] _hitMeta_T_4 = waymask[0] ? io_md_0 : 121'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [120:0] _hitMeta_T_5 = waymask[1] ? io_md_1 : 121'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [120:0] _hitMeta_T_6 = waymask[2] ? io_md_2 : 121'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [120:0] _hitMeta_T_7 = waymask[3] ? io_md_3 : 121'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [120:0] _hitMeta_T_8 = _hitMeta_T_4 | _hitMeta_T_5; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [120:0] _hitMeta_T_9 = _hitMeta_T_8 | _hitMeta_T_6; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [120:0] _hitMeta_T_10 = _hitMeta_T_9 | _hitMeta_T_7; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [7:0] hitMeta_flag = _hitMeta_T_10[59:52]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 220:70]
  wire [17:0] hitMeta_mask = _hitMeta_T_10[77:60]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 220:70]
  wire [15:0] hitMeta_asid = _hitMeta_T_10[93:78]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 220:70]
  wire [26:0] hitMeta_vpn = _hitMeta_T_10[120:94]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 220:70]
  wire [31:0] hitData_pteaddr = _hitMeta_T_10[31:0]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:70]
  wire [19:0] hitData_ppn = _hitMeta_T_10[51:32]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:70]
  wire  hitFlag_v = hitMeta_flag[0]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 222:38]
  wire  hitFlag_r = hitMeta_flag[1]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 222:38]
  wire  hitFlag_w = hitMeta_flag[2]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 222:38]
  wire  hitFlag_x = hitMeta_flag[3]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 222:38]
  wire  hitFlag_u = hitMeta_flag[4]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 222:38]
  wire  hitFlag_g = hitMeta_flag[5]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 222:38]
  wire  hitFlag_a = hitMeta_flag[6]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 222:38]
  wire  hitFlag_d = hitMeta_flag[7]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 222:38]
  wire  _hitWB_T_4 = ~hitFlag_a | ~hitFlag_d & io_in_bits_cmd[0]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 226:34]
  reg [2:0] state; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 253:22]
  wire  _T_4 = 3'h0 == state; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 275:18]
  wire  _hitCheck_T = io_pf_priviledgeMode == 2'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 231:62]
  wire  _hitCheck_T_5 = io_pf_priviledgeMode == 2'h1; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 231:110]
  wire  _hitCheck_T_7 = ~io_pf_status_sum; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 231:137]
  wire  hitCheck = hit & ~(io_pf_priviledgeMode == 2'h0 & ~hitFlag_u) & ~(io_pf_priviledgeMode == 2'h1 & hitFlag_u & ~
    io_pf_status_sum); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 231:87]
  wire  _hitLoad_T_1 = hitCheck & ~_hitWB_T_4; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 234:26]
  wire  hitLoad = hitCheck & ~_hitWB_T_4 & (hitFlag_r | io_pf_status_mxr & hitFlag_x); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 234:41]
  wire  _loadPF_T_5 = ~io_in_bits_cmd[0] & ~io_in_bits_cmd[3]; // @[src/main/scala/bus/simplebus/SimpleBus.scala 73:26]
  wire  _loadPF_T_7 = ~hitLoad & _loadPF_T_5 & hit; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 247:40]
  wire  _loadPF_T_8 = ~ISAMO; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 247:50]
  wire  _T_9 = 3'h1 == state; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 275:18]
  wire  _T_11 = 3'h2 == state; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 275:18]
  wire  _T_12 = io_mem_resp_ready & io_mem_resp_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  wire  memRdata_flag_d = io_mem_resp_bits_rdata[7]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 261:49]
  wire  memRdata_flag_a = io_mem_resp_bits_rdata[6]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 261:49]
  wire  memRdata_flag_g = io_mem_resp_bits_rdata[5]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 261:49]
  wire  memRdata_flag_u = io_mem_resp_bits_rdata[4]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 261:49]
  wire  memRdata_flag_x = io_mem_resp_bits_rdata[3]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 261:49]
  wire  memRdata_flag_w = io_mem_resp_bits_rdata[2]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 261:49]
  wire  memRdata_flag_r = io_mem_resp_bits_rdata[1]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 261:49]
  wire  memRdata_flag_v = io_mem_resp_bits_rdata[0]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 261:49]
  wire [7:0] _missflag_T = {memRdata_flag_d,memRdata_flag_a,memRdata_flag_g,memRdata_flag_u,memRdata_flag_x,
    memRdata_flag_w,memRdata_flag_r,memRdata_flag_v}; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 298:44]
  wire  missflag_r = _missflag_T[1]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 298:44]
  wire  missflag_x = _missflag_T[3]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 298:44]
  reg [1:0] level; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 254:22]
  wire  _T_15 = level == 2'h3; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 303:58]
  wire  _T_16 = level == 2'h2; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 303:73]
  wire  _T_18 = ~(missflag_r | missflag_x) & (level == 2'h3 | level == 2'h2); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 303:49]
  wire  missflag_v = _missflag_T[0]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 298:44]
  wire  missflag_w = _missflag_T[2]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 298:44]
  wire  _T_22 = ~missflag_v | ~missflag_r & missflag_w; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 304:28]
  wire  _loadPF_T_16 = _loadPF_T_5 & _loadPF_T_8; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 308:38]
  wire  _GEN_19 = ~missflag_v | ~missflag_r & missflag_w ? _loadPF_T_5 & _loadPF_T_8 : ~hitLoad & _loadPF_T_5 & hit & ~
    ISAMO; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 247:12 304:60 308:22]
  wire  missflag_u = _missflag_T[4]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 298:44]
  wire  permCheck = missflag_v & ~(_hitCheck_T & ~missflag_u) & ~(_hitCheck_T_5 & missflag_u & _hitCheck_T_7); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 320:87]
  wire  missflag_a = _missflag_T[6]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 298:44]
  wire  missflag_d = _missflag_T[7]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 298:44]
  wire  permAD = ~missflag_a | ~missflag_d & io_in_bits_cmd[0]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 321:83]
  wire  _permLoad_T_1 = permCheck & ~permAD; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 323:36]
  wire  permLoad = permCheck & ~permAD & (missflag_r | io_pf_status_mxr & missflag_x); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 323:47]
  wire  permStore = _permLoad_T_1 & missflag_w; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 324:48]
  wire  _GEN_23 = ~permLoad & _loadPF_T_5 | ~permStore & io_in_bits_cmd[0] ? _loadPF_T_16 : ~hitLoad & _loadPF_T_5 & hit
     & ~ISAMO; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 247:12 337:80 339:22]
  wire  _GEN_29 = level != 2'h0 ? _GEN_23 : ~hitLoad & _loadPF_T_5 & hit & ~ISAMO; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 247:12 319:36]
  wire  _GEN_35 = ~(missflag_r | missflag_x) & (level == 2'h3 | level == 2'h2) ? _GEN_19 : _GEN_29; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 303:82]
  wire  _GEN_54 = _T_12 ? _GEN_35 : ~hitLoad & _loadPF_T_5 & hit & ~ISAMO; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 247:12 299:31]
  wire  _GEN_78 = 3'h2 == state ? _GEN_54 : ~hitLoad & _loadPF_T_5 & hit & ~ISAMO; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 247:12 275:18]
  wire  _GEN_91 = 3'h1 == state ? ~hitLoad & _loadPF_T_5 & hit & ~ISAMO : _GEN_78; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 247:12 275:18]
  wire  loadPF = 3'h0 == state ? ~hitLoad & _loadPF_T_5 & hit & ~ISAMO : _GEN_91; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 247:12 275:18]
  wire  hitStore = _hitLoad_T_1 & hitFlag_w; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 235:42]
  wire  _storePF_T_15 = io_in_bits_cmd[0] | ISAMO; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 309:40]
  wire  _GEN_20 = ~missflag_v | ~missflag_r & missflag_w ? io_in_bits_cmd[0] | ISAMO : ~hitStore & io_in_bits_cmd[0] &
    hit | _loadPF_T_7 & ISAMO; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 248:13 304:60 309:23]
  wire  _GEN_24 = ~permLoad & _loadPF_T_5 | ~permStore & io_in_bits_cmd[0] ? _storePF_T_15 : ~hitStore & io_in_bits_cmd[
    0] & hit | _loadPF_T_7 & ISAMO; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 248:13 337:80 340:23]
  wire  _GEN_30 = level != 2'h0 ? _GEN_24 : ~hitStore & io_in_bits_cmd[0] & hit | _loadPF_T_7 & ISAMO; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 248:13 319:36]
  wire  _GEN_36 = ~(missflag_r | missflag_x) & (level == 2'h3 | level == 2'h2) ? _GEN_20 : _GEN_30; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 303:82]
  wire  _GEN_55 = _T_12 ? _GEN_36 : ~hitStore & io_in_bits_cmd[0] & hit | _loadPF_T_7 & ISAMO; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 248:13 299:31]
  wire  _GEN_79 = 3'h2 == state ? _GEN_55 : ~hitStore & io_in_bits_cmd[0] & hit | _loadPF_T_7 & ISAMO; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 248:13 275:18]
  wire  _GEN_92 = 3'h1 == state ? ~hitStore & io_in_bits_cmd[0] & hit | _loadPF_T_7 & ISAMO : _GEN_79; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 248:13 275:18]
  wire  storePF = 3'h0 == state ? ~hitStore & io_in_bits_cmd[0] & hit | _loadPF_T_7 & ISAMO : _GEN_92; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 248:13 275:18]
  wire  _hitWB_T_9 = io_pf_loadPF | io_pf_storePF; // @[src/main/scala/nutcore/Bundle.scala 131:23]
  wire  hitWB = hit & (~hitFlag_a | ~hitFlag_d & io_in_bits_cmd[0]) & ~(loadPF | storePF | _hitWB_T_9); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 226:81]
  wire [7:0] _hitRefillFlag_T_1 = {io_in_bits_cmd[0],1'h1,6'h0}; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 227:26]
  wire [7:0] _hitRefillFlag_T_2 = {hitFlag_d,hitFlag_a,hitFlag_g,hitFlag_u,hitFlag_x,hitFlag_w,hitFlag_r,hitFlag_v}; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 227:79]
  wire [7:0] hitRefillFlag = _hitRefillFlag_T_1 | _hitRefillFlag_T_2; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 227:69]
  wire [39:0] _hitWBStore_T = {10'h0,hitData_ppn,2'h0,hitRefillFlag}; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 228:33]
  reg [39:0] hitWBStore; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 228:29]
  wire  hitExec = _hitLoad_T_1 & hitFlag_x; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 233:41]
  reg  io_pf_loadPF_REG; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 242:26]
  reg  io_pf_storePF_REG; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 243:27]
  reg [63:0] memRespStore; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 256:25]
  reg [17:0] missMaskStore; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 258:26]
  wire [1:0] memRdata_rsw = io_mem_resp_bits_rdata[9:8]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 261:49]
  wire [19:0] memRdata_ppn = io_mem_resp_bits_rdata[29:10]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 261:49]
  wire [33:0] memRdata_reserved = io_mem_resp_bits_rdata[63:30]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 261:49]
  reg [31:0] raddr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 262:18]
  wire  _alreadyOutFire_T = io_out_ready & io_out_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  reg  alreadyOutFire; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 263:33]
  wire  _GEN_2 = _alreadyOutFire_T | alreadyOutFire; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 263:{33,33,33}]
  wire [31:0] _raddr_T_1 = {satp_ppn,vpn_vpn2,3'h0}; // @[src/main/scala/nutcore/mem/TLB.scala 89:8]
  wire  _T_10 = io_mem_req_ready & io_mem_req_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  wire  missflag_g = _missflag_T[5]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 298:44]
  reg [63:0] c; // @[src/main/scala/utils/GTimer.scala 24:20]
  wire [63:0] _c_T_1 = c + 64'h1; // @[src/main/scala/utils/GTimer.scala 25:12]
  wire  _T_25 = ~reset; // @[src/main/scala/utils/Debug.scala 56:24]
  wire [8:0] _raddr_T_3 = _T_15 ? vpn_vpn1 : vpn_vpn0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 317:50]
  wire [31:0] _raddr_T_5 = {memRdata_ppn,_raddr_T_3,3'h0}; // @[src/main/scala/nutcore/mem/TLB.scala 89:8]
  wire [2:0] _GEN_18 = ~missflag_v | ~missflag_r & missflag_w ? 3'h5 : 3'h1; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 304:60 305:73 316:19]
  wire [31:0] _GEN_21 = ~missflag_v | ~missflag_r & missflag_w ? raddr : _raddr_T_5; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 262:18 304:60 317:19]
  wire [63:0] updateData = {56'h0,io_in_bits_cmd[0],7'h40}; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 326:31]
  wire [7:0] _missRefillFlag_T_2 = {missflag_d,missflag_a,missflag_g,missflag_u,missflag_x,missflag_w,missflag_r,
    missflag_v}; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 327:79]
  wire [7:0] _missRefillFlag_T_3 = _hitRefillFlag_T_1 | _missRefillFlag_T_2; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 327:68]
  wire [63:0] _memRespStore_T = io_mem_resp_bits_rdata | updateData; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 328:50]
  wire [2:0] _GEN_22 = ~permLoad & _loadPF_T_5 | ~permStore & io_in_bits_cmd[0] ? 3'h5 : 3'h4; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 337:80 338:21 342:21]
  wire  _GEN_25 = ~permLoad & _loadPF_T_5 | ~permStore & io_in_bits_cmd[0] ? 1'h0 : 1'h1; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 259:32 337:80 343:30]
  wire [17:0] _missMask_T_2 = _T_16 ? 18'h3fe00 : 18'h3ffff; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 346:59]
  wire [17:0] _missMask_T_3 = _T_15 ? 18'h0 : _missMask_T_2; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 346:26]
  wire [7:0] _GEN_26 = level != 2'h0 ? _missRefillFlag_T_3 : 8'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 319:36 327:26 260:32]
  wire [63:0] _GEN_27 = level != 2'h0 ? _memRespStore_T : memRespStore; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 319:36 328:24 256:25]
  wire [2:0] _GEN_28 = level != 2'h0 ? _GEN_22 : state; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 253:22 319:36]
  wire  _GEN_31 = level != 2'h0 & _GEN_25; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 259:32 319:36]
  wire [17:0] _GEN_32 = level != 2'h0 ? _missMask_T_3 : 18'h3ffff; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 319:36 346:20 257:26]
  wire [17:0] _GEN_41 = ~(missflag_r | missflag_x) & (level == 2'h3 | level == 2'h2) ? 18'h3ffff : _GEN_32; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 257:26 303:82]
  wire [17:0] _GEN_60 = _T_12 ? _GEN_41 : 18'h3ffff; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 257:26 299:31]
  wire [17:0] _GEN_84 = 3'h2 == state ? _GEN_60 : 18'h3ffff; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 275:18 257:26]
  wire [17:0] _GEN_97 = 3'h1 == state ? 18'h3ffff : _GEN_84; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 275:18 257:26]
  wire [17:0] missMask = 3'h0 == state ? 18'h3ffff : _GEN_97; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 275:18 257:26]
  wire [17:0] _GEN_33 = level != 2'h0 ? missMask : missMaskStore; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 319:36 347:25 258:26]
  wire [2:0] _GEN_34 = ~(missflag_r | missflag_x) & (level == 2'h3 | level == 2'h2) ? _GEN_18 : _GEN_28; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 303:82]
  wire [31:0] _GEN_37 = ~(missflag_r | missflag_x) & (level == 2'h3 | level == 2'h2) ? _GEN_21 : raddr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 262:18 303:82]
  wire [7:0] _GEN_38 = ~(missflag_r | missflag_x) & (level == 2'h3 | level == 2'h2) ? 8'h0 : _GEN_26; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 260:32 303:82]
  wire [63:0] _GEN_39 = ~(missflag_r | missflag_x) & (level == 2'h3 | level == 2'h2) ? memRespStore : _GEN_27; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 256:25 303:82]
  wire  _GEN_40 = ~(missflag_r | missflag_x) & (level == 2'h3 | level == 2'h2) ? 1'h0 : _GEN_31; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 259:32 303:82]
  wire [17:0] _GEN_42 = ~(missflag_r | missflag_x) & (level == 2'h3 | level == 2'h2) ? missMaskStore : _GEN_33; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 258:26 303:82]
  wire [1:0] _level_T_1 = level - 2'h1; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 349:24]
  wire [2:0] _GEN_52 = _T_12 ? _GEN_34 : state; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 253:22 299:31]
  wire [7:0] _GEN_57 = _T_12 ? _GEN_38 : 8'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 299:31 260:32]
  wire  _GEN_59 = _T_12 & _GEN_40; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 299:31 259:32]
  wire [1:0] _GEN_62 = _T_12 ? _level_T_1 : level; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 299:31 349:15 254:22]
  wire [2:0] _GEN_63 = _T_10 ? 3'h4 : state; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 253:22 357:{36,44}]
  wire [2:0] _GEN_65 = _GEN_2 ? 3'h0 : state; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 360:71 361:13 253:22]
  wire  _GEN_67 = _GEN_2 ? 1'h0 : _GEN_2; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 360:71 363:22]
  wire [2:0] _GEN_68 = 3'h5 == state ? 3'h0 : state; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 275:18 367:13 253:22]
  wire [2:0] _GEN_69 = 3'h4 == state ? _GEN_65 : _GEN_68; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 275:18]
  wire  _GEN_71 = 3'h4 == state ? _GEN_67 : _GEN_2; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 275:18]
  wire [2:0] _GEN_72 = 3'h3 == state ? _GEN_63 : _GEN_69; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 275:18]
  wire  _GEN_75 = 3'h3 == state ? _GEN_2 : _GEN_71; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 275:18]
  wire [7:0] _GEN_81 = 3'h2 == state ? _GEN_57 : 8'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 275:18 260:32]
  wire [7:0] _GEN_94 = 3'h1 == state ? 8'h0 : _GEN_81; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 275:18 260:32]
  wire  _GEN_96 = 3'h1 == state ? 1'h0 : 3'h2 == state & _GEN_59; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 275:18 259:32]
  wire [7:0] missRefillFlag = 3'h0 == state ? 8'h0 : _GEN_94; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 275:18 260:32]
  wire  missMetaRefill = 3'h0 == state ? 1'h0 : _GEN_96; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 275:18 259:32]
  wire  cmd = state == 3'h3; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 372:23]
  wire  _T_60 = state == 3'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 378:82]
  reg  REG; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 378:33]
  reg [3:0] REG_1; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 379:21]
  reg [3:0] REG_2; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 379:60]
  reg [26:0] REG_3; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 379:84]
  reg [15:0] REG_4; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 380:19]
  reg [17:0] REG_5; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 380:72]
  reg [7:0] REG_6; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 381:19]
  reg [19:0] REG_7; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 381:77]
  reg [31:0] REG_8; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 382:22]
  wire [59:0] io_mdWrite_wdata_lo = {REG_6,REG_7,REG_8}; // @[src/main/scala/nutcore/mem/TLB.scala 217:22]
  wire [60:0] io_mdWrite_wdata_hi = {REG_3,REG_4,REG_5}; // @[src/main/scala/nutcore/mem/TLB.scala 217:22]
  wire [31:0] _io_out_bits_addr_T_1 = {hitData_ppn,12'h0}; // @[src/main/scala/nutcore/mem/TLB.scala 127:24]
  wire [31:0] _io_out_bits_addr_T_3 = {2'h3,hitMeta_mask,12'h0}; // @[src/main/scala/nutcore/mem/TLB.scala 127:49]
  wire [31:0] _io_out_bits_addr_T_4 = _io_out_bits_addr_T_1 & _io_out_bits_addr_T_3; // @[src/main/scala/utils/BitUtils.scala 34:14]
  wire [31:0] _io_out_bits_addr_T_5 = ~_io_out_bits_addr_T_3; // @[src/main/scala/utils/BitUtils.scala 34:39]
  wire [31:0] _io_out_bits_addr_T_6 = io_in_bits_addr[31:0] & _io_out_bits_addr_T_5; // @[src/main/scala/utils/BitUtils.scala 34:37]
  wire [31:0] _io_out_bits_addr_T_7 = _io_out_bits_addr_T_4 | _io_out_bits_addr_T_6; // @[src/main/scala/utils/BitUtils.scala 34:26]
  wire [31:0] _io_out_bits_addr_T_20 = {memRespStore[29:10],12'h0}; // @[src/main/scala/nutcore/mem/TLB.scala 127:24]
  wire [31:0] _io_out_bits_addr_T_22 = {2'h3,missMaskStore,12'h0}; // @[src/main/scala/nutcore/mem/TLB.scala 127:49]
  wire [31:0] _io_out_bits_addr_T_23 = _io_out_bits_addr_T_20 & _io_out_bits_addr_T_22; // @[src/main/scala/utils/BitUtils.scala 34:14]
  wire [31:0] _io_out_bits_addr_T_24 = ~_io_out_bits_addr_T_22; // @[src/main/scala/utils/BitUtils.scala 34:39]
  wire [31:0] _io_out_bits_addr_T_25 = io_in_bits_addr[31:0] & _io_out_bits_addr_T_24; // @[src/main/scala/utils/BitUtils.scala 34:37]
  wire [31:0] _io_out_bits_addr_T_26 = _io_out_bits_addr_T_23 | _io_out_bits_addr_T_25; // @[src/main/scala/utils/BitUtils.scala 34:26]
  wire  _io_out_valid_T = ~hitWB; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 387:45]
  wire  _io_out_valid_T_7 = hit & ~hitWB ? ~(_hitWB_T_9 | loadPF | storePF) : state == 3'h4; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 387:37]
  reg [63:0] c_4; // @[src/main/scala/utils/GTimer.scala 24:20]
  wire [63:0] _c_T_9 = c_4 + 64'h1; // @[src/main/scala/utils/GTimer.scala 25:12]
  reg [63:0] c_5; // @[src/main/scala/utils/GTimer.scala 24:20]
  wire [63:0] _c_T_11 = c_5 + 64'h1; // @[src/main/scala/utils/GTimer.scala 25:12]
  reg [63:0] c_6; // @[src/main/scala/utils/GTimer.scala 24:20]
  wire [63:0] _c_T_13 = c_6 + 64'h1; // @[src/main/scala/utils/GTimer.scala 25:12]
  wire [4:0] lo_1 = {memRdata_flag_u,memRdata_flag_x,memRdata_flag_w,memRdata_flag_r,memRdata_flag_v}; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 397:145]
  wire [63:0] _T_90 = {memRdata_reserved,memRdata_ppn,memRdata_rsw,memRdata_flag_d,memRdata_flag_a,memRdata_flag_g,lo_1}
    ; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 397:145]
  reg [63:0] c_7; // @[src/main/scala/utils/GTimer.scala 24:20]
  wire [63:0] _c_T_15 = c_7 + 64'h1; // @[src/main/scala/utils/GTimer.scala 25:12]
  reg [63:0] c_8; // @[src/main/scala/utils/GTimer.scala 24:20]
  wire [63:0] _c_T_17 = c_8 + 64'h1; // @[src/main/scala/utils/GTimer.scala 25:12]
  reg [63:0] c_9; // @[src/main/scala/utils/GTimer.scala 24:20]
  wire [63:0] _c_T_19 = c_9 + 64'h1; // @[src/main/scala/utils/GTimer.scala 25:12]
  reg [63:0] c_10; // @[src/main/scala/utils/GTimer.scala 24:20]
  wire [63:0] _c_T_21 = c_10 + 64'h1; // @[src/main/scala/utils/GTimer.scala 25:12]
  reg [63:0] c_11; // @[src/main/scala/utils/GTimer.scala 24:20]
  wire [63:0] _c_T_23 = c_11 + 64'h1; // @[src/main/scala/utils/GTimer.scala 25:12]
  wire  _GEN_122 = ~_T_4 & ~_T_9 & _T_11 & _T_12 & _T_18 & _T_22 & DISPLAY_ENABLE; // @[src/main/scala/utils/Debug.scala 56:24]
  assign io_in_ready = io_out_ready & _T_60 & ~miss & _io_out_valid_T & io_mdReady & (~_hitWB_T_9 & ~loadPF & ~storePF); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 389:86]
  assign io_out_valid = io_in_valid & _io_out_valid_T_7; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 387:31]
  assign io_out_bits_addr = hit ? _io_out_bits_addr_T_7 : _io_out_bits_addr_T_26; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 386:26]
  assign io_out_bits_size = io_in_bits_size; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 385:15]
  assign io_out_bits_cmd = io_in_bits_cmd; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 385:15]
  assign io_out_bits_wmask = io_in_bits_wmask; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 385:15]
  assign io_out_bits_wdata = io_in_bits_wdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 385:15]
  assign io_mdWrite_wen = REG; // @[src/main/scala/nutcore/mem/TLB.scala 214:14]
  assign io_mdWrite_windex = REG_1; // @[src/main/scala/nutcore/mem/TLB.scala 215:17]
  assign io_mdWrite_waymask = REG_2; // @[src/main/scala/nutcore/mem/TLB.scala 216:18]
  assign io_mdWrite_wdata = {io_mdWrite_wdata_hi,io_mdWrite_wdata_lo}; // @[src/main/scala/nutcore/mem/TLB.scala 217:22]
  assign io_mem_req_valid = state == 3'h1 | cmd; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 374:48]
  assign io_mem_req_bits_addr = hitWB ? hitData_pteaddr : raddr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 373:35]
  assign io_mem_req_bits_size = 3'h3; // @[src/main/scala/bus/simplebus/SimpleBus.scala 66:15]
  assign io_mem_req_bits_cmd = {{3'd0}, cmd}; // @[src/main/scala/bus/simplebus/SimpleBus.scala 65:14]
  assign io_mem_req_bits_wmask = 8'hff; // @[src/main/scala/bus/simplebus/SimpleBus.scala 68:16]
  assign io_mem_req_bits_wdata = hitWB ? {{24'd0}, hitWBStore} : memRespStore; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 373:138]
  assign io_mem_resp_ready = 1'h1; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 375:21]
  assign io_pf_loadPF = io_pf_loadPF_REG; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 242:16]
  assign io_pf_storePF = io_pf_storePF_REG; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 243:17]
  assign io_pf_addr = io_in_bits_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 206:11]
  assign io_ipf = 1'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 391:16]
  assign io_isFinish = _alreadyOutFire_T | _hitWB_T_9; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 392:30]
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/utils/LFSR64.scala 25:23]
      victimWaymask_lfsr <= 64'h1234567887654321; // @[src/main/scala/utils/LFSR64.scala 25:23]
    end else if (victimWaymask_lfsr == 64'h0) begin // @[src/main/scala/utils/LFSR64.scala 28:18]
      victimWaymask_lfsr <= 64'h1;
    end else begin
      victimWaymask_lfsr <= _victimWaymask_lfsr_T_2;
    end
    if (reset) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 253:22]
      state <= 3'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 253:22]
    end else if (3'h0 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 275:18]
      if (hitWB) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 277:32]
        state <= 3'h3; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 278:15]
      end else if (miss) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 281:37]
        state <= 3'h1; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 282:15]
      end
    end else if (3'h1 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 275:18]
      if (_T_10) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 294:36]
        state <= 3'h2; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 294:44]
      end
    end else if (3'h2 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 275:18]
      state <= _GEN_52;
    end else begin
      state <= _GEN_72;
    end
    if (reset) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 254:22]
      level <= 2'h3; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 254:22]
    end else if (3'h0 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 275:18]
      if (!(hitWB)) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 277:32]
        if (miss) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 281:37]
          level <= 2'h3; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 284:15]
        end
      end
    end else if (!(3'h1 == state)) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 275:18]
      if (3'h2 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 275:18]
        level <= _GEN_62;
      end
    end
    if (hitWB) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 228:29]
      hitWBStore <= _hitWBStore_T; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 228:29]
    end
    if (reset) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 242:26]
      io_pf_loadPF_REG <= 1'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 242:26]
    end else if (3'h0 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 275:18]
      io_pf_loadPF_REG <= ~hitLoad & _loadPF_T_5 & hit & ~ISAMO; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 247:12]
    end else if (3'h1 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 275:18]
      io_pf_loadPF_REG <= ~hitLoad & _loadPF_T_5 & hit & ~ISAMO; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 247:12]
    end else if (3'h2 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 275:18]
      io_pf_loadPF_REG <= _GEN_54;
    end else begin
      io_pf_loadPF_REG <= ~hitLoad & _loadPF_T_5 & hit & ~ISAMO; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 247:12]
    end
    if (reset) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 243:27]
      io_pf_storePF_REG <= 1'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 243:27]
    end else if (3'h0 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 275:18]
      io_pf_storePF_REG <= ~hitStore & io_in_bits_cmd[0] & hit | _loadPF_T_7 & ISAMO; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 248:13]
    end else if (3'h1 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 275:18]
      io_pf_storePF_REG <= ~hitStore & io_in_bits_cmd[0] & hit | _loadPF_T_7 & ISAMO; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 248:13]
    end else if (3'h2 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 275:18]
      io_pf_storePF_REG <= _GEN_55;
    end else begin
      io_pf_storePF_REG <= ~hitStore & io_in_bits_cmd[0] & hit | _loadPF_T_7 & ISAMO; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 248:13]
    end
    if (!(3'h0 == state)) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 275:18]
      if (!(3'h1 == state)) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 275:18]
        if (3'h2 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 275:18]
          if (_T_12) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 299:31]
            memRespStore <= _GEN_39;
          end
        end
      end
    end
    if (!(3'h0 == state)) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 275:18]
      if (!(3'h1 == state)) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 275:18]
        if (3'h2 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 275:18]
          if (_T_12) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 299:31]
            missMaskStore <= _GEN_42;
          end
        end
      end
    end
    if (3'h0 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 275:18]
      if (!(hitWB)) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 277:32]
        if (miss) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 281:37]
          raddr <= _raddr_T_1; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 283:15]
        end
      end
    end else if (!(3'h1 == state)) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 275:18]
      if (3'h2 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 275:18]
        if (_T_12) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 299:31]
          raddr <= _GEN_37;
        end
      end
    end
    if (reset) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 263:33]
      alreadyOutFire <= 1'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 263:33]
    end else if (3'h0 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 275:18]
      if (hitWB) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 277:32]
        alreadyOutFire <= 1'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 280:24]
      end else if (miss) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 281:37]
        alreadyOutFire <= 1'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 286:24]
      end else begin
        alreadyOutFire <= _GEN_2;
      end
    end else if (3'h1 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 275:18]
      alreadyOutFire <= _GEN_2;
    end else if (3'h2 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 275:18]
      alreadyOutFire <= _GEN_2;
    end else begin
      alreadyOutFire <= _GEN_75;
    end
    if (reset) begin // @[src/main/scala/utils/GTimer.scala 24:20]
      c <= 64'h0; // @[src/main/scala/utils/GTimer.scala 24:20]
    end else begin
      c <= _c_T_1; // @[src/main/scala/utils/GTimer.scala 25:7]
    end
    if (reset) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 378:33]
      REG <= 1'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 378:33]
    end else begin
      REG <= missMetaRefill | hitWB & state == 3'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 378:33]
    end
    REG_1 <= io_in_bits_addr[15:12]; // @[src/main/scala/nutcore/mem/TLB.scala 200:19]
    if (hit) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 214:20]
      REG_2 <= hitVec;
    end else begin
      REG_2 <= victimWaymask;
    end
    REG_3 <= {hitVec_hi,vpn_vpn0}; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 379:89]
    if (hitWB) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 380:23]
      REG_4 <= hitMeta_asid;
    end else begin
      REG_4 <= satp_asid;
    end
    if (hitWB) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 380:76]
      REG_5 <= hitMeta_mask;
    end else if (3'h0 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 275:18]
      REG_5 <= 18'h3ffff; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 257:26]
    end else if (3'h1 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 275:18]
      REG_5 <= 18'h3ffff; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 257:26]
    end else if (3'h2 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 275:18]
      REG_5 <= _GEN_60;
    end else begin
      REG_5 <= 18'h3ffff; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 257:26]
    end
    if (hitWB) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 381:23]
      REG_6 <= hitRefillFlag;
    end else if (3'h0 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 275:18]
      REG_6 <= 8'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 260:32]
    end else if (3'h1 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 275:18]
      REG_6 <= 8'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 260:32]
    end else if (3'h2 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 275:18]
      REG_6 <= _GEN_57;
    end else begin
      REG_6 <= 8'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 260:32]
    end
    if (hitWB) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 381:81]
      REG_7 <= hitData_ppn;
    end else begin
      REG_7 <= memRdata_ppn;
    end
    if (hitWB) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 382:27]
      REG_8 <= hitData_pteaddr;
    end else begin
      REG_8 <= raddr;
    end
    if (reset) begin // @[src/main/scala/utils/GTimer.scala 24:20]
      c_4 <= 64'h0; // @[src/main/scala/utils/GTimer.scala 24:20]
    end else begin
      c_4 <= _c_T_9; // @[src/main/scala/utils/GTimer.scala 25:7]
    end
    if (reset) begin // @[src/main/scala/utils/GTimer.scala 24:20]
      c_5 <= 64'h0; // @[src/main/scala/utils/GTimer.scala 24:20]
    end else begin
      c_5 <= _c_T_11; // @[src/main/scala/utils/GTimer.scala 25:7]
    end
    if (reset) begin // @[src/main/scala/utils/GTimer.scala 24:20]
      c_6 <= 64'h0; // @[src/main/scala/utils/GTimer.scala 24:20]
    end else begin
      c_6 <= _c_T_13; // @[src/main/scala/utils/GTimer.scala 25:7]
    end
    if (reset) begin // @[src/main/scala/utils/GTimer.scala 24:20]
      c_7 <= 64'h0; // @[src/main/scala/utils/GTimer.scala 24:20]
    end else begin
      c_7 <= _c_T_15; // @[src/main/scala/utils/GTimer.scala 25:7]
    end
    if (reset) begin // @[src/main/scala/utils/GTimer.scala 24:20]
      c_8 <= 64'h0; // @[src/main/scala/utils/GTimer.scala 24:20]
    end else begin
      c_8 <= _c_T_17; // @[src/main/scala/utils/GTimer.scala 25:7]
    end
    if (reset) begin // @[src/main/scala/utils/GTimer.scala 24:20]
      c_9 <= 64'h0; // @[src/main/scala/utils/GTimer.scala 24:20]
    end else begin
      c_9 <= _c_T_19; // @[src/main/scala/utils/GTimer.scala 25:7]
    end
    if (reset) begin // @[src/main/scala/utils/GTimer.scala 24:20]
      c_10 <= 64'h0; // @[src/main/scala/utils/GTimer.scala 24:20]
    end else begin
      c_10 <= _c_T_21; // @[src/main/scala/utils/GTimer.scala 25:7]
    end
    if (reset) begin // @[src/main/scala/utils/GTimer.scala 24:20]
      c_11 <= 64'h0; // @[src/main/scala/utils/GTimer.scala 24:20]
    end else begin
      c_11 <= _c_T_23; // @[src/main/scala/utils/GTimer.scala 25:7]
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~_T_4 & ~_T_9 & _T_11 & _T_12 & _T_18 & _T_22 & DISPLAY_ENABLE & ~reset) begin
          $fwrite(32'h80000002,"[%d] EmbeddedTLBExec_1: ",c); // @[src/main/scala/utils/Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_122 & _T_25) begin
          $fwrite(32'h80000002,"tlbException!!! "); // @[src/main/scala/utils/Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_122 & _T_25) begin
          $fwrite(32'h80000002,
            " req:addr = 0x%x, cmd = %d, size = %d, wmask = 0x%x, wdata = 0x%x  Memreq:DecoupledIO(ready -> %d, valid -> %d, bits -> addr = 0x%x, cmd = %d, size = %d, wmask = 0x%x, wdata = 0x%x)  MemResp:DecoupledIO(ready -> %d, valid -> %d, bits -> rdata = %x, cmd = %d)"
            ,io_in_bits_addr,io_in_bits_cmd,io_in_bits_size,io_in_bits_wmask,io_in_bits_wdata,io_mem_req_ready,
            io_mem_req_valid,io_mem_req_bits_addr,io_mem_req_bits_cmd,io_mem_req_bits_size,io_mem_req_bits_wmask,
            io_mem_req_bits_wdata,io_mem_resp_ready,io_mem_resp_valid,io_mem_resp_bits_rdata,io_mem_resp_bits_cmd); // @[src/main/scala/utils/Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_122 & _T_25) begin
          $fwrite(32'h80000002," level:%d",level); // @[src/main/scala/utils/Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_122 & _T_25) begin
          $fwrite(32'h80000002,"\n"); // @[src/main/scala/utils/Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & ~reset) begin
          $fwrite(32'h80000002,"[%d] EmbeddedTLBExec_1: ",c_4); // @[src/main/scala/utils/Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_25) begin
          $fwrite(32'h80000002,"In(%d, %d) Out(%d, %d) InAddr:%x OutAddr:%x cmd:%d \n",io_in_valid,io_in_ready,
            io_out_valid,io_out_ready,io_in_bits_addr,io_out_bits_addr,io_in_bits_cmd); // @[src/main/scala/utils/Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & ~reset) begin
          $fwrite(32'h80000002,"[%d] EmbeddedTLBExec_1: ",c_5); // @[src/main/scala/utils/Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_25) begin
          $fwrite(32'h80000002,"isAMO:%d io.Flush:%d needFlush:%d alreadyOutFire:%d isFinish:%d\n",ISAMO,1'h0,1'h0,
            alreadyOutFire,io_isFinish); // @[src/main/scala/utils/Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & ~reset) begin
          $fwrite(32'h80000002,"[%d] EmbeddedTLBExec_1: ",c_6); // @[src/main/scala/utils/Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_25) begin
          $fwrite(32'h80000002,
            "hit:%d hitWB:%d hitVPN:%x hitFlag:%x hitPPN:%x hitRefillFlag:%x hitWBStore:%x hitCheck:%d hitExec:%d hitLoad:%d hitStore:%d\n"
            ,hit,hitWB,hitMeta_vpn,_hitRefillFlag_T_2,hitData_ppn,hitRefillFlag,hitWBStore,hitCheck,hitExec,hitLoad,
            hitStore); // @[src/main/scala/utils/Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & ~reset) begin
          $fwrite(32'h80000002,"[%d] EmbeddedTLBExec_1: ",c_7); // @[src/main/scala/utils/Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_25) begin
          $fwrite(32'h80000002,
            "miss:%d state:%d level:%d raddr:%x memRdata:%x missMask:%x missRefillFlag:%x missMetaRefill:%d\n",miss,
            state,level,raddr,_T_90,missMask,missRefillFlag,missMetaRefill); // @[src/main/scala/utils/Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & ~reset) begin
          $fwrite(32'h80000002,"[%d] EmbeddedTLBExec_1: ",c_8); // @[src/main/scala/utils/Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_25) begin
          $fwrite(32'h80000002,"meta/data: (0)%x|%b|%x (1)%x|%b|%x (2)%x|%b|%x (3)%x|%b|%x rread:%d\n",io_md_0[120:94],
            io_md_0[59:52],io_md_0[51:32],io_md_1[120:94],io_md_1[59:52],io_md_1[51:32],io_md_2[120:94],io_md_2[59:52],
            io_md_2[51:32],io_md_3[120:94],io_md_3[59:52],io_md_3[51:32],io_mdReady); // @[src/main/scala/utils/Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & ~reset) begin
          $fwrite(32'h80000002,"[%d] EmbeddedTLBExec_1: ",c_9); // @[src/main/scala/utils/Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_25) begin
          $fwrite(32'h80000002,
            "md: wen:%d windex:%x waymask:%x vpn:%x asid:%x mask:%x flag:%x asid:%x ppn:%x pteaddr:%x\n",io_mdWrite_wen,
            io_mdWrite_windex,io_mdWrite_waymask,io_mdWrite_wdata[120:94],io_mdWrite_wdata[93:78],io_mdWrite_wdata[77:60
            ],io_mdWrite_wdata[59:52],io_mdWrite_wdata[93:78],io_mdWrite_wdata[51:32],io_mdWrite_wdata[31:0]); // @[src/main/scala/utils/Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & ~reset) begin
          $fwrite(32'h80000002,"[%d] EmbeddedTLBExec_1: ",c_10); // @[src/main/scala/utils/Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_25) begin
          $fwrite(32'h80000002,"MemReq(%d, %d) MemResp(%d, %d) addr:%x cmd:%d rdata:%x cmd:%d\n",io_mem_req_valid,
            io_mem_req_ready,io_mem_resp_valid,io_mem_resp_ready,io_mem_req_bits_addr,io_mem_req_bits_cmd,
            io_mem_resp_bits_rdata,io_mem_resp_bits_cmd); // @[src/main/scala/utils/Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & ~reset) begin
          $fwrite(32'h80000002,"[%d] EmbeddedTLBExec_1: ",c_11); // @[src/main/scala/utils/Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_25) begin
          $fwrite(32'h80000002,"io.ipf:%d hitinstrPF:%d missIPF:%d pf.loadPF:%d pf.storePF:%d loadPF:%d storePF:%d\n",
            io_ipf,1'h0,1'h0,io_pf_loadPF,io_pf_storePF,loadPF,storePF); // @[src/main/scala/utils/Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  victimWaymask_lfsr = _RAND_0[63:0];
  _RAND_1 = {1{`RANDOM}};
  state = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  level = _RAND_2[1:0];
  _RAND_3 = {2{`RANDOM}};
  hitWBStore = _RAND_3[39:0];
  _RAND_4 = {1{`RANDOM}};
  io_pf_loadPF_REG = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  io_pf_storePF_REG = _RAND_5[0:0];
  _RAND_6 = {2{`RANDOM}};
  memRespStore = _RAND_6[63:0];
  _RAND_7 = {1{`RANDOM}};
  missMaskStore = _RAND_7[17:0];
  _RAND_8 = {1{`RANDOM}};
  raddr = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  alreadyOutFire = _RAND_9[0:0];
  _RAND_10 = {2{`RANDOM}};
  c = _RAND_10[63:0];
  _RAND_11 = {1{`RANDOM}};
  REG = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  REG_1 = _RAND_12[3:0];
  _RAND_13 = {1{`RANDOM}};
  REG_2 = _RAND_13[3:0];
  _RAND_14 = {1{`RANDOM}};
  REG_3 = _RAND_14[26:0];
  _RAND_15 = {1{`RANDOM}};
  REG_4 = _RAND_15[15:0];
  _RAND_16 = {1{`RANDOM}};
  REG_5 = _RAND_16[17:0];
  _RAND_17 = {1{`RANDOM}};
  REG_6 = _RAND_17[7:0];
  _RAND_18 = {1{`RANDOM}};
  REG_7 = _RAND_18[19:0];
  _RAND_19 = {1{`RANDOM}};
  REG_8 = _RAND_19[31:0];
  _RAND_20 = {2{`RANDOM}};
  c_4 = _RAND_20[63:0];
  _RAND_21 = {2{`RANDOM}};
  c_5 = _RAND_21[63:0];
  _RAND_22 = {2{`RANDOM}};
  c_6 = _RAND_22[63:0];
  _RAND_23 = {2{`RANDOM}};
  c_7 = _RAND_23[63:0];
  _RAND_24 = {2{`RANDOM}};
  c_8 = _RAND_24[63:0];
  _RAND_25 = {2{`RANDOM}};
  c_9 = _RAND_25[63:0];
  _RAND_26 = {2{`RANDOM}};
  c_10 = _RAND_26[63:0];
  _RAND_27 = {2{`RANDOM}};
  c_11 = _RAND_27[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module EmbeddedTLBEmpty_1(
  output        io_in_ready, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 405:14]
  input         io_in_valid, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 405:14]
  input  [31:0] io_in_bits_addr, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 405:14]
  input  [2:0]  io_in_bits_size, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 405:14]
  input  [3:0]  io_in_bits_cmd, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 405:14]
  input  [7:0]  io_in_bits_wmask, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 405:14]
  input  [63:0] io_in_bits_wdata, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 405:14]
  input         io_out_ready, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 405:14]
  output        io_out_valid, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 405:14]
  output [31:0] io_out_bits_addr, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 405:14]
  output [2:0]  io_out_bits_size, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 405:14]
  output [3:0]  io_out_bits_cmd, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 405:14]
  output [7:0]  io_out_bits_wmask, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 405:14]
  output [63:0] io_out_bits_wdata // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 405:14]
);
  assign io_in_ready = io_out_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 410:10]
  assign io_out_valid = io_in_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 410:10]
  assign io_out_bits_addr = io_in_bits_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 410:10]
  assign io_out_bits_size = io_in_bits_size; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 410:10]
  assign io_out_bits_cmd = io_in_bits_cmd; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 410:10]
  assign io_out_bits_wmask = io_in_bits_wmask; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 410:10]
  assign io_out_bits_wdata = io_in_bits_wdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 410:10]
endmodule
module EmbeddedTLBMD_1(
  input          clock,
  input          reset,
  output [120:0] io_tlbmd_0, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 41:14]
  output [120:0] io_tlbmd_1, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 41:14]
  output [120:0] io_tlbmd_2, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 41:14]
  output [120:0] io_tlbmd_3, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 41:14]
  input          io_write_wen, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 41:14]
  input  [3:0]   io_write_windex, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 41:14]
  input  [3:0]   io_write_waymask, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 41:14]
  input  [120:0] io_write_wdata, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 41:14]
  input  [3:0]   io_rindex, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 41:14]
  output         io_ready // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 41:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [127:0] _RAND_0;
  reg [127:0] _RAND_1;
  reg [127:0] _RAND_2;
  reg [127:0] _RAND_3;
  reg [127:0] _RAND_4;
  reg [127:0] _RAND_5;
  reg [127:0] _RAND_6;
  reg [127:0] _RAND_7;
  reg [127:0] _RAND_8;
  reg [127:0] _RAND_9;
  reg [127:0] _RAND_10;
  reg [127:0] _RAND_11;
  reg [127:0] _RAND_12;
  reg [127:0] _RAND_13;
  reg [127:0] _RAND_14;
  reg [127:0] _RAND_15;
  reg [127:0] _RAND_16;
  reg [127:0] _RAND_17;
  reg [127:0] _RAND_18;
  reg [127:0] _RAND_19;
  reg [127:0] _RAND_20;
  reg [127:0] _RAND_21;
  reg [127:0] _RAND_22;
  reg [127:0] _RAND_23;
  reg [127:0] _RAND_24;
  reg [127:0] _RAND_25;
  reg [127:0] _RAND_26;
  reg [127:0] _RAND_27;
  reg [127:0] _RAND_28;
  reg [127:0] _RAND_29;
  reg [127:0] _RAND_30;
  reg [127:0] _RAND_31;
  reg [127:0] _RAND_32;
  reg [127:0] _RAND_33;
  reg [127:0] _RAND_34;
  reg [127:0] _RAND_35;
  reg [127:0] _RAND_36;
  reg [127:0] _RAND_37;
  reg [127:0] _RAND_38;
  reg [127:0] _RAND_39;
  reg [127:0] _RAND_40;
  reg [127:0] _RAND_41;
  reg [127:0] _RAND_42;
  reg [127:0] _RAND_43;
  reg [127:0] _RAND_44;
  reg [127:0] _RAND_45;
  reg [127:0] _RAND_46;
  reg [127:0] _RAND_47;
  reg [127:0] _RAND_48;
  reg [127:0] _RAND_49;
  reg [127:0] _RAND_50;
  reg [127:0] _RAND_51;
  reg [127:0] _RAND_52;
  reg [127:0] _RAND_53;
  reg [127:0] _RAND_54;
  reg [127:0] _RAND_55;
  reg [127:0] _RAND_56;
  reg [127:0] _RAND_57;
  reg [127:0] _RAND_58;
  reg [127:0] _RAND_59;
  reg [127:0] _RAND_60;
  reg [127:0] _RAND_61;
  reg [127:0] _RAND_62;
  reg [127:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
`endif // RANDOMIZE_REG_INIT
  reg [120:0] tlbmd_0_0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 49:18]
  reg [120:0] tlbmd_0_1; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 49:18]
  reg [120:0] tlbmd_0_2; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 49:18]
  reg [120:0] tlbmd_0_3; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 49:18]
  reg [120:0] tlbmd_1_0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 49:18]
  reg [120:0] tlbmd_1_1; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 49:18]
  reg [120:0] tlbmd_1_2; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 49:18]
  reg [120:0] tlbmd_1_3; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 49:18]
  reg [120:0] tlbmd_2_0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 49:18]
  reg [120:0] tlbmd_2_1; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 49:18]
  reg [120:0] tlbmd_2_2; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 49:18]
  reg [120:0] tlbmd_2_3; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 49:18]
  reg [120:0] tlbmd_3_0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 49:18]
  reg [120:0] tlbmd_3_1; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 49:18]
  reg [120:0] tlbmd_3_2; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 49:18]
  reg [120:0] tlbmd_3_3; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 49:18]
  reg [120:0] tlbmd_4_0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 49:18]
  reg [120:0] tlbmd_4_1; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 49:18]
  reg [120:0] tlbmd_4_2; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 49:18]
  reg [120:0] tlbmd_4_3; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 49:18]
  reg [120:0] tlbmd_5_0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 49:18]
  reg [120:0] tlbmd_5_1; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 49:18]
  reg [120:0] tlbmd_5_2; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 49:18]
  reg [120:0] tlbmd_5_3; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 49:18]
  reg [120:0] tlbmd_6_0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 49:18]
  reg [120:0] tlbmd_6_1; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 49:18]
  reg [120:0] tlbmd_6_2; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 49:18]
  reg [120:0] tlbmd_6_3; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 49:18]
  reg [120:0] tlbmd_7_0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 49:18]
  reg [120:0] tlbmd_7_1; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 49:18]
  reg [120:0] tlbmd_7_2; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 49:18]
  reg [120:0] tlbmd_7_3; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 49:18]
  reg [120:0] tlbmd_8_0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 49:18]
  reg [120:0] tlbmd_8_1; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 49:18]
  reg [120:0] tlbmd_8_2; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 49:18]
  reg [120:0] tlbmd_8_3; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 49:18]
  reg [120:0] tlbmd_9_0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 49:18]
  reg [120:0] tlbmd_9_1; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 49:18]
  reg [120:0] tlbmd_9_2; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 49:18]
  reg [120:0] tlbmd_9_3; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 49:18]
  reg [120:0] tlbmd_10_0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 49:18]
  reg [120:0] tlbmd_10_1; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 49:18]
  reg [120:0] tlbmd_10_2; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 49:18]
  reg [120:0] tlbmd_10_3; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 49:18]
  reg [120:0] tlbmd_11_0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 49:18]
  reg [120:0] tlbmd_11_1; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 49:18]
  reg [120:0] tlbmd_11_2; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 49:18]
  reg [120:0] tlbmd_11_3; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 49:18]
  reg [120:0] tlbmd_12_0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 49:18]
  reg [120:0] tlbmd_12_1; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 49:18]
  reg [120:0] tlbmd_12_2; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 49:18]
  reg [120:0] tlbmd_12_3; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 49:18]
  reg [120:0] tlbmd_13_0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 49:18]
  reg [120:0] tlbmd_13_1; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 49:18]
  reg [120:0] tlbmd_13_2; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 49:18]
  reg [120:0] tlbmd_13_3; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 49:18]
  reg [120:0] tlbmd_14_0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 49:18]
  reg [120:0] tlbmd_14_1; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 49:18]
  reg [120:0] tlbmd_14_2; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 49:18]
  reg [120:0] tlbmd_14_3; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 49:18]
  reg [120:0] tlbmd_15_0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 49:18]
  reg [120:0] tlbmd_15_1; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 49:18]
  reg [120:0] tlbmd_15_2; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 49:18]
  reg [120:0] tlbmd_15_3; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 49:18]
  wire [120:0] _GEN_1 = 4'h1 == io_rindex ? tlbmd_1_0 : tlbmd_0_0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 50:{12,12}]
  wire [120:0] _GEN_2 = 4'h2 == io_rindex ? tlbmd_2_0 : _GEN_1; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 50:{12,12}]
  wire [120:0] _GEN_3 = 4'h3 == io_rindex ? tlbmd_3_0 : _GEN_2; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 50:{12,12}]
  wire [120:0] _GEN_4 = 4'h4 == io_rindex ? tlbmd_4_0 : _GEN_3; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 50:{12,12}]
  wire [120:0] _GEN_5 = 4'h5 == io_rindex ? tlbmd_5_0 : _GEN_4; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 50:{12,12}]
  wire [120:0] _GEN_6 = 4'h6 == io_rindex ? tlbmd_6_0 : _GEN_5; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 50:{12,12}]
  wire [120:0] _GEN_7 = 4'h7 == io_rindex ? tlbmd_7_0 : _GEN_6; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 50:{12,12}]
  wire [120:0] _GEN_8 = 4'h8 == io_rindex ? tlbmd_8_0 : _GEN_7; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 50:{12,12}]
  wire [120:0] _GEN_9 = 4'h9 == io_rindex ? tlbmd_9_0 : _GEN_8; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 50:{12,12}]
  wire [120:0] _GEN_10 = 4'ha == io_rindex ? tlbmd_10_0 : _GEN_9; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 50:{12,12}]
  wire [120:0] _GEN_11 = 4'hb == io_rindex ? tlbmd_11_0 : _GEN_10; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 50:{12,12}]
  wire [120:0] _GEN_12 = 4'hc == io_rindex ? tlbmd_12_0 : _GEN_11; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 50:{12,12}]
  wire [120:0] _GEN_13 = 4'hd == io_rindex ? tlbmd_13_0 : _GEN_12; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 50:{12,12}]
  wire [120:0] _GEN_14 = 4'he == io_rindex ? tlbmd_14_0 : _GEN_13; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 50:{12,12}]
  wire [120:0] _GEN_17 = 4'h1 == io_rindex ? tlbmd_1_1 : tlbmd_0_1; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 50:{12,12}]
  wire [120:0] _GEN_18 = 4'h2 == io_rindex ? tlbmd_2_1 : _GEN_17; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 50:{12,12}]
  wire [120:0] _GEN_19 = 4'h3 == io_rindex ? tlbmd_3_1 : _GEN_18; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 50:{12,12}]
  wire [120:0] _GEN_20 = 4'h4 == io_rindex ? tlbmd_4_1 : _GEN_19; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 50:{12,12}]
  wire [120:0] _GEN_21 = 4'h5 == io_rindex ? tlbmd_5_1 : _GEN_20; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 50:{12,12}]
  wire [120:0] _GEN_22 = 4'h6 == io_rindex ? tlbmd_6_1 : _GEN_21; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 50:{12,12}]
  wire [120:0] _GEN_23 = 4'h7 == io_rindex ? tlbmd_7_1 : _GEN_22; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 50:{12,12}]
  wire [120:0] _GEN_24 = 4'h8 == io_rindex ? tlbmd_8_1 : _GEN_23; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 50:{12,12}]
  wire [120:0] _GEN_25 = 4'h9 == io_rindex ? tlbmd_9_1 : _GEN_24; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 50:{12,12}]
  wire [120:0] _GEN_26 = 4'ha == io_rindex ? tlbmd_10_1 : _GEN_25; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 50:{12,12}]
  wire [120:0] _GEN_27 = 4'hb == io_rindex ? tlbmd_11_1 : _GEN_26; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 50:{12,12}]
  wire [120:0] _GEN_28 = 4'hc == io_rindex ? tlbmd_12_1 : _GEN_27; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 50:{12,12}]
  wire [120:0] _GEN_29 = 4'hd == io_rindex ? tlbmd_13_1 : _GEN_28; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 50:{12,12}]
  wire [120:0] _GEN_30 = 4'he == io_rindex ? tlbmd_14_1 : _GEN_29; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 50:{12,12}]
  wire [120:0] _GEN_33 = 4'h1 == io_rindex ? tlbmd_1_2 : tlbmd_0_2; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 50:{12,12}]
  wire [120:0] _GEN_34 = 4'h2 == io_rindex ? tlbmd_2_2 : _GEN_33; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 50:{12,12}]
  wire [120:0] _GEN_35 = 4'h3 == io_rindex ? tlbmd_3_2 : _GEN_34; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 50:{12,12}]
  wire [120:0] _GEN_36 = 4'h4 == io_rindex ? tlbmd_4_2 : _GEN_35; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 50:{12,12}]
  wire [120:0] _GEN_37 = 4'h5 == io_rindex ? tlbmd_5_2 : _GEN_36; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 50:{12,12}]
  wire [120:0] _GEN_38 = 4'h6 == io_rindex ? tlbmd_6_2 : _GEN_37; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 50:{12,12}]
  wire [120:0] _GEN_39 = 4'h7 == io_rindex ? tlbmd_7_2 : _GEN_38; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 50:{12,12}]
  wire [120:0] _GEN_40 = 4'h8 == io_rindex ? tlbmd_8_2 : _GEN_39; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 50:{12,12}]
  wire [120:0] _GEN_41 = 4'h9 == io_rindex ? tlbmd_9_2 : _GEN_40; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 50:{12,12}]
  wire [120:0] _GEN_42 = 4'ha == io_rindex ? tlbmd_10_2 : _GEN_41; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 50:{12,12}]
  wire [120:0] _GEN_43 = 4'hb == io_rindex ? tlbmd_11_2 : _GEN_42; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 50:{12,12}]
  wire [120:0] _GEN_44 = 4'hc == io_rindex ? tlbmd_12_2 : _GEN_43; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 50:{12,12}]
  wire [120:0] _GEN_45 = 4'hd == io_rindex ? tlbmd_13_2 : _GEN_44; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 50:{12,12}]
  wire [120:0] _GEN_46 = 4'he == io_rindex ? tlbmd_14_2 : _GEN_45; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 50:{12,12}]
  wire [120:0] _GEN_49 = 4'h1 == io_rindex ? tlbmd_1_3 : tlbmd_0_3; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 50:{12,12}]
  wire [120:0] _GEN_50 = 4'h2 == io_rindex ? tlbmd_2_3 : _GEN_49; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 50:{12,12}]
  wire [120:0] _GEN_51 = 4'h3 == io_rindex ? tlbmd_3_3 : _GEN_50; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 50:{12,12}]
  wire [120:0] _GEN_52 = 4'h4 == io_rindex ? tlbmd_4_3 : _GEN_51; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 50:{12,12}]
  wire [120:0] _GEN_53 = 4'h5 == io_rindex ? tlbmd_5_3 : _GEN_52; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 50:{12,12}]
  wire [120:0] _GEN_54 = 4'h6 == io_rindex ? tlbmd_6_3 : _GEN_53; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 50:{12,12}]
  wire [120:0] _GEN_55 = 4'h7 == io_rindex ? tlbmd_7_3 : _GEN_54; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 50:{12,12}]
  wire [120:0] _GEN_56 = 4'h8 == io_rindex ? tlbmd_8_3 : _GEN_55; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 50:{12,12}]
  wire [120:0] _GEN_57 = 4'h9 == io_rindex ? tlbmd_9_3 : _GEN_56; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 50:{12,12}]
  wire [120:0] _GEN_58 = 4'ha == io_rindex ? tlbmd_10_3 : _GEN_57; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 50:{12,12}]
  wire [120:0] _GEN_59 = 4'hb == io_rindex ? tlbmd_11_3 : _GEN_58; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 50:{12,12}]
  wire [120:0] _GEN_60 = 4'hc == io_rindex ? tlbmd_12_3 : _GEN_59; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 50:{12,12}]
  wire [120:0] _GEN_61 = 4'hd == io_rindex ? tlbmd_13_3 : _GEN_60; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 50:{12,12}]
  wire [120:0] _GEN_62 = 4'he == io_rindex ? tlbmd_14_3 : _GEN_61; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 50:{12,12}]
  reg  resetState; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 53:27]
  reg [3:0] resetSet; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
  wire  wrap_wrap = resetSet == 4'hf; // @[src/main/scala/chisel3/util/Counter.scala 73:24]
  wire [3:0] _wrap_value_T_1 = resetSet + 4'h1; // @[src/main/scala/chisel3/util/Counter.scala 77:24]
  wire  resetFinish = resetState & wrap_wrap; // @[src/main/scala/chisel3/util/Counter.scala 118:{16,23} 117:24]
  wire  _GEN_66 = resetFinish ? 1'h0 : resetState; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 55:22 53:27 55:35]
  wire  wen = resetState | io_write_wen; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 62:16]
  wire [3:0] setIdx = resetState ? resetSet : io_write_windex; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 63:19]
  wire [3:0] waymask = resetState ? 4'hf : io_write_waymask; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 64:20]
  assign io_tlbmd_0 = 4'hf == io_rindex ? tlbmd_15_0 : _GEN_14; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 50:{12,12}]
  assign io_tlbmd_1 = 4'hf == io_rindex ? tlbmd_15_1 : _GEN_30; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 50:{12,12}]
  assign io_tlbmd_2 = 4'hf == io_rindex ? tlbmd_15_2 : _GEN_46; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 50:{12,12}]
  assign io_tlbmd_3 = 4'hf == io_rindex ? tlbmd_15_3 : _GEN_62; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 50:{12,12}]
  assign io_ready = ~resetState; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 74:15]
  always @(posedge clock) begin
    if (wen & waymask[0]) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 69:21]
      if (4'h0 == setIdx) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 70:24]
        if (resetState) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 65:21]
          tlbmd_0_0 <= 121'h0;
        end else begin
          tlbmd_0_0 <= io_write_wdata;
        end
      end
    end
    if (wen & waymask[1]) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 69:21]
      if (4'h0 == setIdx) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 70:24]
        if (resetState) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 65:21]
          tlbmd_0_1 <= 121'h0;
        end else begin
          tlbmd_0_1 <= io_write_wdata;
        end
      end
    end
    if (wen & waymask[2]) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 69:21]
      if (4'h0 == setIdx) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 70:24]
        if (resetState) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 65:21]
          tlbmd_0_2 <= 121'h0;
        end else begin
          tlbmd_0_2 <= io_write_wdata;
        end
      end
    end
    if (wen & waymask[3]) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 69:21]
      if (4'h0 == setIdx) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 70:24]
        if (resetState) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 65:21]
          tlbmd_0_3 <= 121'h0;
        end else begin
          tlbmd_0_3 <= io_write_wdata;
        end
      end
    end
    if (wen & waymask[0]) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 69:21]
      if (4'h1 == setIdx) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 70:24]
        if (resetState) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 65:21]
          tlbmd_1_0 <= 121'h0;
        end else begin
          tlbmd_1_0 <= io_write_wdata;
        end
      end
    end
    if (wen & waymask[1]) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 69:21]
      if (4'h1 == setIdx) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 70:24]
        if (resetState) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 65:21]
          tlbmd_1_1 <= 121'h0;
        end else begin
          tlbmd_1_1 <= io_write_wdata;
        end
      end
    end
    if (wen & waymask[2]) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 69:21]
      if (4'h1 == setIdx) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 70:24]
        if (resetState) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 65:21]
          tlbmd_1_2 <= 121'h0;
        end else begin
          tlbmd_1_2 <= io_write_wdata;
        end
      end
    end
    if (wen & waymask[3]) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 69:21]
      if (4'h1 == setIdx) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 70:24]
        if (resetState) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 65:21]
          tlbmd_1_3 <= 121'h0;
        end else begin
          tlbmd_1_3 <= io_write_wdata;
        end
      end
    end
    if (wen & waymask[0]) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 69:21]
      if (4'h2 == setIdx) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 70:24]
        if (resetState) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 65:21]
          tlbmd_2_0 <= 121'h0;
        end else begin
          tlbmd_2_0 <= io_write_wdata;
        end
      end
    end
    if (wen & waymask[1]) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 69:21]
      if (4'h2 == setIdx) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 70:24]
        if (resetState) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 65:21]
          tlbmd_2_1 <= 121'h0;
        end else begin
          tlbmd_2_1 <= io_write_wdata;
        end
      end
    end
    if (wen & waymask[2]) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 69:21]
      if (4'h2 == setIdx) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 70:24]
        if (resetState) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 65:21]
          tlbmd_2_2 <= 121'h0;
        end else begin
          tlbmd_2_2 <= io_write_wdata;
        end
      end
    end
    if (wen & waymask[3]) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 69:21]
      if (4'h2 == setIdx) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 70:24]
        if (resetState) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 65:21]
          tlbmd_2_3 <= 121'h0;
        end else begin
          tlbmd_2_3 <= io_write_wdata;
        end
      end
    end
    if (wen & waymask[0]) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 69:21]
      if (4'h3 == setIdx) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 70:24]
        if (resetState) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 65:21]
          tlbmd_3_0 <= 121'h0;
        end else begin
          tlbmd_3_0 <= io_write_wdata;
        end
      end
    end
    if (wen & waymask[1]) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 69:21]
      if (4'h3 == setIdx) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 70:24]
        if (resetState) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 65:21]
          tlbmd_3_1 <= 121'h0;
        end else begin
          tlbmd_3_1 <= io_write_wdata;
        end
      end
    end
    if (wen & waymask[2]) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 69:21]
      if (4'h3 == setIdx) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 70:24]
        if (resetState) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 65:21]
          tlbmd_3_2 <= 121'h0;
        end else begin
          tlbmd_3_2 <= io_write_wdata;
        end
      end
    end
    if (wen & waymask[3]) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 69:21]
      if (4'h3 == setIdx) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 70:24]
        if (resetState) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 65:21]
          tlbmd_3_3 <= 121'h0;
        end else begin
          tlbmd_3_3 <= io_write_wdata;
        end
      end
    end
    if (wen & waymask[0]) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 69:21]
      if (4'h4 == setIdx) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 70:24]
        if (resetState) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 65:21]
          tlbmd_4_0 <= 121'h0;
        end else begin
          tlbmd_4_0 <= io_write_wdata;
        end
      end
    end
    if (wen & waymask[1]) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 69:21]
      if (4'h4 == setIdx) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 70:24]
        if (resetState) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 65:21]
          tlbmd_4_1 <= 121'h0;
        end else begin
          tlbmd_4_1 <= io_write_wdata;
        end
      end
    end
    if (wen & waymask[2]) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 69:21]
      if (4'h4 == setIdx) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 70:24]
        if (resetState) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 65:21]
          tlbmd_4_2 <= 121'h0;
        end else begin
          tlbmd_4_2 <= io_write_wdata;
        end
      end
    end
    if (wen & waymask[3]) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 69:21]
      if (4'h4 == setIdx) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 70:24]
        if (resetState) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 65:21]
          tlbmd_4_3 <= 121'h0;
        end else begin
          tlbmd_4_3 <= io_write_wdata;
        end
      end
    end
    if (wen & waymask[0]) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 69:21]
      if (4'h5 == setIdx) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 70:24]
        if (resetState) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 65:21]
          tlbmd_5_0 <= 121'h0;
        end else begin
          tlbmd_5_0 <= io_write_wdata;
        end
      end
    end
    if (wen & waymask[1]) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 69:21]
      if (4'h5 == setIdx) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 70:24]
        if (resetState) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 65:21]
          tlbmd_5_1 <= 121'h0;
        end else begin
          tlbmd_5_1 <= io_write_wdata;
        end
      end
    end
    if (wen & waymask[2]) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 69:21]
      if (4'h5 == setIdx) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 70:24]
        if (resetState) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 65:21]
          tlbmd_5_2 <= 121'h0;
        end else begin
          tlbmd_5_2 <= io_write_wdata;
        end
      end
    end
    if (wen & waymask[3]) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 69:21]
      if (4'h5 == setIdx) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 70:24]
        if (resetState) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 65:21]
          tlbmd_5_3 <= 121'h0;
        end else begin
          tlbmd_5_3 <= io_write_wdata;
        end
      end
    end
    if (wen & waymask[0]) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 69:21]
      if (4'h6 == setIdx) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 70:24]
        if (resetState) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 65:21]
          tlbmd_6_0 <= 121'h0;
        end else begin
          tlbmd_6_0 <= io_write_wdata;
        end
      end
    end
    if (wen & waymask[1]) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 69:21]
      if (4'h6 == setIdx) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 70:24]
        if (resetState) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 65:21]
          tlbmd_6_1 <= 121'h0;
        end else begin
          tlbmd_6_1 <= io_write_wdata;
        end
      end
    end
    if (wen & waymask[2]) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 69:21]
      if (4'h6 == setIdx) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 70:24]
        if (resetState) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 65:21]
          tlbmd_6_2 <= 121'h0;
        end else begin
          tlbmd_6_2 <= io_write_wdata;
        end
      end
    end
    if (wen & waymask[3]) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 69:21]
      if (4'h6 == setIdx) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 70:24]
        if (resetState) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 65:21]
          tlbmd_6_3 <= 121'h0;
        end else begin
          tlbmd_6_3 <= io_write_wdata;
        end
      end
    end
    if (wen & waymask[0]) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 69:21]
      if (4'h7 == setIdx) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 70:24]
        if (resetState) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 65:21]
          tlbmd_7_0 <= 121'h0;
        end else begin
          tlbmd_7_0 <= io_write_wdata;
        end
      end
    end
    if (wen & waymask[1]) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 69:21]
      if (4'h7 == setIdx) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 70:24]
        if (resetState) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 65:21]
          tlbmd_7_1 <= 121'h0;
        end else begin
          tlbmd_7_1 <= io_write_wdata;
        end
      end
    end
    if (wen & waymask[2]) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 69:21]
      if (4'h7 == setIdx) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 70:24]
        if (resetState) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 65:21]
          tlbmd_7_2 <= 121'h0;
        end else begin
          tlbmd_7_2 <= io_write_wdata;
        end
      end
    end
    if (wen & waymask[3]) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 69:21]
      if (4'h7 == setIdx) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 70:24]
        if (resetState) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 65:21]
          tlbmd_7_3 <= 121'h0;
        end else begin
          tlbmd_7_3 <= io_write_wdata;
        end
      end
    end
    if (wen & waymask[0]) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 69:21]
      if (4'h8 == setIdx) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 70:24]
        if (resetState) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 65:21]
          tlbmd_8_0 <= 121'h0;
        end else begin
          tlbmd_8_0 <= io_write_wdata;
        end
      end
    end
    if (wen & waymask[1]) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 69:21]
      if (4'h8 == setIdx) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 70:24]
        if (resetState) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 65:21]
          tlbmd_8_1 <= 121'h0;
        end else begin
          tlbmd_8_1 <= io_write_wdata;
        end
      end
    end
    if (wen & waymask[2]) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 69:21]
      if (4'h8 == setIdx) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 70:24]
        if (resetState) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 65:21]
          tlbmd_8_2 <= 121'h0;
        end else begin
          tlbmd_8_2 <= io_write_wdata;
        end
      end
    end
    if (wen & waymask[3]) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 69:21]
      if (4'h8 == setIdx) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 70:24]
        if (resetState) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 65:21]
          tlbmd_8_3 <= 121'h0;
        end else begin
          tlbmd_8_3 <= io_write_wdata;
        end
      end
    end
    if (wen & waymask[0]) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 69:21]
      if (4'h9 == setIdx) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 70:24]
        if (resetState) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 65:21]
          tlbmd_9_0 <= 121'h0;
        end else begin
          tlbmd_9_0 <= io_write_wdata;
        end
      end
    end
    if (wen & waymask[1]) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 69:21]
      if (4'h9 == setIdx) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 70:24]
        if (resetState) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 65:21]
          tlbmd_9_1 <= 121'h0;
        end else begin
          tlbmd_9_1 <= io_write_wdata;
        end
      end
    end
    if (wen & waymask[2]) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 69:21]
      if (4'h9 == setIdx) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 70:24]
        if (resetState) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 65:21]
          tlbmd_9_2 <= 121'h0;
        end else begin
          tlbmd_9_2 <= io_write_wdata;
        end
      end
    end
    if (wen & waymask[3]) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 69:21]
      if (4'h9 == setIdx) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 70:24]
        if (resetState) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 65:21]
          tlbmd_9_3 <= 121'h0;
        end else begin
          tlbmd_9_3 <= io_write_wdata;
        end
      end
    end
    if (wen & waymask[0]) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 69:21]
      if (4'ha == setIdx) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 70:24]
        if (resetState) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 65:21]
          tlbmd_10_0 <= 121'h0;
        end else begin
          tlbmd_10_0 <= io_write_wdata;
        end
      end
    end
    if (wen & waymask[1]) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 69:21]
      if (4'ha == setIdx) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 70:24]
        if (resetState) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 65:21]
          tlbmd_10_1 <= 121'h0;
        end else begin
          tlbmd_10_1 <= io_write_wdata;
        end
      end
    end
    if (wen & waymask[2]) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 69:21]
      if (4'ha == setIdx) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 70:24]
        if (resetState) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 65:21]
          tlbmd_10_2 <= 121'h0;
        end else begin
          tlbmd_10_2 <= io_write_wdata;
        end
      end
    end
    if (wen & waymask[3]) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 69:21]
      if (4'ha == setIdx) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 70:24]
        if (resetState) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 65:21]
          tlbmd_10_3 <= 121'h0;
        end else begin
          tlbmd_10_3 <= io_write_wdata;
        end
      end
    end
    if (wen & waymask[0]) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 69:21]
      if (4'hb == setIdx) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 70:24]
        if (resetState) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 65:21]
          tlbmd_11_0 <= 121'h0;
        end else begin
          tlbmd_11_0 <= io_write_wdata;
        end
      end
    end
    if (wen & waymask[1]) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 69:21]
      if (4'hb == setIdx) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 70:24]
        if (resetState) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 65:21]
          tlbmd_11_1 <= 121'h0;
        end else begin
          tlbmd_11_1 <= io_write_wdata;
        end
      end
    end
    if (wen & waymask[2]) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 69:21]
      if (4'hb == setIdx) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 70:24]
        if (resetState) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 65:21]
          tlbmd_11_2 <= 121'h0;
        end else begin
          tlbmd_11_2 <= io_write_wdata;
        end
      end
    end
    if (wen & waymask[3]) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 69:21]
      if (4'hb == setIdx) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 70:24]
        if (resetState) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 65:21]
          tlbmd_11_3 <= 121'h0;
        end else begin
          tlbmd_11_3 <= io_write_wdata;
        end
      end
    end
    if (wen & waymask[0]) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 69:21]
      if (4'hc == setIdx) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 70:24]
        if (resetState) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 65:21]
          tlbmd_12_0 <= 121'h0;
        end else begin
          tlbmd_12_0 <= io_write_wdata;
        end
      end
    end
    if (wen & waymask[1]) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 69:21]
      if (4'hc == setIdx) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 70:24]
        if (resetState) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 65:21]
          tlbmd_12_1 <= 121'h0;
        end else begin
          tlbmd_12_1 <= io_write_wdata;
        end
      end
    end
    if (wen & waymask[2]) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 69:21]
      if (4'hc == setIdx) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 70:24]
        if (resetState) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 65:21]
          tlbmd_12_2 <= 121'h0;
        end else begin
          tlbmd_12_2 <= io_write_wdata;
        end
      end
    end
    if (wen & waymask[3]) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 69:21]
      if (4'hc == setIdx) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 70:24]
        if (resetState) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 65:21]
          tlbmd_12_3 <= 121'h0;
        end else begin
          tlbmd_12_3 <= io_write_wdata;
        end
      end
    end
    if (wen & waymask[0]) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 69:21]
      if (4'hd == setIdx) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 70:24]
        if (resetState) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 65:21]
          tlbmd_13_0 <= 121'h0;
        end else begin
          tlbmd_13_0 <= io_write_wdata;
        end
      end
    end
    if (wen & waymask[1]) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 69:21]
      if (4'hd == setIdx) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 70:24]
        if (resetState) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 65:21]
          tlbmd_13_1 <= 121'h0;
        end else begin
          tlbmd_13_1 <= io_write_wdata;
        end
      end
    end
    if (wen & waymask[2]) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 69:21]
      if (4'hd == setIdx) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 70:24]
        if (resetState) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 65:21]
          tlbmd_13_2 <= 121'h0;
        end else begin
          tlbmd_13_2 <= io_write_wdata;
        end
      end
    end
    if (wen & waymask[3]) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 69:21]
      if (4'hd == setIdx) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 70:24]
        if (resetState) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 65:21]
          tlbmd_13_3 <= 121'h0;
        end else begin
          tlbmd_13_3 <= io_write_wdata;
        end
      end
    end
    if (wen & waymask[0]) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 69:21]
      if (4'he == setIdx) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 70:24]
        if (resetState) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 65:21]
          tlbmd_14_0 <= 121'h0;
        end else begin
          tlbmd_14_0 <= io_write_wdata;
        end
      end
    end
    if (wen & waymask[1]) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 69:21]
      if (4'he == setIdx) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 70:24]
        if (resetState) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 65:21]
          tlbmd_14_1 <= 121'h0;
        end else begin
          tlbmd_14_1 <= io_write_wdata;
        end
      end
    end
    if (wen & waymask[2]) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 69:21]
      if (4'he == setIdx) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 70:24]
        if (resetState) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 65:21]
          tlbmd_14_2 <= 121'h0;
        end else begin
          tlbmd_14_2 <= io_write_wdata;
        end
      end
    end
    if (wen & waymask[3]) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 69:21]
      if (4'he == setIdx) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 70:24]
        if (resetState) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 65:21]
          tlbmd_14_3 <= 121'h0;
        end else begin
          tlbmd_14_3 <= io_write_wdata;
        end
      end
    end
    if (wen & waymask[0]) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 69:21]
      if (4'hf == setIdx) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 70:24]
        if (resetState) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 65:21]
          tlbmd_15_0 <= 121'h0;
        end else begin
          tlbmd_15_0 <= io_write_wdata;
        end
      end
    end
    if (wen & waymask[1]) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 69:21]
      if (4'hf == setIdx) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 70:24]
        if (resetState) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 65:21]
          tlbmd_15_1 <= 121'h0;
        end else begin
          tlbmd_15_1 <= io_write_wdata;
        end
      end
    end
    if (wen & waymask[2]) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 69:21]
      if (4'hf == setIdx) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 70:24]
        if (resetState) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 65:21]
          tlbmd_15_2 <= 121'h0;
        end else begin
          tlbmd_15_2 <= io_write_wdata;
        end
      end
    end
    if (wen & waymask[3]) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 69:21]
      if (4'hf == setIdx) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 70:24]
        if (resetState) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 65:21]
          tlbmd_15_3 <= 121'h0;
        end else begin
          tlbmd_15_3 <= io_write_wdata;
        end
      end
    end
    resetState <= reset | _GEN_66; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 53:{27,27}]
    if (reset) begin // @[src/main/scala/chisel3/util/Counter.scala 61:40]
      resetSet <= 4'h0; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end else if (resetState) begin // @[src/main/scala/chisel3/util/Counter.scala 118:16]
      resetSet <= _wrap_value_T_1; // @[src/main/scala/chisel3/util/Counter.scala 77:15]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {4{`RANDOM}};
  tlbmd_0_0 = _RAND_0[120:0];
  _RAND_1 = {4{`RANDOM}};
  tlbmd_0_1 = _RAND_1[120:0];
  _RAND_2 = {4{`RANDOM}};
  tlbmd_0_2 = _RAND_2[120:0];
  _RAND_3 = {4{`RANDOM}};
  tlbmd_0_3 = _RAND_3[120:0];
  _RAND_4 = {4{`RANDOM}};
  tlbmd_1_0 = _RAND_4[120:0];
  _RAND_5 = {4{`RANDOM}};
  tlbmd_1_1 = _RAND_5[120:0];
  _RAND_6 = {4{`RANDOM}};
  tlbmd_1_2 = _RAND_6[120:0];
  _RAND_7 = {4{`RANDOM}};
  tlbmd_1_3 = _RAND_7[120:0];
  _RAND_8 = {4{`RANDOM}};
  tlbmd_2_0 = _RAND_8[120:0];
  _RAND_9 = {4{`RANDOM}};
  tlbmd_2_1 = _RAND_9[120:0];
  _RAND_10 = {4{`RANDOM}};
  tlbmd_2_2 = _RAND_10[120:0];
  _RAND_11 = {4{`RANDOM}};
  tlbmd_2_3 = _RAND_11[120:0];
  _RAND_12 = {4{`RANDOM}};
  tlbmd_3_0 = _RAND_12[120:0];
  _RAND_13 = {4{`RANDOM}};
  tlbmd_3_1 = _RAND_13[120:0];
  _RAND_14 = {4{`RANDOM}};
  tlbmd_3_2 = _RAND_14[120:0];
  _RAND_15 = {4{`RANDOM}};
  tlbmd_3_3 = _RAND_15[120:0];
  _RAND_16 = {4{`RANDOM}};
  tlbmd_4_0 = _RAND_16[120:0];
  _RAND_17 = {4{`RANDOM}};
  tlbmd_4_1 = _RAND_17[120:0];
  _RAND_18 = {4{`RANDOM}};
  tlbmd_4_2 = _RAND_18[120:0];
  _RAND_19 = {4{`RANDOM}};
  tlbmd_4_3 = _RAND_19[120:0];
  _RAND_20 = {4{`RANDOM}};
  tlbmd_5_0 = _RAND_20[120:0];
  _RAND_21 = {4{`RANDOM}};
  tlbmd_5_1 = _RAND_21[120:0];
  _RAND_22 = {4{`RANDOM}};
  tlbmd_5_2 = _RAND_22[120:0];
  _RAND_23 = {4{`RANDOM}};
  tlbmd_5_3 = _RAND_23[120:0];
  _RAND_24 = {4{`RANDOM}};
  tlbmd_6_0 = _RAND_24[120:0];
  _RAND_25 = {4{`RANDOM}};
  tlbmd_6_1 = _RAND_25[120:0];
  _RAND_26 = {4{`RANDOM}};
  tlbmd_6_2 = _RAND_26[120:0];
  _RAND_27 = {4{`RANDOM}};
  tlbmd_6_3 = _RAND_27[120:0];
  _RAND_28 = {4{`RANDOM}};
  tlbmd_7_0 = _RAND_28[120:0];
  _RAND_29 = {4{`RANDOM}};
  tlbmd_7_1 = _RAND_29[120:0];
  _RAND_30 = {4{`RANDOM}};
  tlbmd_7_2 = _RAND_30[120:0];
  _RAND_31 = {4{`RANDOM}};
  tlbmd_7_3 = _RAND_31[120:0];
  _RAND_32 = {4{`RANDOM}};
  tlbmd_8_0 = _RAND_32[120:0];
  _RAND_33 = {4{`RANDOM}};
  tlbmd_8_1 = _RAND_33[120:0];
  _RAND_34 = {4{`RANDOM}};
  tlbmd_8_2 = _RAND_34[120:0];
  _RAND_35 = {4{`RANDOM}};
  tlbmd_8_3 = _RAND_35[120:0];
  _RAND_36 = {4{`RANDOM}};
  tlbmd_9_0 = _RAND_36[120:0];
  _RAND_37 = {4{`RANDOM}};
  tlbmd_9_1 = _RAND_37[120:0];
  _RAND_38 = {4{`RANDOM}};
  tlbmd_9_2 = _RAND_38[120:0];
  _RAND_39 = {4{`RANDOM}};
  tlbmd_9_3 = _RAND_39[120:0];
  _RAND_40 = {4{`RANDOM}};
  tlbmd_10_0 = _RAND_40[120:0];
  _RAND_41 = {4{`RANDOM}};
  tlbmd_10_1 = _RAND_41[120:0];
  _RAND_42 = {4{`RANDOM}};
  tlbmd_10_2 = _RAND_42[120:0];
  _RAND_43 = {4{`RANDOM}};
  tlbmd_10_3 = _RAND_43[120:0];
  _RAND_44 = {4{`RANDOM}};
  tlbmd_11_0 = _RAND_44[120:0];
  _RAND_45 = {4{`RANDOM}};
  tlbmd_11_1 = _RAND_45[120:0];
  _RAND_46 = {4{`RANDOM}};
  tlbmd_11_2 = _RAND_46[120:0];
  _RAND_47 = {4{`RANDOM}};
  tlbmd_11_3 = _RAND_47[120:0];
  _RAND_48 = {4{`RANDOM}};
  tlbmd_12_0 = _RAND_48[120:0];
  _RAND_49 = {4{`RANDOM}};
  tlbmd_12_1 = _RAND_49[120:0];
  _RAND_50 = {4{`RANDOM}};
  tlbmd_12_2 = _RAND_50[120:0];
  _RAND_51 = {4{`RANDOM}};
  tlbmd_12_3 = _RAND_51[120:0];
  _RAND_52 = {4{`RANDOM}};
  tlbmd_13_0 = _RAND_52[120:0];
  _RAND_53 = {4{`RANDOM}};
  tlbmd_13_1 = _RAND_53[120:0];
  _RAND_54 = {4{`RANDOM}};
  tlbmd_13_2 = _RAND_54[120:0];
  _RAND_55 = {4{`RANDOM}};
  tlbmd_13_3 = _RAND_55[120:0];
  _RAND_56 = {4{`RANDOM}};
  tlbmd_14_0 = _RAND_56[120:0];
  _RAND_57 = {4{`RANDOM}};
  tlbmd_14_1 = _RAND_57[120:0];
  _RAND_58 = {4{`RANDOM}};
  tlbmd_14_2 = _RAND_58[120:0];
  _RAND_59 = {4{`RANDOM}};
  tlbmd_14_3 = _RAND_59[120:0];
  _RAND_60 = {4{`RANDOM}};
  tlbmd_15_0 = _RAND_60[120:0];
  _RAND_61 = {4{`RANDOM}};
  tlbmd_15_1 = _RAND_61[120:0];
  _RAND_62 = {4{`RANDOM}};
  tlbmd_15_2 = _RAND_62[120:0];
  _RAND_63 = {4{`RANDOM}};
  tlbmd_15_3 = _RAND_63[120:0];
  _RAND_64 = {1{`RANDOM}};
  resetState = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  resetSet = _RAND_65[3:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module EmbeddedTLB_1(
  input         clock,
  input         reset,
  output        io_in_req_ready, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 37:14]
  input         io_in_req_valid, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 37:14]
  input  [38:0] io_in_req_bits_addr, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 37:14]
  input  [2:0]  io_in_req_bits_size, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 37:14]
  input  [3:0]  io_in_req_bits_cmd, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 37:14]
  input  [7:0]  io_in_req_bits_wmask, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 37:14]
  input  [63:0] io_in_req_bits_wdata, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 37:14]
  output        io_in_resp_valid, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 37:14]
  output [3:0]  io_in_resp_bits_cmd, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 37:14]
  output [63:0] io_in_resp_bits_rdata, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 37:14]
  input         io_out_req_ready, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 37:14]
  output        io_out_req_valid, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 37:14]
  output [31:0] io_out_req_bits_addr, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 37:14]
  output [2:0]  io_out_req_bits_size, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 37:14]
  output [3:0]  io_out_req_bits_cmd, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 37:14]
  output [7:0]  io_out_req_bits_wmask, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 37:14]
  output [63:0] io_out_req_bits_wdata, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 37:14]
  output        io_out_resp_ready, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 37:14]
  input         io_out_resp_valid, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 37:14]
  input  [3:0]  io_out_resp_bits_cmd, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 37:14]
  input  [63:0] io_out_resp_bits_rdata, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 37:14]
  input         io_mem_req_ready, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 37:14]
  output        io_mem_req_valid, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 37:14]
  output [31:0] io_mem_req_bits_addr, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 37:14]
  output [3:0]  io_mem_req_bits_cmd, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 37:14]
  output [63:0] io_mem_req_bits_wdata, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 37:14]
  input         io_mem_resp_valid, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 37:14]
  input  [3:0]  io_mem_resp_bits_cmd, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 37:14]
  input  [63:0] io_mem_resp_bits_rdata, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 37:14]
  input  [1:0]  io_csrMMU_priviledgeMode, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 37:14]
  input         io_csrMMU_status_sum, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 37:14]
  input         io_csrMMU_status_mxr, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 37:14]
  output        io_csrMMU_loadPF, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 37:14]
  output        io_csrMMU_storePF, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 37:14]
  output [38:0] io_csrMMU_addr, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 37:14]
  input         io_cacheEmpty, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 37:14]
  output        io_ipf, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 37:14]
  input         _WIRE_4,
  input  [63:0] CSRSATP,
  input         DISPLAY_ENABLE,
  output        _WIRE_1_1,
  input         MOUFlushTLB,
  output        _WIRE_2_3,
  output        _WIRE_16
);
`ifdef RANDOMIZE_REG_INIT
  reg [127:0] _RAND_0;
  reg [127:0] _RAND_1;
  reg [127:0] _RAND_2;
  reg [127:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [63:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [63:0] _RAND_17;
  reg [63:0] _RAND_18;
  reg [63:0] _RAND_19;
  reg [63:0] _RAND_20;
`endif // RANDOMIZE_REG_INIT
  wire  tlbExec_clock; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 85:23]
  wire  tlbExec_reset; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 85:23]
  wire  tlbExec_io_in_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 85:23]
  wire  tlbExec_io_in_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 85:23]
  wire [38:0] tlbExec_io_in_bits_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 85:23]
  wire [2:0] tlbExec_io_in_bits_size; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 85:23]
  wire [3:0] tlbExec_io_in_bits_cmd; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 85:23]
  wire [7:0] tlbExec_io_in_bits_wmask; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 85:23]
  wire [63:0] tlbExec_io_in_bits_wdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 85:23]
  wire  tlbExec_io_out_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 85:23]
  wire  tlbExec_io_out_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 85:23]
  wire [31:0] tlbExec_io_out_bits_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 85:23]
  wire [2:0] tlbExec_io_out_bits_size; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 85:23]
  wire [3:0] tlbExec_io_out_bits_cmd; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 85:23]
  wire [7:0] tlbExec_io_out_bits_wmask; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 85:23]
  wire [63:0] tlbExec_io_out_bits_wdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 85:23]
  wire [120:0] tlbExec_io_md_0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 85:23]
  wire [120:0] tlbExec_io_md_1; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 85:23]
  wire [120:0] tlbExec_io_md_2; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 85:23]
  wire [120:0] tlbExec_io_md_3; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 85:23]
  wire  tlbExec_io_mdWrite_wen; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 85:23]
  wire [3:0] tlbExec_io_mdWrite_windex; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 85:23]
  wire [3:0] tlbExec_io_mdWrite_waymask; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 85:23]
  wire [120:0] tlbExec_io_mdWrite_wdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 85:23]
  wire  tlbExec_io_mdReady; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 85:23]
  wire  tlbExec_io_mem_req_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 85:23]
  wire  tlbExec_io_mem_req_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 85:23]
  wire [31:0] tlbExec_io_mem_req_bits_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 85:23]
  wire [2:0] tlbExec_io_mem_req_bits_size; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 85:23]
  wire [3:0] tlbExec_io_mem_req_bits_cmd; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 85:23]
  wire [7:0] tlbExec_io_mem_req_bits_wmask; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 85:23]
  wire [63:0] tlbExec_io_mem_req_bits_wdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 85:23]
  wire  tlbExec_io_mem_resp_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 85:23]
  wire  tlbExec_io_mem_resp_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 85:23]
  wire [3:0] tlbExec_io_mem_resp_bits_cmd; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 85:23]
  wire [63:0] tlbExec_io_mem_resp_bits_rdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 85:23]
  wire [63:0] tlbExec_io_satp; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 85:23]
  wire [1:0] tlbExec_io_pf_priviledgeMode; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 85:23]
  wire  tlbExec_io_pf_status_sum; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 85:23]
  wire  tlbExec_io_pf_status_mxr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 85:23]
  wire  tlbExec_io_pf_loadPF; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 85:23]
  wire  tlbExec_io_pf_storePF; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 85:23]
  wire [38:0] tlbExec_io_pf_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 85:23]
  wire  tlbExec_io_ipf; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 85:23]
  wire  tlbExec_io_isFinish; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 85:23]
  wire  tlbExec_ISAMO; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 85:23]
  wire  tlbExec_DISPLAY_ENABLE; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 85:23]
  wire  tlbEmpty_io_in_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 86:24]
  wire  tlbEmpty_io_in_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 86:24]
  wire [31:0] tlbEmpty_io_in_bits_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 86:24]
  wire [2:0] tlbEmpty_io_in_bits_size; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 86:24]
  wire [3:0] tlbEmpty_io_in_bits_cmd; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 86:24]
  wire [7:0] tlbEmpty_io_in_bits_wmask; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 86:24]
  wire [63:0] tlbEmpty_io_in_bits_wdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 86:24]
  wire  tlbEmpty_io_out_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 86:24]
  wire  tlbEmpty_io_out_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 86:24]
  wire [31:0] tlbEmpty_io_out_bits_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 86:24]
  wire [2:0] tlbEmpty_io_out_bits_size; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 86:24]
  wire [3:0] tlbEmpty_io_out_bits_cmd; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 86:24]
  wire [7:0] tlbEmpty_io_out_bits_wmask; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 86:24]
  wire [63:0] tlbEmpty_io_out_bits_wdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 86:24]
  wire  mdTLB_clock; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 87:21]
  wire  mdTLB_reset; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 87:21]
  wire [120:0] mdTLB_io_tlbmd_0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 87:21]
  wire [120:0] mdTLB_io_tlbmd_1; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 87:21]
  wire [120:0] mdTLB_io_tlbmd_2; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 87:21]
  wire [120:0] mdTLB_io_tlbmd_3; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 87:21]
  wire  mdTLB_io_write_wen; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 87:21]
  wire [3:0] mdTLB_io_write_windex; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 87:21]
  wire [3:0] mdTLB_io_write_waymask; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 87:21]
  wire [120:0] mdTLB_io_write_wdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 87:21]
  wire [3:0] mdTLB_io_rindex; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 87:21]
  wire  mdTLB_io_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 87:21]
  reg [120:0] r_0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 94:29]
  reg [120:0] r_1; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 94:29]
  reg [120:0] r_2; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 94:29]
  reg [120:0] r_3; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 94:29]
  wire  mdUpdate = io_in_req_valid & tlbExec_io_in_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 119:26]
  wire  vmEnable = CSRSATP[63:60] == 4'h8 & io_csrMMU_priviledgeMode < 2'h3; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 107:57]
  reg  valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 110:24]
  wire  _GEN_4 = tlbExec_io_isFinish ? 1'h0 : valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 110:24 111:{25,33}]
  wire  _GEN_5 = mdUpdate & vmEnable | _GEN_4; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 112:{50,58}]
  reg [38:0] tlbExec_io_in_bits_r_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 116:28]
  reg [2:0] tlbExec_io_in_bits_r_size; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 116:28]
  reg [3:0] tlbExec_io_in_bits_r_cmd; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 116:28]
  reg [7:0] tlbExec_io_in_bits_r_wmask; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 116:28]
  reg [63:0] tlbExec_io_in_bits_r_wdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 116:28]
  wire  _T_2 = tlbEmpty_io_out_ready & tlbEmpty_io_out_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  reg  valid_1; // @[src/main/scala/utils/Pipeline.scala 24:24]
  wire  _GEN_12 = _T_2 ? 1'h0 : valid_1; // @[src/main/scala/utils/Pipeline.scala 24:24 25:{25,33}]
  wire  _T_3 = tlbExec_io_out_valid & tlbEmpty_io_in_ready; // @[src/main/scala/utils/Pipeline.scala 26:22]
  wire  _GEN_13 = tlbExec_io_out_valid & tlbEmpty_io_in_ready | _GEN_12; // @[src/main/scala/utils/Pipeline.scala 26:{38,46}]
  reg [31:0] tlbEmpty_io_in_bits_r_addr; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg [2:0] tlbEmpty_io_in_bits_r_size; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg [3:0] tlbEmpty_io_in_bits_r_cmd; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg [7:0] tlbEmpty_io_in_bits_r_wmask; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg [63:0] tlbEmpty_io_in_bits_r_wdata; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg  alreadyOutFinish; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 147:37]
  wire  _GEN_29 = tlbExec_io_out_valid & ~tlbExec_io_out_ready | alreadyOutFinish; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 147:{37,37,37}]
  wire  _T_5 = tlbExec_io_out_ready & tlbExec_io_out_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  wire  _tlbFinish_T_2 = tlbExec_io_pf_loadPF | tlbExec_io_pf_storePF; // @[src/main/scala/nutcore/Bundle.scala 131:23]
  wire  tlbFinish = tlbExec_io_out_valid & ~alreadyOutFinish | _tlbFinish_T_2; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 149:65]
  reg [63:0] c; // @[src/main/scala/utils/GTimer.scala 24:20]
  wire [63:0] _c_T_1 = c + 64'h1; // @[src/main/scala/utils/GTimer.scala 25:12]
  wire  _T_10 = ~reset; // @[src/main/scala/utils/Debug.scala 56:24]
  reg [63:0] c_1; // @[src/main/scala/utils/GTimer.scala 24:20]
  wire [63:0] _c_T_3 = c_1 + 64'h1; // @[src/main/scala/utils/GTimer.scala 25:12]
  reg [63:0] c_2; // @[src/main/scala/utils/GTimer.scala 24:20]
  wire [63:0] _c_T_5 = c_2 + 64'h1; // @[src/main/scala/utils/GTimer.scala 25:12]
  reg [63:0] c_3; // @[src/main/scala/utils/GTimer.scala 24:20]
  wire [63:0] _c_T_7 = c_3 + 64'h1; // @[src/main/scala/utils/GTimer.scala 25:12]
  wire  _WIRE = tlbFinish; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 149:65]
  wire  _WIRE_1 = io_csrMMU_loadPF | io_csrMMU_storePF; // @[src/main/scala/nutcore/Bundle.scala 131:23]
  wire  _WIRE_2 = vmEnable; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 107:57]
  EmbeddedTLBExec_1 tlbExec ( // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 85:23]
    .clock(tlbExec_clock),
    .reset(tlbExec_reset),
    .io_in_ready(tlbExec_io_in_ready),
    .io_in_valid(tlbExec_io_in_valid),
    .io_in_bits_addr(tlbExec_io_in_bits_addr),
    .io_in_bits_size(tlbExec_io_in_bits_size),
    .io_in_bits_cmd(tlbExec_io_in_bits_cmd),
    .io_in_bits_wmask(tlbExec_io_in_bits_wmask),
    .io_in_bits_wdata(tlbExec_io_in_bits_wdata),
    .io_out_ready(tlbExec_io_out_ready),
    .io_out_valid(tlbExec_io_out_valid),
    .io_out_bits_addr(tlbExec_io_out_bits_addr),
    .io_out_bits_size(tlbExec_io_out_bits_size),
    .io_out_bits_cmd(tlbExec_io_out_bits_cmd),
    .io_out_bits_wmask(tlbExec_io_out_bits_wmask),
    .io_out_bits_wdata(tlbExec_io_out_bits_wdata),
    .io_md_0(tlbExec_io_md_0),
    .io_md_1(tlbExec_io_md_1),
    .io_md_2(tlbExec_io_md_2),
    .io_md_3(tlbExec_io_md_3),
    .io_mdWrite_wen(tlbExec_io_mdWrite_wen),
    .io_mdWrite_windex(tlbExec_io_mdWrite_windex),
    .io_mdWrite_waymask(tlbExec_io_mdWrite_waymask),
    .io_mdWrite_wdata(tlbExec_io_mdWrite_wdata),
    .io_mdReady(tlbExec_io_mdReady),
    .io_mem_req_ready(tlbExec_io_mem_req_ready),
    .io_mem_req_valid(tlbExec_io_mem_req_valid),
    .io_mem_req_bits_addr(tlbExec_io_mem_req_bits_addr),
    .io_mem_req_bits_size(tlbExec_io_mem_req_bits_size),
    .io_mem_req_bits_cmd(tlbExec_io_mem_req_bits_cmd),
    .io_mem_req_bits_wmask(tlbExec_io_mem_req_bits_wmask),
    .io_mem_req_bits_wdata(tlbExec_io_mem_req_bits_wdata),
    .io_mem_resp_ready(tlbExec_io_mem_resp_ready),
    .io_mem_resp_valid(tlbExec_io_mem_resp_valid),
    .io_mem_resp_bits_cmd(tlbExec_io_mem_resp_bits_cmd),
    .io_mem_resp_bits_rdata(tlbExec_io_mem_resp_bits_rdata),
    .io_satp(tlbExec_io_satp),
    .io_pf_priviledgeMode(tlbExec_io_pf_priviledgeMode),
    .io_pf_status_sum(tlbExec_io_pf_status_sum),
    .io_pf_status_mxr(tlbExec_io_pf_status_mxr),
    .io_pf_loadPF(tlbExec_io_pf_loadPF),
    .io_pf_storePF(tlbExec_io_pf_storePF),
    .io_pf_addr(tlbExec_io_pf_addr),
    .io_ipf(tlbExec_io_ipf),
    .io_isFinish(tlbExec_io_isFinish),
    .ISAMO(tlbExec_ISAMO),
    .DISPLAY_ENABLE(tlbExec_DISPLAY_ENABLE)
  );
  EmbeddedTLBEmpty_1 tlbEmpty ( // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 86:24]
    .io_in_ready(tlbEmpty_io_in_ready),
    .io_in_valid(tlbEmpty_io_in_valid),
    .io_in_bits_addr(tlbEmpty_io_in_bits_addr),
    .io_in_bits_size(tlbEmpty_io_in_bits_size),
    .io_in_bits_cmd(tlbEmpty_io_in_bits_cmd),
    .io_in_bits_wmask(tlbEmpty_io_in_bits_wmask),
    .io_in_bits_wdata(tlbEmpty_io_in_bits_wdata),
    .io_out_ready(tlbEmpty_io_out_ready),
    .io_out_valid(tlbEmpty_io_out_valid),
    .io_out_bits_addr(tlbEmpty_io_out_bits_addr),
    .io_out_bits_size(tlbEmpty_io_out_bits_size),
    .io_out_bits_cmd(tlbEmpty_io_out_bits_cmd),
    .io_out_bits_wmask(tlbEmpty_io_out_bits_wmask),
    .io_out_bits_wdata(tlbEmpty_io_out_bits_wdata)
  );
  EmbeddedTLBMD_1 mdTLB ( // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 87:21]
    .clock(mdTLB_clock),
    .reset(mdTLB_reset),
    .io_tlbmd_0(mdTLB_io_tlbmd_0),
    .io_tlbmd_1(mdTLB_io_tlbmd_1),
    .io_tlbmd_2(mdTLB_io_tlbmd_2),
    .io_tlbmd_3(mdTLB_io_tlbmd_3),
    .io_write_wen(mdTLB_io_write_wen),
    .io_write_windex(mdTLB_io_write_windex),
    .io_write_waymask(mdTLB_io_write_waymask),
    .io_write_wdata(mdTLB_io_write_wdata),
    .io_rindex(mdTLB_io_rindex),
    .io_ready(mdTLB_io_ready)
  );
  assign io_in_req_ready = ~vmEnable ? io_out_req_ready : tlbExec_io_in_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 115:16 128:19 132:21]
  assign io_in_resp_valid = io_out_resp_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 143:15]
  assign io_in_resp_bits_cmd = io_out_resp_bits_cmd; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 143:15]
  assign io_in_resp_bits_rdata = io_out_resp_bits_rdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 143:15]
  assign io_out_req_valid = ~vmEnable ? io_in_req_valid : tlbEmpty_io_out_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 128:19 131:22 140:41]
  assign io_out_req_bits_addr = ~vmEnable ? io_in_req_bits_addr[31:0] : tlbEmpty_io_out_bits_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 128:19 133:26 140:41]
  assign io_out_req_bits_size = ~vmEnable ? io_in_req_bits_size : tlbEmpty_io_out_bits_size; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 128:19 134:26 140:41]
  assign io_out_req_bits_cmd = ~vmEnable ? io_in_req_bits_cmd : tlbEmpty_io_out_bits_cmd; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 128:19 135:25 140:41]
  assign io_out_req_bits_wmask = ~vmEnable ? io_in_req_bits_wmask : tlbEmpty_io_out_bits_wmask; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 128:19 136:27 140:41]
  assign io_out_req_bits_wdata = ~vmEnable ? io_in_req_bits_wdata : tlbEmpty_io_out_bits_wdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 128:19 137:27 140:41]
  assign io_out_resp_ready = 1'h1; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 143:15]
  assign io_mem_req_valid = tlbExec_io_mem_req_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 92:18]
  assign io_mem_req_bits_addr = tlbExec_io_mem_req_bits_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 92:18]
  assign io_mem_req_bits_cmd = tlbExec_io_mem_req_bits_cmd; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 92:18]
  assign io_mem_req_bits_wdata = tlbExec_io_mem_req_bits_wdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 92:18]
  assign io_csrMMU_loadPF = tlbExec_io_pf_loadPF; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 93:17]
  assign io_csrMMU_storePF = tlbExec_io_pf_storePF; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 93:17]
  assign io_csrMMU_addr = tlbExec_io_pf_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 93:17]
  assign io_ipf = 1'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 99:10]
  assign _WIRE_1_1 = _WIRE_1;
  assign _WIRE_2_3 = _WIRE_2;
  assign _WIRE_16 = _WIRE;
  assign tlbExec_clock = clock;
  assign tlbExec_reset = reset;
  assign tlbExec_io_in_valid = valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 117:17]
  assign tlbExec_io_in_bits_addr = tlbExec_io_in_bits_r_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 116:16]
  assign tlbExec_io_in_bits_size = tlbExec_io_in_bits_r_size; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 116:16]
  assign tlbExec_io_in_bits_cmd = tlbExec_io_in_bits_r_cmd; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 116:16]
  assign tlbExec_io_in_bits_wmask = tlbExec_io_in_bits_r_wmask; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 116:16]
  assign tlbExec_io_in_bits_wdata = tlbExec_io_in_bits_r_wdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 116:16]
  assign tlbExec_io_out_ready = ~vmEnable | tlbEmpty_io_in_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 128:19 129:26 src/main/scala/utils/Pipeline.scala 29:16]
  assign tlbExec_io_md_0 = r_0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 94:17]
  assign tlbExec_io_md_1 = r_1; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 94:17]
  assign tlbExec_io_md_2 = r_2; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 94:17]
  assign tlbExec_io_md_3 = r_3; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 94:17]
  assign tlbExec_io_mdReady = mdTLB_io_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 95:22]
  assign tlbExec_io_mem_req_ready = io_mem_req_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 92:18]
  assign tlbExec_io_mem_resp_valid = io_mem_resp_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 92:18]
  assign tlbExec_io_mem_resp_bits_cmd = io_mem_resp_bits_cmd; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 92:18]
  assign tlbExec_io_mem_resp_bits_rdata = io_mem_resp_bits_rdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 92:18]
  assign tlbExec_io_satp = CSRSATP; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 81:22]
  assign tlbExec_io_pf_priviledgeMode = io_csrMMU_priviledgeMode; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 93:17]
  assign tlbExec_io_pf_status_sum = io_csrMMU_status_sum; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 93:17]
  assign tlbExec_io_pf_status_mxr = io_csrMMU_status_mxr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 93:17]
  assign tlbExec_ISAMO = _WIRE_4;
  assign tlbExec_DISPLAY_ENABLE = DISPLAY_ENABLE;
  assign tlbEmpty_io_in_valid = valid_1; // @[src/main/scala/utils/Pipeline.scala 31:17]
  assign tlbEmpty_io_in_bits_addr = tlbEmpty_io_in_bits_r_addr; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign tlbEmpty_io_in_bits_size = tlbEmpty_io_in_bits_r_size; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign tlbEmpty_io_in_bits_cmd = tlbEmpty_io_in_bits_r_cmd; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign tlbEmpty_io_in_bits_wmask = tlbEmpty_io_in_bits_r_wmask; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign tlbEmpty_io_in_bits_wdata = tlbEmpty_io_in_bits_r_wdata; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign tlbEmpty_io_out_ready = ~vmEnable | io_out_req_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 128:19 130:52 140:41]
  assign mdTLB_clock = clock;
  assign mdTLB_reset = reset | MOUFlushTLB; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 104:31]
  assign mdTLB_io_write_wen = tlbExec_io_mdWrite_wen; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 97:18]
  assign mdTLB_io_write_windex = tlbExec_io_mdWrite_windex; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 97:18]
  assign mdTLB_io_write_waymask = tlbExec_io_mdWrite_waymask; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 97:18]
  assign mdTLB_io_write_wdata = tlbExec_io_mdWrite_wdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 97:18]
  assign mdTLB_io_rindex = io_in_req_bits_addr[15:12]; // @[src/main/scala/nutcore/mem/TLB.scala 200:19]
  always @(posedge clock) begin
    if (mdUpdate) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 94:29]
      r_0 <= mdTLB_io_tlbmd_0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 94:29]
    end
    if (mdUpdate) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 94:29]
      r_1 <= mdTLB_io_tlbmd_1; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 94:29]
    end
    if (mdUpdate) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 94:29]
      r_2 <= mdTLB_io_tlbmd_2; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 94:29]
    end
    if (mdUpdate) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 94:29]
      r_3 <= mdTLB_io_tlbmd_3; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 94:29]
    end
    if (reset) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 110:24]
      valid <= 1'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 110:24]
    end else begin
      valid <= _GEN_5;
    end
    if (mdUpdate) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 116:28]
      tlbExec_io_in_bits_r_addr <= io_in_req_bits_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 116:28]
    end
    if (mdUpdate) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 116:28]
      tlbExec_io_in_bits_r_size <= io_in_req_bits_size; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 116:28]
    end
    if (mdUpdate) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 116:28]
      tlbExec_io_in_bits_r_cmd <= io_in_req_bits_cmd; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 116:28]
    end
    if (mdUpdate) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 116:28]
      tlbExec_io_in_bits_r_wmask <= io_in_req_bits_wmask; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 116:28]
    end
    if (mdUpdate) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 116:28]
      tlbExec_io_in_bits_r_wdata <= io_in_req_bits_wdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 116:28]
    end
    if (reset) begin // @[src/main/scala/utils/Pipeline.scala 24:24]
      valid_1 <= 1'h0; // @[src/main/scala/utils/Pipeline.scala 24:24]
    end else begin
      valid_1 <= _GEN_13;
    end
    if (_T_3) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      tlbEmpty_io_in_bits_r_addr <= tlbExec_io_out_bits_addr; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_3) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      tlbEmpty_io_in_bits_r_size <= tlbExec_io_out_bits_size; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_3) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      tlbEmpty_io_in_bits_r_cmd <= tlbExec_io_out_bits_cmd; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_3) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      tlbEmpty_io_in_bits_r_wmask <= tlbExec_io_out_bits_wmask; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_3) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      tlbEmpty_io_in_bits_r_wdata <= tlbExec_io_out_bits_wdata; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (reset) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 147:37]
      alreadyOutFinish <= 1'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 147:37]
    end else if (alreadyOutFinish & _T_5) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 148:51]
      alreadyOutFinish <= 1'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 148:70]
    end else begin
      alreadyOutFinish <= _GEN_29;
    end
    if (reset) begin // @[src/main/scala/utils/GTimer.scala 24:20]
      c <= 64'h0; // @[src/main/scala/utils/GTimer.scala 24:20]
    end else begin
      c <= _c_T_1; // @[src/main/scala/utils/GTimer.scala 25:7]
    end
    if (reset) begin // @[src/main/scala/utils/GTimer.scala 24:20]
      c_1 <= 64'h0; // @[src/main/scala/utils/GTimer.scala 24:20]
    end else begin
      c_1 <= _c_T_3; // @[src/main/scala/utils/GTimer.scala 25:7]
    end
    if (reset) begin // @[src/main/scala/utils/GTimer.scala 24:20]
      c_2 <= 64'h0; // @[src/main/scala/utils/GTimer.scala 24:20]
    end else begin
      c_2 <= _c_T_5; // @[src/main/scala/utils/GTimer.scala 25:7]
    end
    if (reset) begin // @[src/main/scala/utils/GTimer.scala 24:20]
      c_3 <= 64'h0; // @[src/main/scala/utils/GTimer.scala 24:20]
    end else begin
      c_3 <= _c_T_7; // @[src/main/scala/utils/GTimer.scala 25:7]
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & ~reset) begin
          $fwrite(32'h80000002,"[%d] EmbeddedTLB_1: ",c); // @[src/main/scala/utils/Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_10) begin
          $fwrite(32'h80000002,"InReq(%d, %d) InResp(%d, %d) OutReq(%d, %d) OutResp(%d, %d) vmEnable:%d mode:%d\n",
            io_in_req_valid,io_in_req_ready,io_in_resp_valid,1'h1,io_out_req_valid,io_out_req_ready,io_out_resp_valid,
            io_out_resp_ready,vmEnable,io_csrMMU_priviledgeMode); // @[src/main/scala/utils/Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & ~reset) begin
          $fwrite(32'h80000002,"[%d] EmbeddedTLB_1: ",c_1); // @[src/main/scala/utils/Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_10) begin
          $fwrite(32'h80000002,"InReq: addr:%x cmd:%d wdata:%x OutReq: addr:%x cmd:%x wdata:%x\n",io_in_req_bits_addr,
            io_in_req_bits_cmd,io_in_req_bits_wdata,io_out_req_bits_addr,io_out_req_bits_cmd,io_out_req_bits_wdata); // @[src/main/scala/utils/Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & ~reset) begin
          $fwrite(32'h80000002,"[%d] EmbeddedTLB_1: ",c_2); // @[src/main/scala/utils/Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_10) begin
          $fwrite(32'h80000002,"OutResp: rdata:%x cmd:%x Inresp: rdata:%x cmd:%x\n",io_out_resp_bits_rdata,
            io_out_resp_bits_cmd,io_in_resp_bits_rdata,io_in_resp_bits_cmd); // @[src/main/scala/utils/Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & ~reset) begin
          $fwrite(32'h80000002,"[%d] EmbeddedTLB_1: ",c_3); // @[src/main/scala/utils/Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_10) begin
          $fwrite(32'h80000002,"satp:%x flush:%d cacheEmpty:%d instrPF:%d loadPF:%d storePF:%d \n",CSRSATP,1'h0,
            io_cacheEmpty,io_ipf,io_csrMMU_loadPF,io_csrMMU_storePF); // @[src/main/scala/utils/Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {4{`RANDOM}};
  r_0 = _RAND_0[120:0];
  _RAND_1 = {4{`RANDOM}};
  r_1 = _RAND_1[120:0];
  _RAND_2 = {4{`RANDOM}};
  r_2 = _RAND_2[120:0];
  _RAND_3 = {4{`RANDOM}};
  r_3 = _RAND_3[120:0];
  _RAND_4 = {1{`RANDOM}};
  valid = _RAND_4[0:0];
  _RAND_5 = {2{`RANDOM}};
  tlbExec_io_in_bits_r_addr = _RAND_5[38:0];
  _RAND_6 = {1{`RANDOM}};
  tlbExec_io_in_bits_r_size = _RAND_6[2:0];
  _RAND_7 = {1{`RANDOM}};
  tlbExec_io_in_bits_r_cmd = _RAND_7[3:0];
  _RAND_8 = {1{`RANDOM}};
  tlbExec_io_in_bits_r_wmask = _RAND_8[7:0];
  _RAND_9 = {2{`RANDOM}};
  tlbExec_io_in_bits_r_wdata = _RAND_9[63:0];
  _RAND_10 = {1{`RANDOM}};
  valid_1 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  tlbEmpty_io_in_bits_r_addr = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  tlbEmpty_io_in_bits_r_size = _RAND_12[2:0];
  _RAND_13 = {1{`RANDOM}};
  tlbEmpty_io_in_bits_r_cmd = _RAND_13[3:0];
  _RAND_14 = {1{`RANDOM}};
  tlbEmpty_io_in_bits_r_wmask = _RAND_14[7:0];
  _RAND_15 = {2{`RANDOM}};
  tlbEmpty_io_in_bits_r_wdata = _RAND_15[63:0];
  _RAND_16 = {1{`RANDOM}};
  alreadyOutFinish = _RAND_16[0:0];
  _RAND_17 = {2{`RANDOM}};
  c = _RAND_17[63:0];
  _RAND_18 = {2{`RANDOM}};
  c_1 = _RAND_18[63:0];
  _RAND_19 = {2{`RANDOM}};
  c_2 = _RAND_19[63:0];
  _RAND_20 = {2{`RANDOM}};
  c_3 = _RAND_20[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module CacheStage1_1(
  input         clock,
  input         reset,
  output        io_in_ready, // @[src/main/scala/nutcore/mem/Cache.scala 133:14]
  input         io_in_valid, // @[src/main/scala/nutcore/mem/Cache.scala 133:14]
  input  [31:0] io_in_bits_addr, // @[src/main/scala/nutcore/mem/Cache.scala 133:14]
  input  [2:0]  io_in_bits_size, // @[src/main/scala/nutcore/mem/Cache.scala 133:14]
  input  [3:0]  io_in_bits_cmd, // @[src/main/scala/nutcore/mem/Cache.scala 133:14]
  input  [7:0]  io_in_bits_wmask, // @[src/main/scala/nutcore/mem/Cache.scala 133:14]
  input  [63:0] io_in_bits_wdata, // @[src/main/scala/nutcore/mem/Cache.scala 133:14]
  input         io_out_ready, // @[src/main/scala/nutcore/mem/Cache.scala 133:14]
  output        io_out_valid, // @[src/main/scala/nutcore/mem/Cache.scala 133:14]
  output [31:0] io_out_bits_req_addr, // @[src/main/scala/nutcore/mem/Cache.scala 133:14]
  output [2:0]  io_out_bits_req_size, // @[src/main/scala/nutcore/mem/Cache.scala 133:14]
  output [3:0]  io_out_bits_req_cmd, // @[src/main/scala/nutcore/mem/Cache.scala 133:14]
  output [7:0]  io_out_bits_req_wmask, // @[src/main/scala/nutcore/mem/Cache.scala 133:14]
  output [63:0] io_out_bits_req_wdata, // @[src/main/scala/nutcore/mem/Cache.scala 133:14]
  input         io_metaReadBus_req_ready, // @[src/main/scala/nutcore/mem/Cache.scala 133:14]
  output        io_metaReadBus_req_valid, // @[src/main/scala/nutcore/mem/Cache.scala 133:14]
  output [6:0]  io_metaReadBus_req_bits_setIdx, // @[src/main/scala/nutcore/mem/Cache.scala 133:14]
  input  [18:0] io_metaReadBus_resp_data_0_tag, // @[src/main/scala/nutcore/mem/Cache.scala 133:14]
  input         io_metaReadBus_resp_data_0_valid, // @[src/main/scala/nutcore/mem/Cache.scala 133:14]
  input         io_metaReadBus_resp_data_0_dirty, // @[src/main/scala/nutcore/mem/Cache.scala 133:14]
  input  [18:0] io_metaReadBus_resp_data_1_tag, // @[src/main/scala/nutcore/mem/Cache.scala 133:14]
  input         io_metaReadBus_resp_data_1_valid, // @[src/main/scala/nutcore/mem/Cache.scala 133:14]
  input         io_metaReadBus_resp_data_1_dirty, // @[src/main/scala/nutcore/mem/Cache.scala 133:14]
  input  [18:0] io_metaReadBus_resp_data_2_tag, // @[src/main/scala/nutcore/mem/Cache.scala 133:14]
  input         io_metaReadBus_resp_data_2_valid, // @[src/main/scala/nutcore/mem/Cache.scala 133:14]
  input         io_metaReadBus_resp_data_2_dirty, // @[src/main/scala/nutcore/mem/Cache.scala 133:14]
  input  [18:0] io_metaReadBus_resp_data_3_tag, // @[src/main/scala/nutcore/mem/Cache.scala 133:14]
  input         io_metaReadBus_resp_data_3_valid, // @[src/main/scala/nutcore/mem/Cache.scala 133:14]
  input         io_metaReadBus_resp_data_3_dirty, // @[src/main/scala/nutcore/mem/Cache.scala 133:14]
  input         io_dataReadBus_req_ready, // @[src/main/scala/nutcore/mem/Cache.scala 133:14]
  output        io_dataReadBus_req_valid, // @[src/main/scala/nutcore/mem/Cache.scala 133:14]
  output [9:0]  io_dataReadBus_req_bits_setIdx, // @[src/main/scala/nutcore/mem/Cache.scala 133:14]
  input  [63:0] io_dataReadBus_resp_data_0_data, // @[src/main/scala/nutcore/mem/Cache.scala 133:14]
  input  [63:0] io_dataReadBus_resp_data_1_data, // @[src/main/scala/nutcore/mem/Cache.scala 133:14]
  input  [63:0] io_dataReadBus_resp_data_2_data, // @[src/main/scala/nutcore/mem/Cache.scala 133:14]
  input  [63:0] io_dataReadBus_resp_data_3_data, // @[src/main/scala/nutcore/mem/Cache.scala 133:14]
  input         DISPLAY_ENABLE
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  wire  _T = io_in_ready & io_in_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  reg [63:0] c; // @[src/main/scala/utils/GTimer.scala 24:20]
  wire [63:0] _c_T_1 = c + 64'h1; // @[src/main/scala/utils/GTimer.scala 25:12]
  wire  _T_1 = _T & DISPLAY_ENABLE; // @[src/main/scala/utils/Debug.scala 55:16]
  wire  _T_3 = ~reset; // @[src/main/scala/utils/Debug.scala 56:24]
  wire  _io_in_ready_T_1 = io_out_ready & io_out_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  reg [63:0] c_1; // @[src/main/scala/utils/GTimer.scala 24:20]
  wire [63:0] _c_T_3 = c_1 + 64'h1; // @[src/main/scala/utils/GTimer.scala 25:12]
  assign io_in_ready = (~io_in_valid | _io_in_ready_T_1) & io_metaReadBus_req_ready & io_dataReadBus_req_ready; // @[src/main/scala/nutcore/mem/Cache.scala 145:76]
  assign io_out_valid = io_in_valid & io_metaReadBus_req_ready & io_dataReadBus_req_ready; // @[src/main/scala/nutcore/mem/Cache.scala 144:59]
  assign io_out_bits_req_addr = io_in_bits_addr; // @[src/main/scala/nutcore/mem/Cache.scala 143:19]
  assign io_out_bits_req_size = io_in_bits_size; // @[src/main/scala/nutcore/mem/Cache.scala 143:19]
  assign io_out_bits_req_cmd = io_in_bits_cmd; // @[src/main/scala/nutcore/mem/Cache.scala 143:19]
  assign io_out_bits_req_wmask = io_in_bits_wmask; // @[src/main/scala/nutcore/mem/Cache.scala 143:19]
  assign io_out_bits_req_wdata = io_in_bits_wdata; // @[src/main/scala/nutcore/mem/Cache.scala 143:19]
  assign io_metaReadBus_req_valid = io_in_valid & io_out_ready; // @[src/main/scala/nutcore/mem/Cache.scala 139:34]
  assign io_metaReadBus_req_bits_setIdx = io_in_bits_addr[12:6]; // @[src/main/scala/nutcore/mem/Cache.scala 77:45]
  assign io_dataReadBus_req_valid = io_in_valid & io_out_ready; // @[src/main/scala/nutcore/mem/Cache.scala 139:34]
  assign io_dataReadBus_req_bits_setIdx = {io_in_bits_addr[12:6],io_in_bits_addr[5:3]}; // @[src/main/scala/nutcore/mem/Cache.scala 78:35]
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/utils/GTimer.scala 24:20]
      c <= 64'h0; // @[src/main/scala/utils/GTimer.scala 24:20]
    end else begin
      c <= _c_T_1; // @[src/main/scala/utils/GTimer.scala 25:7]
    end
    if (reset) begin // @[src/main/scala/utils/GTimer.scala 24:20]
      c_1 <= 64'h0; // @[src/main/scala/utils/GTimer.scala 24:20]
    end else begin
      c_1 <= _c_T_3; // @[src/main/scala/utils/GTimer.scala 25:7]
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1 & ~reset) begin
          $fwrite(32'h80000002,"[%d] CacheStage1_1: ",c); // @[src/main/scala/utils/Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1 & _T_3) begin
          $fwrite(32'h80000002,"[L1$] cache stage1, addr in: %x, user: %x id: %x\n",io_in_bits_addr,1'h0,1'h0); // @[src/main/scala/utils/Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & ~reset) begin
          $fwrite(32'h80000002,"[%d] CacheStage1_1: ",c_1); // @[src/main/scala/utils/Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_3) begin
          $fwrite(32'h80000002,
            "in.ready = %d, in.valid = %d, out.valid = %d, out.ready = %d, addr = %x, cmd = %x, dataReadBus.req.valid = %d\n"
            ,io_in_ready,io_in_valid,io_out_valid,io_out_ready,io_in_bits_addr,io_in_bits_cmd,io_dataReadBus_req_valid); // @[src/main/scala/utils/Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  c = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  c_1 = _RAND_1[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module CacheStage2_1(
  input         clock,
  input         reset,
  output        io_in_ready, // @[src/main/scala/nutcore/mem/Cache.scala 171:14]
  input         io_in_valid, // @[src/main/scala/nutcore/mem/Cache.scala 171:14]
  input  [31:0] io_in_bits_req_addr, // @[src/main/scala/nutcore/mem/Cache.scala 171:14]
  input  [2:0]  io_in_bits_req_size, // @[src/main/scala/nutcore/mem/Cache.scala 171:14]
  input  [3:0]  io_in_bits_req_cmd, // @[src/main/scala/nutcore/mem/Cache.scala 171:14]
  input  [7:0]  io_in_bits_req_wmask, // @[src/main/scala/nutcore/mem/Cache.scala 171:14]
  input  [63:0] io_in_bits_req_wdata, // @[src/main/scala/nutcore/mem/Cache.scala 171:14]
  input         io_out_ready, // @[src/main/scala/nutcore/mem/Cache.scala 171:14]
  output        io_out_valid, // @[src/main/scala/nutcore/mem/Cache.scala 171:14]
  output [31:0] io_out_bits_req_addr, // @[src/main/scala/nutcore/mem/Cache.scala 171:14]
  output [2:0]  io_out_bits_req_size, // @[src/main/scala/nutcore/mem/Cache.scala 171:14]
  output [3:0]  io_out_bits_req_cmd, // @[src/main/scala/nutcore/mem/Cache.scala 171:14]
  output [7:0]  io_out_bits_req_wmask, // @[src/main/scala/nutcore/mem/Cache.scala 171:14]
  output [63:0] io_out_bits_req_wdata, // @[src/main/scala/nutcore/mem/Cache.scala 171:14]
  output [18:0] io_out_bits_metas_0_tag, // @[src/main/scala/nutcore/mem/Cache.scala 171:14]
  output        io_out_bits_metas_0_valid, // @[src/main/scala/nutcore/mem/Cache.scala 171:14]
  output        io_out_bits_metas_0_dirty, // @[src/main/scala/nutcore/mem/Cache.scala 171:14]
  output [18:0] io_out_bits_metas_1_tag, // @[src/main/scala/nutcore/mem/Cache.scala 171:14]
  output        io_out_bits_metas_1_valid, // @[src/main/scala/nutcore/mem/Cache.scala 171:14]
  output        io_out_bits_metas_1_dirty, // @[src/main/scala/nutcore/mem/Cache.scala 171:14]
  output [18:0] io_out_bits_metas_2_tag, // @[src/main/scala/nutcore/mem/Cache.scala 171:14]
  output        io_out_bits_metas_2_valid, // @[src/main/scala/nutcore/mem/Cache.scala 171:14]
  output        io_out_bits_metas_2_dirty, // @[src/main/scala/nutcore/mem/Cache.scala 171:14]
  output [18:0] io_out_bits_metas_3_tag, // @[src/main/scala/nutcore/mem/Cache.scala 171:14]
  output        io_out_bits_metas_3_valid, // @[src/main/scala/nutcore/mem/Cache.scala 171:14]
  output        io_out_bits_metas_3_dirty, // @[src/main/scala/nutcore/mem/Cache.scala 171:14]
  output [63:0] io_out_bits_datas_0_data, // @[src/main/scala/nutcore/mem/Cache.scala 171:14]
  output [63:0] io_out_bits_datas_1_data, // @[src/main/scala/nutcore/mem/Cache.scala 171:14]
  output [63:0] io_out_bits_datas_2_data, // @[src/main/scala/nutcore/mem/Cache.scala 171:14]
  output [63:0] io_out_bits_datas_3_data, // @[src/main/scala/nutcore/mem/Cache.scala 171:14]
  output        io_out_bits_hit, // @[src/main/scala/nutcore/mem/Cache.scala 171:14]
  output [3:0]  io_out_bits_waymask, // @[src/main/scala/nutcore/mem/Cache.scala 171:14]
  output        io_out_bits_mmio, // @[src/main/scala/nutcore/mem/Cache.scala 171:14]
  output        io_out_bits_isForwardData, // @[src/main/scala/nutcore/mem/Cache.scala 171:14]
  output [63:0] io_out_bits_forwardData_data_data, // @[src/main/scala/nutcore/mem/Cache.scala 171:14]
  output [3:0]  io_out_bits_forwardData_waymask, // @[src/main/scala/nutcore/mem/Cache.scala 171:14]
  input  [18:0] io_metaReadResp_0_tag, // @[src/main/scala/nutcore/mem/Cache.scala 171:14]
  input         io_metaReadResp_0_valid, // @[src/main/scala/nutcore/mem/Cache.scala 171:14]
  input         io_metaReadResp_0_dirty, // @[src/main/scala/nutcore/mem/Cache.scala 171:14]
  input  [18:0] io_metaReadResp_1_tag, // @[src/main/scala/nutcore/mem/Cache.scala 171:14]
  input         io_metaReadResp_1_valid, // @[src/main/scala/nutcore/mem/Cache.scala 171:14]
  input         io_metaReadResp_1_dirty, // @[src/main/scala/nutcore/mem/Cache.scala 171:14]
  input  [18:0] io_metaReadResp_2_tag, // @[src/main/scala/nutcore/mem/Cache.scala 171:14]
  input         io_metaReadResp_2_valid, // @[src/main/scala/nutcore/mem/Cache.scala 171:14]
  input         io_metaReadResp_2_dirty, // @[src/main/scala/nutcore/mem/Cache.scala 171:14]
  input  [18:0] io_metaReadResp_3_tag, // @[src/main/scala/nutcore/mem/Cache.scala 171:14]
  input         io_metaReadResp_3_valid, // @[src/main/scala/nutcore/mem/Cache.scala 171:14]
  input         io_metaReadResp_3_dirty, // @[src/main/scala/nutcore/mem/Cache.scala 171:14]
  input  [63:0] io_dataReadResp_0_data, // @[src/main/scala/nutcore/mem/Cache.scala 171:14]
  input  [63:0] io_dataReadResp_1_data, // @[src/main/scala/nutcore/mem/Cache.scala 171:14]
  input  [63:0] io_dataReadResp_2_data, // @[src/main/scala/nutcore/mem/Cache.scala 171:14]
  input  [63:0] io_dataReadResp_3_data, // @[src/main/scala/nutcore/mem/Cache.scala 171:14]
  input         io_metaWriteBus_req_valid, // @[src/main/scala/nutcore/mem/Cache.scala 171:14]
  input  [6:0]  io_metaWriteBus_req_bits_setIdx, // @[src/main/scala/nutcore/mem/Cache.scala 171:14]
  input  [18:0] io_metaWriteBus_req_bits_data_tag, // @[src/main/scala/nutcore/mem/Cache.scala 171:14]
  input         io_metaWriteBus_req_bits_data_dirty, // @[src/main/scala/nutcore/mem/Cache.scala 171:14]
  input  [3:0]  io_metaWriteBus_req_bits_waymask, // @[src/main/scala/nutcore/mem/Cache.scala 171:14]
  input         io_dataWriteBus_req_valid, // @[src/main/scala/nutcore/mem/Cache.scala 171:14]
  input  [9:0]  io_dataWriteBus_req_bits_setIdx, // @[src/main/scala/nutcore/mem/Cache.scala 171:14]
  input  [63:0] io_dataWriteBus_req_bits_data_data, // @[src/main/scala/nutcore/mem/Cache.scala 171:14]
  input  [3:0]  io_dataWriteBus_req_bits_waymask, // @[src/main/scala/nutcore/mem/Cache.scala 171:14]
  input         DISPLAY_ENABLE
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [63:0] _RAND_12;
  reg [63:0] _RAND_13;
  reg [63:0] _RAND_14;
  reg [63:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [63:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [63:0] _RAND_19;
  reg [63:0] _RAND_20;
`endif // RANDOMIZE_REG_INIT
  wire [2:0] addr_wordIndex = io_in_bits_req_addr[5:3]; // @[src/main/scala/nutcore/mem/Cache.scala 174:31]
  wire [6:0] addr_index = io_in_bits_req_addr[12:6]; // @[src/main/scala/nutcore/mem/Cache.scala 174:31]
  wire [18:0] addr_tag = io_in_bits_req_addr[31:13]; // @[src/main/scala/nutcore/mem/Cache.scala 174:31]
  wire  isForwardMeta = io_in_valid & io_metaWriteBus_req_valid & io_metaWriteBus_req_bits_setIdx == addr_index; // @[src/main/scala/nutcore/mem/Cache.scala 176:64]
  reg  isForwardMetaReg; // @[src/main/scala/nutcore/mem/Cache.scala 177:33]
  wire  _GEN_0 = isForwardMeta | isForwardMetaReg; // @[src/main/scala/nutcore/mem/Cache.scala 178:24 177:33 178:43]
  wire  _T = io_in_ready & io_in_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  wire  _T_1 = ~io_in_valid; // @[src/main/scala/nutcore/mem/Cache.scala 179:23]
  wire  _T_2 = _T | ~io_in_valid; // @[src/main/scala/nutcore/mem/Cache.scala 179:20]
  reg [18:0] forwardMetaReg_data_tag; // @[src/main/scala/nutcore/mem/Cache.scala 180:33]
  reg  forwardMetaReg_data_dirty; // @[src/main/scala/nutcore/mem/Cache.scala 180:33]
  reg [3:0] forwardMetaReg_waymask; // @[src/main/scala/nutcore/mem/Cache.scala 180:33]
  wire [18:0] _GEN_3 = isForwardMeta ? io_metaWriteBus_req_bits_data_tag : forwardMetaReg_data_tag; // @[src/main/scala/nutcore/mem/Cache.scala 180:{33,33,33}]
  wire  _GEN_5 = isForwardMeta ? io_metaWriteBus_req_bits_data_dirty : forwardMetaReg_data_dirty; // @[src/main/scala/nutcore/mem/Cache.scala 180:{33,33,33}]
  wire [3:0] _GEN_6 = isForwardMeta ? io_metaWriteBus_req_bits_waymask : forwardMetaReg_waymask; // @[src/main/scala/nutcore/mem/Cache.scala 180:{33,33,33}]
  wire  pickForwardMeta = isForwardMetaReg | isForwardMeta; // @[src/main/scala/nutcore/mem/Cache.scala 183:42]
  wire  forwardWaymask_0 = _GEN_6[0]; // @[src/main/scala/nutcore/mem/Cache.scala 185:61]
  wire  forwardWaymask_1 = _GEN_6[1]; // @[src/main/scala/nutcore/mem/Cache.scala 185:61]
  wire  forwardWaymask_2 = _GEN_6[2]; // @[src/main/scala/nutcore/mem/Cache.scala 185:61]
  wire  forwardWaymask_3 = _GEN_6[3]; // @[src/main/scala/nutcore/mem/Cache.scala 185:61]
  wire [18:0] metaWay_0_tag = pickForwardMeta & forwardWaymask_0 ? _GEN_3 : io_metaReadResp_0_tag; // @[src/main/scala/nutcore/mem/Cache.scala 187:22]
  wire  metaWay_0_valid = pickForwardMeta & forwardWaymask_0 | io_metaReadResp_0_valid; // @[src/main/scala/nutcore/mem/Cache.scala 187:22]
  wire [18:0] metaWay_1_tag = pickForwardMeta & forwardWaymask_1 ? _GEN_3 : io_metaReadResp_1_tag; // @[src/main/scala/nutcore/mem/Cache.scala 187:22]
  wire  metaWay_1_valid = pickForwardMeta & forwardWaymask_1 | io_metaReadResp_1_valid; // @[src/main/scala/nutcore/mem/Cache.scala 187:22]
  wire [18:0] metaWay_2_tag = pickForwardMeta & forwardWaymask_2 ? _GEN_3 : io_metaReadResp_2_tag; // @[src/main/scala/nutcore/mem/Cache.scala 187:22]
  wire  metaWay_2_valid = pickForwardMeta & forwardWaymask_2 | io_metaReadResp_2_valid; // @[src/main/scala/nutcore/mem/Cache.scala 187:22]
  wire [18:0] metaWay_3_tag = pickForwardMeta & forwardWaymask_3 ? _GEN_3 : io_metaReadResp_3_tag; // @[src/main/scala/nutcore/mem/Cache.scala 187:22]
  wire  metaWay_3_valid = pickForwardMeta & forwardWaymask_3 | io_metaReadResp_3_valid; // @[src/main/scala/nutcore/mem/Cache.scala 187:22]
  wire  _hitVec_T_2 = metaWay_0_valid & metaWay_0_tag == addr_tag & io_in_valid; // @[src/main/scala/nutcore/mem/Cache.scala 190:73]
  wire  _hitVec_T_5 = metaWay_1_valid & metaWay_1_tag == addr_tag & io_in_valid; // @[src/main/scala/nutcore/mem/Cache.scala 190:73]
  wire  _hitVec_T_8 = metaWay_2_valid & metaWay_2_tag == addr_tag & io_in_valid; // @[src/main/scala/nutcore/mem/Cache.scala 190:73]
  wire  _hitVec_T_11 = metaWay_3_valid & metaWay_3_tag == addr_tag & io_in_valid; // @[src/main/scala/nutcore/mem/Cache.scala 190:73]
  wire [3:0] hitVec = {_hitVec_T_11,_hitVec_T_8,_hitVec_T_5,_hitVec_T_2}; // @[src/main/scala/nutcore/mem/Cache.scala 190:90]
  reg [63:0] victimWaymask_lfsr; // @[src/main/scala/utils/LFSR64.scala 25:23]
  wire  victimWaymask_xor = victimWaymask_lfsr[0] ^ victimWaymask_lfsr[1] ^ victimWaymask_lfsr[3] ^ victimWaymask_lfsr[4
    ]; // @[src/main/scala/utils/LFSR64.scala 26:43]
  wire [63:0] _victimWaymask_lfsr_T_2 = {victimWaymask_xor,victimWaymask_lfsr[63:1]}; // @[src/main/scala/utils/LFSR64.scala 28:41]
  wire [3:0] victimWaymask = 4'h1 << victimWaymask_lfsr[1:0]; // @[src/main/scala/nutcore/mem/Cache.scala 191:42]
  wire  _invalidVec_T = ~metaWay_0_valid; // @[src/main/scala/nutcore/mem/Cache.scala 193:45]
  wire  _invalidVec_T_1 = ~metaWay_1_valid; // @[src/main/scala/nutcore/mem/Cache.scala 193:45]
  wire  _invalidVec_T_2 = ~metaWay_2_valid; // @[src/main/scala/nutcore/mem/Cache.scala 193:45]
  wire  _invalidVec_T_3 = ~metaWay_3_valid; // @[src/main/scala/nutcore/mem/Cache.scala 193:45]
  wire [3:0] invalidVec = {_invalidVec_T_3,_invalidVec_T_2,_invalidVec_T_1,_invalidVec_T}; // @[src/main/scala/nutcore/mem/Cache.scala 193:56]
  wire  hasInvalidWay = |invalidVec; // @[src/main/scala/nutcore/mem/Cache.scala 194:34]
  wire [1:0] _refillInvalidWaymask_T_3 = invalidVec >= 4'h2 ? 2'h2 : 2'h1; // @[src/main/scala/nutcore/mem/Cache.scala 197:8]
  wire [2:0] _refillInvalidWaymask_T_4 = invalidVec >= 4'h4 ? 3'h4 : {{1'd0}, _refillInvalidWaymask_T_3}; // @[src/main/scala/nutcore/mem/Cache.scala 196:8]
  wire [3:0] refillInvalidWaymask = invalidVec >= 4'h8 ? 4'h8 : {{1'd0}, _refillInvalidWaymask_T_4}; // @[src/main/scala/nutcore/mem/Cache.scala 195:33]
  wire [3:0] _waymask_T = hasInvalidWay ? refillInvalidWaymask : victimWaymask; // @[src/main/scala/nutcore/mem/Cache.scala 200:49]
  wire [3:0] waymask = io_out_bits_hit ? hitVec : _waymask_T; // @[src/main/scala/nutcore/mem/Cache.scala 200:20]
  wire [1:0] _T_7 = waymask[0] + waymask[1]; // @[src/main/scala/nutcore/mem/Cache.scala 201:16]
  wire [1:0] _T_9 = waymask[2] + waymask[3]; // @[src/main/scala/nutcore/mem/Cache.scala 201:16]
  wire [2:0] _T_11 = _T_7 + _T_9; // @[src/main/scala/nutcore/mem/Cache.scala 201:16]
  wire  _T_13 = _T_11 > 3'h1; // @[src/main/scala/nutcore/mem/Cache.scala 201:26]
  reg [63:0] c; // @[src/main/scala/utils/GTimer.scala 24:20]
  wire [63:0] _c_T_1 = c + 64'h1; // @[src/main/scala/utils/GTimer.scala 25:12]
  wire  _T_16 = ~reset; // @[src/main/scala/utils/Debug.scala 56:24]
  reg [63:0] c_1; // @[src/main/scala/utils/GTimer.scala 24:20]
  wire [63:0] _c_T_3 = c_1 + 64'h1; // @[src/main/scala/utils/GTimer.scala 25:12]
  reg [63:0] c_2; // @[src/main/scala/utils/GTimer.scala 24:20]
  wire [63:0] _c_T_5 = c_2 + 64'h1; // @[src/main/scala/utils/GTimer.scala 25:12]
  reg [63:0] c_3; // @[src/main/scala/utils/GTimer.scala 24:20]
  wire [63:0] _c_T_7 = c_3 + 64'h1; // @[src/main/scala/utils/GTimer.scala 25:12]
  reg [63:0] c_4; // @[src/main/scala/utils/GTimer.scala 24:20]
  wire [63:0] _c_T_9 = c_4 + 64'h1; // @[src/main/scala/utils/GTimer.scala 25:12]
  reg [63:0] c_5; // @[src/main/scala/utils/GTimer.scala 24:20]
  wire [63:0] _c_T_11 = c_5 + 64'h1; // @[src/main/scala/utils/GTimer.scala 25:12]
  reg [63:0] c_6; // @[src/main/scala/utils/GTimer.scala 24:20]
  wire [63:0] _c_T_13 = c_6 + 64'h1; // @[src/main/scala/utils/GTimer.scala 25:12]
  reg [63:0] c_7; // @[src/main/scala/utils/GTimer.scala 24:20]
  wire [63:0] _c_T_15 = c_7 + 64'h1; // @[src/main/scala/utils/GTimer.scala 25:12]
  reg [63:0] c_8; // @[src/main/scala/utils/GTimer.scala 24:20]
  wire [63:0] _c_T_17 = c_8 + 64'h1; // @[src/main/scala/utils/GTimer.scala 25:12]
  reg [63:0] c_9; // @[src/main/scala/utils/GTimer.scala 24:20]
  wire [63:0] _c_T_19 = c_9 + 64'h1; // @[src/main/scala/utils/GTimer.scala 25:12]
  reg [63:0] c_10; // @[src/main/scala/utils/GTimer.scala 24:20]
  wire [63:0] _c_T_21 = c_10 + 64'h1; // @[src/main/scala/utils/GTimer.scala 25:12]
  wire [31:0] _io_out_bits_mmio_T = io_in_bits_req_addr ^ 32'h30000000; // @[src/main/scala/nutcore/NutCore.scala 87:11]
  wire  _io_out_bits_mmio_T_2 = _io_out_bits_mmio_T[31:28] == 4'h0; // @[src/main/scala/nutcore/NutCore.scala 87:44]
  wire [31:0] _io_out_bits_mmio_T_3 = io_in_bits_req_addr ^ 32'h40000000; // @[src/main/scala/nutcore/NutCore.scala 87:11]
  wire  _io_out_bits_mmio_T_5 = _io_out_bits_mmio_T_3[31:30] == 2'h0; // @[src/main/scala/nutcore/NutCore.scala 87:44]
  wire [9:0] _isForwardData_T_8 = {addr_index,addr_wordIndex}; // @[src/main/scala/nutcore/mem/Cache.scala 78:35]
  wire  _isForwardData_T_10 = io_dataWriteBus_req_valid & io_dataWriteBus_req_bits_setIdx == _isForwardData_T_8; // @[src/main/scala/nutcore/mem/Cache.scala 217:13]
  wire  isForwardData = io_in_valid & _isForwardData_T_10; // @[src/main/scala/nutcore/mem/Cache.scala 216:35]
  reg  isForwardDataReg; // @[src/main/scala/nutcore/mem/Cache.scala 219:33]
  wire  _GEN_8 = isForwardData | isForwardDataReg; // @[src/main/scala/nutcore/mem/Cache.scala 220:24 219:33 220:43]
  reg [63:0] forwardDataReg_data_data; // @[src/main/scala/nutcore/mem/Cache.scala 222:33]
  reg [3:0] forwardDataReg_waymask; // @[src/main/scala/nutcore/mem/Cache.scala 222:33]
  wire  _io_in_ready_T_1 = io_out_ready & io_out_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  reg [63:0] c_11; // @[src/main/scala/utils/GTimer.scala 24:20]
  wire [63:0] _c_T_23 = c_11 + 64'h1; // @[src/main/scala/utils/GTimer.scala 25:12]
  reg [63:0] c_12; // @[src/main/scala/utils/GTimer.scala 24:20]
  wire [63:0] _c_T_25 = c_12 + 64'h1; // @[src/main/scala/utils/GTimer.scala 25:12]
  wire  _GEN_13 = _T_13 & DISPLAY_ENABLE; // @[src/main/scala/utils/Debug.scala 56:24]
  assign io_in_ready = _T_1 | _io_in_ready_T_1; // @[src/main/scala/nutcore/mem/Cache.scala 228:31]
  assign io_out_valid = io_in_valid; // @[src/main/scala/nutcore/mem/Cache.scala 227:16]
  assign io_out_bits_req_addr = io_in_bits_req_addr; // @[src/main/scala/nutcore/mem/Cache.scala 226:19]
  assign io_out_bits_req_size = io_in_bits_req_size; // @[src/main/scala/nutcore/mem/Cache.scala 226:19]
  assign io_out_bits_req_cmd = io_in_bits_req_cmd; // @[src/main/scala/nutcore/mem/Cache.scala 226:19]
  assign io_out_bits_req_wmask = io_in_bits_req_wmask; // @[src/main/scala/nutcore/mem/Cache.scala 226:19]
  assign io_out_bits_req_wdata = io_in_bits_req_wdata; // @[src/main/scala/nutcore/mem/Cache.scala 226:19]
  assign io_out_bits_metas_0_tag = pickForwardMeta & forwardWaymask_0 ? _GEN_3 : io_metaReadResp_0_tag; // @[src/main/scala/nutcore/mem/Cache.scala 187:22]
  assign io_out_bits_metas_0_valid = pickForwardMeta & forwardWaymask_0 | io_metaReadResp_0_valid; // @[src/main/scala/nutcore/mem/Cache.scala 187:22]
  assign io_out_bits_metas_0_dirty = pickForwardMeta & forwardWaymask_0 ? _GEN_5 : io_metaReadResp_0_dirty; // @[src/main/scala/nutcore/mem/Cache.scala 187:22]
  assign io_out_bits_metas_1_tag = pickForwardMeta & forwardWaymask_1 ? _GEN_3 : io_metaReadResp_1_tag; // @[src/main/scala/nutcore/mem/Cache.scala 187:22]
  assign io_out_bits_metas_1_valid = pickForwardMeta & forwardWaymask_1 | io_metaReadResp_1_valid; // @[src/main/scala/nutcore/mem/Cache.scala 187:22]
  assign io_out_bits_metas_1_dirty = pickForwardMeta & forwardWaymask_1 ? _GEN_5 : io_metaReadResp_1_dirty; // @[src/main/scala/nutcore/mem/Cache.scala 187:22]
  assign io_out_bits_metas_2_tag = pickForwardMeta & forwardWaymask_2 ? _GEN_3 : io_metaReadResp_2_tag; // @[src/main/scala/nutcore/mem/Cache.scala 187:22]
  assign io_out_bits_metas_2_valid = pickForwardMeta & forwardWaymask_2 | io_metaReadResp_2_valid; // @[src/main/scala/nutcore/mem/Cache.scala 187:22]
  assign io_out_bits_metas_2_dirty = pickForwardMeta & forwardWaymask_2 ? _GEN_5 : io_metaReadResp_2_dirty; // @[src/main/scala/nutcore/mem/Cache.scala 187:22]
  assign io_out_bits_metas_3_tag = pickForwardMeta & forwardWaymask_3 ? _GEN_3 : io_metaReadResp_3_tag; // @[src/main/scala/nutcore/mem/Cache.scala 187:22]
  assign io_out_bits_metas_3_valid = pickForwardMeta & forwardWaymask_3 | io_metaReadResp_3_valid; // @[src/main/scala/nutcore/mem/Cache.scala 187:22]
  assign io_out_bits_metas_3_dirty = pickForwardMeta & forwardWaymask_3 ? _GEN_5 : io_metaReadResp_3_dirty; // @[src/main/scala/nutcore/mem/Cache.scala 187:22]
  assign io_out_bits_datas_0_data = io_dataReadResp_0_data; // @[src/main/scala/nutcore/mem/Cache.scala 213:21]
  assign io_out_bits_datas_1_data = io_dataReadResp_1_data; // @[src/main/scala/nutcore/mem/Cache.scala 213:21]
  assign io_out_bits_datas_2_data = io_dataReadResp_2_data; // @[src/main/scala/nutcore/mem/Cache.scala 213:21]
  assign io_out_bits_datas_3_data = io_dataReadResp_3_data; // @[src/main/scala/nutcore/mem/Cache.scala 213:21]
  assign io_out_bits_hit = io_in_valid & |hitVec; // @[src/main/scala/nutcore/mem/Cache.scala 211:34]
  assign io_out_bits_waymask = io_out_bits_hit ? hitVec : _waymask_T; // @[src/main/scala/nutcore/mem/Cache.scala 200:20]
  assign io_out_bits_mmio = _io_out_bits_mmio_T_2 | _io_out_bits_mmio_T_5; // @[src/main/scala/nutcore/NutCore.scala 88:15]
  assign io_out_bits_isForwardData = isForwardDataReg | isForwardData; // @[src/main/scala/nutcore/mem/Cache.scala 223:49]
  assign io_out_bits_forwardData_data_data = isForwardData ? io_dataWriteBus_req_bits_data_data :
    forwardDataReg_data_data; // @[src/main/scala/nutcore/mem/Cache.scala 224:33]
  assign io_out_bits_forwardData_waymask = isForwardData ? io_dataWriteBus_req_bits_waymask : forwardDataReg_waymask; // @[src/main/scala/nutcore/mem/Cache.scala 224:33]
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/nutcore/mem/Cache.scala 177:33]
      isForwardMetaReg <= 1'h0; // @[src/main/scala/nutcore/mem/Cache.scala 177:33]
    end else if (_T | ~io_in_valid) begin // @[src/main/scala/nutcore/mem/Cache.scala 179:37]
      isForwardMetaReg <= 1'h0; // @[src/main/scala/nutcore/mem/Cache.scala 179:56]
    end else begin
      isForwardMetaReg <= _GEN_0;
    end
    if (isForwardMeta) begin // @[src/main/scala/nutcore/mem/Cache.scala 180:33]
      forwardMetaReg_data_tag <= io_metaWriteBus_req_bits_data_tag; // @[src/main/scala/nutcore/mem/Cache.scala 180:33]
    end
    if (isForwardMeta) begin // @[src/main/scala/nutcore/mem/Cache.scala 180:33]
      forwardMetaReg_data_dirty <= io_metaWriteBus_req_bits_data_dirty; // @[src/main/scala/nutcore/mem/Cache.scala 180:33]
    end
    if (isForwardMeta) begin // @[src/main/scala/nutcore/mem/Cache.scala 180:33]
      forwardMetaReg_waymask <= io_metaWriteBus_req_bits_waymask; // @[src/main/scala/nutcore/mem/Cache.scala 180:33]
    end
    if (reset) begin // @[src/main/scala/utils/LFSR64.scala 25:23]
      victimWaymask_lfsr <= 64'h1234567887654321; // @[src/main/scala/utils/LFSR64.scala 25:23]
    end else if (victimWaymask_lfsr == 64'h0) begin // @[src/main/scala/utils/LFSR64.scala 28:18]
      victimWaymask_lfsr <= 64'h1;
    end else begin
      victimWaymask_lfsr <= _victimWaymask_lfsr_T_2;
    end
    if (reset) begin // @[src/main/scala/utils/GTimer.scala 24:20]
      c <= 64'h0; // @[src/main/scala/utils/GTimer.scala 24:20]
    end else begin
      c <= _c_T_1; // @[src/main/scala/utils/GTimer.scala 25:7]
    end
    if (reset) begin // @[src/main/scala/utils/GTimer.scala 24:20]
      c_1 <= 64'h0; // @[src/main/scala/utils/GTimer.scala 24:20]
    end else begin
      c_1 <= _c_T_3; // @[src/main/scala/utils/GTimer.scala 25:7]
    end
    if (reset) begin // @[src/main/scala/utils/GTimer.scala 24:20]
      c_2 <= 64'h0; // @[src/main/scala/utils/GTimer.scala 24:20]
    end else begin
      c_2 <= _c_T_5; // @[src/main/scala/utils/GTimer.scala 25:7]
    end
    if (reset) begin // @[src/main/scala/utils/GTimer.scala 24:20]
      c_3 <= 64'h0; // @[src/main/scala/utils/GTimer.scala 24:20]
    end else begin
      c_3 <= _c_T_7; // @[src/main/scala/utils/GTimer.scala 25:7]
    end
    if (reset) begin // @[src/main/scala/utils/GTimer.scala 24:20]
      c_4 <= 64'h0; // @[src/main/scala/utils/GTimer.scala 24:20]
    end else begin
      c_4 <= _c_T_9; // @[src/main/scala/utils/GTimer.scala 25:7]
    end
    if (reset) begin // @[src/main/scala/utils/GTimer.scala 24:20]
      c_5 <= 64'h0; // @[src/main/scala/utils/GTimer.scala 24:20]
    end else begin
      c_5 <= _c_T_11; // @[src/main/scala/utils/GTimer.scala 25:7]
    end
    if (reset) begin // @[src/main/scala/utils/GTimer.scala 24:20]
      c_6 <= 64'h0; // @[src/main/scala/utils/GTimer.scala 24:20]
    end else begin
      c_6 <= _c_T_13; // @[src/main/scala/utils/GTimer.scala 25:7]
    end
    if (reset) begin // @[src/main/scala/utils/GTimer.scala 24:20]
      c_7 <= 64'h0; // @[src/main/scala/utils/GTimer.scala 24:20]
    end else begin
      c_7 <= _c_T_15; // @[src/main/scala/utils/GTimer.scala 25:7]
    end
    if (reset) begin // @[src/main/scala/utils/GTimer.scala 24:20]
      c_8 <= 64'h0; // @[src/main/scala/utils/GTimer.scala 24:20]
    end else begin
      c_8 <= _c_T_17; // @[src/main/scala/utils/GTimer.scala 25:7]
    end
    if (reset) begin // @[src/main/scala/utils/GTimer.scala 24:20]
      c_9 <= 64'h0; // @[src/main/scala/utils/GTimer.scala 24:20]
    end else begin
      c_9 <= _c_T_19; // @[src/main/scala/utils/GTimer.scala 25:7]
    end
    if (reset) begin // @[src/main/scala/utils/GTimer.scala 24:20]
      c_10 <= 64'h0; // @[src/main/scala/utils/GTimer.scala 24:20]
    end else begin
      c_10 <= _c_T_21; // @[src/main/scala/utils/GTimer.scala 25:7]
    end
    if (reset) begin // @[src/main/scala/nutcore/mem/Cache.scala 219:33]
      isForwardDataReg <= 1'h0; // @[src/main/scala/nutcore/mem/Cache.scala 219:33]
    end else if (_T_2) begin // @[src/main/scala/nutcore/mem/Cache.scala 221:37]
      isForwardDataReg <= 1'h0; // @[src/main/scala/nutcore/mem/Cache.scala 221:56]
    end else begin
      isForwardDataReg <= _GEN_8;
    end
    if (isForwardData) begin // @[src/main/scala/nutcore/mem/Cache.scala 222:33]
      forwardDataReg_data_data <= io_dataWriteBus_req_bits_data_data; // @[src/main/scala/nutcore/mem/Cache.scala 222:33]
    end
    if (isForwardData) begin // @[src/main/scala/nutcore/mem/Cache.scala 222:33]
      forwardDataReg_waymask <= io_dataWriteBus_req_bits_waymask; // @[src/main/scala/nutcore/mem/Cache.scala 222:33]
    end
    if (reset) begin // @[src/main/scala/utils/GTimer.scala 24:20]
      c_11 <= 64'h0; // @[src/main/scala/utils/GTimer.scala 24:20]
    end else begin
      c_11 <= _c_T_23; // @[src/main/scala/utils/GTimer.scala 25:7]
    end
    if (reset) begin // @[src/main/scala/utils/GTimer.scala 24:20]
      c_12 <= 64'h0; // @[src/main/scala/utils/GTimer.scala 24:20]
    end else begin
      c_12 <= _c_T_25; // @[src/main/scala/utils/GTimer.scala 25:7]
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_13 & DISPLAY_ENABLE & ~reset) begin
          $fwrite(32'h80000002,"[%d] CacheStage2_1: ",c); // @[src/main/scala/utils/Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_13 & _T_16) begin
          $fwrite(32'h80000002,"[ERROR] metaWay %x metat %x reqt %x\n",metaWay_0_valid,metaWay_0_tag,addr_tag); // @[src/main/scala/utils/Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_13 & DISPLAY_ENABLE & ~reset) begin
          $fwrite(32'h80000002,"[%d] CacheStage2_1: ",c_1); // @[src/main/scala/utils/Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_13 & _T_16) begin
          $fwrite(32'h80000002,"[ERROR] metaWay %x metat %x reqt %x\n",metaWay_1_valid,metaWay_1_tag,addr_tag); // @[src/main/scala/utils/Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_13 & DISPLAY_ENABLE & ~reset) begin
          $fwrite(32'h80000002,"[%d] CacheStage2_1: ",c_2); // @[src/main/scala/utils/Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_13 & _T_16) begin
          $fwrite(32'h80000002,"[ERROR] metaWay %x metat %x reqt %x\n",metaWay_2_valid,metaWay_2_tag,addr_tag); // @[src/main/scala/utils/Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_13 & DISPLAY_ENABLE & ~reset) begin
          $fwrite(32'h80000002,"[%d] CacheStage2_1: ",c_3); // @[src/main/scala/utils/Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_13 & _T_16) begin
          $fwrite(32'h80000002,"[ERROR] metaWay %x metat %x reqt %x\n",metaWay_3_valid,metaWay_3_tag,addr_tag); // @[src/main/scala/utils/Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_13 & DISPLAY_ENABLE & ~reset) begin
          $fwrite(32'h80000002,"[%d] CacheStage2_1: ",c_4); // @[src/main/scala/utils/Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_13 & _T_16) begin
          $fwrite(32'h80000002,"[ERROR] metaReadResp %x metat %x reqt %x\n",io_metaReadResp_0_valid,
            io_metaReadResp_0_tag,addr_tag); // @[src/main/scala/utils/Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_13 & DISPLAY_ENABLE & ~reset) begin
          $fwrite(32'h80000002,"[%d] CacheStage2_1: ",c_5); // @[src/main/scala/utils/Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_13 & _T_16) begin
          $fwrite(32'h80000002,"[ERROR] metaReadResp %x metat %x reqt %x\n",io_metaReadResp_1_valid,
            io_metaReadResp_1_tag,addr_tag); // @[src/main/scala/utils/Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_13 & DISPLAY_ENABLE & ~reset) begin
          $fwrite(32'h80000002,"[%d] CacheStage2_1: ",c_6); // @[src/main/scala/utils/Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_13 & _T_16) begin
          $fwrite(32'h80000002,"[ERROR] metaReadResp %x metat %x reqt %x\n",io_metaReadResp_2_valid,
            io_metaReadResp_2_tag,addr_tag); // @[src/main/scala/utils/Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_13 & DISPLAY_ENABLE & ~reset) begin
          $fwrite(32'h80000002,"[%d] CacheStage2_1: ",c_7); // @[src/main/scala/utils/Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_13 & _T_16) begin
          $fwrite(32'h80000002,"[ERROR] metaReadResp %x metat %x reqt %x\n",io_metaReadResp_3_valid,
            io_metaReadResp_3_tag,addr_tag); // @[src/main/scala/utils/Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_13 & DISPLAY_ENABLE & ~reset) begin
          $fwrite(32'h80000002,"[%d] CacheStage2_1: ",c_8); // @[src/main/scala/utils/Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_13 & _T_16) begin
          $fwrite(32'h80000002,"[ERROR] forwardMetaReg isForwardMetaReg %x %x metat %x wm %b\n",isForwardMetaReg,1'h1,
            forwardMetaReg_data_tag,forwardMetaReg_waymask); // @[src/main/scala/utils/Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_13 & DISPLAY_ENABLE & ~reset) begin
          $fwrite(32'h80000002,"[%d] CacheStage2_1: ",c_9); // @[src/main/scala/utils/Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_13 & _T_16) begin
          $fwrite(32'h80000002,"[ERROR] forwardMeta isForwardMeta %x %x metat %x wm %b\n",isForwardMeta,1'h1,
            io_metaWriteBus_req_bits_data_tag,io_metaWriteBus_req_bits_waymask); // @[src/main/scala/utils/Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_13 & DISPLAY_ENABLE & ~reset) begin
          $fwrite(32'h80000002,"[%d] CacheStage2_1: ",c_10); // @[src/main/scala/utils/Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_13 & _T_16) begin
          $fwrite(32'h80000002,"[ERROR] hit %b wmask %b hitvec %b\n",io_out_bits_hit,_GEN_6,hitVec); // @[src/main/scala/utils/Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_16 & ~(~(io_in_valid & _T_13))) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Cache.scala:208 assert(!(io.in.valid && PopCount(waymask) > 1.U))\n"); // @[src/main/scala/nutcore/mem/Cache.scala 208:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~(io_in_valid & _T_13)) & _T_16) begin
          $fatal; // @[src/main/scala/nutcore/mem/Cache.scala 208:9]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & ~reset) begin
          $fwrite(32'h80000002,"[%d] CacheStage2_1: ",c_11); // @[src/main/scala/utils/Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_16) begin
          $fwrite(32'h80000002,"[isFD:%d isFDreg:%d inFire:%d invalid:%d \n",isForwardData,isForwardDataReg,_T,
            io_in_valid); // @[src/main/scala/utils/Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & ~reset) begin
          $fwrite(32'h80000002,"[%d] CacheStage2_1: ",c_12); // @[src/main/scala/utils/Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_16) begin
          $fwrite(32'h80000002,"[isFM:%d isFMreg:%d metawreq:%x widx:%x ridx:%x \n",isForwardMeta,isForwardMetaReg,
            io_metaWriteBus_req_valid,io_metaWriteBus_req_bits_setIdx,addr_index); // @[src/main/scala/utils/Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  isForwardMetaReg = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  forwardMetaReg_data_tag = _RAND_1[18:0];
  _RAND_2 = {1{`RANDOM}};
  forwardMetaReg_data_dirty = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  forwardMetaReg_waymask = _RAND_3[3:0];
  _RAND_4 = {2{`RANDOM}};
  victimWaymask_lfsr = _RAND_4[63:0];
  _RAND_5 = {2{`RANDOM}};
  c = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  c_1 = _RAND_6[63:0];
  _RAND_7 = {2{`RANDOM}};
  c_2 = _RAND_7[63:0];
  _RAND_8 = {2{`RANDOM}};
  c_3 = _RAND_8[63:0];
  _RAND_9 = {2{`RANDOM}};
  c_4 = _RAND_9[63:0];
  _RAND_10 = {2{`RANDOM}};
  c_5 = _RAND_10[63:0];
  _RAND_11 = {2{`RANDOM}};
  c_6 = _RAND_11[63:0];
  _RAND_12 = {2{`RANDOM}};
  c_7 = _RAND_12[63:0];
  _RAND_13 = {2{`RANDOM}};
  c_8 = _RAND_13[63:0];
  _RAND_14 = {2{`RANDOM}};
  c_9 = _RAND_14[63:0];
  _RAND_15 = {2{`RANDOM}};
  c_10 = _RAND_15[63:0];
  _RAND_16 = {1{`RANDOM}};
  isForwardDataReg = _RAND_16[0:0];
  _RAND_17 = {2{`RANDOM}};
  forwardDataReg_data_data = _RAND_17[63:0];
  _RAND_18 = {1{`RANDOM}};
  forwardDataReg_waymask = _RAND_18[3:0];
  _RAND_19 = {2{`RANDOM}};
  c_11 = _RAND_19[63:0];
  _RAND_20 = {2{`RANDOM}};
  c_12 = _RAND_20[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module CacheStage3_1(
  input         clock,
  input         reset,
  output        io_in_ready, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  input         io_in_valid, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  input  [31:0] io_in_bits_req_addr, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  input  [2:0]  io_in_bits_req_size, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  input  [3:0]  io_in_bits_req_cmd, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  input  [7:0]  io_in_bits_req_wmask, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  input  [63:0] io_in_bits_req_wdata, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  input  [18:0] io_in_bits_metas_0_tag, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  input         io_in_bits_metas_0_valid, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  input         io_in_bits_metas_0_dirty, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  input  [18:0] io_in_bits_metas_1_tag, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  input         io_in_bits_metas_1_valid, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  input         io_in_bits_metas_1_dirty, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  input  [18:0] io_in_bits_metas_2_tag, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  input         io_in_bits_metas_2_valid, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  input         io_in_bits_metas_2_dirty, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  input  [18:0] io_in_bits_metas_3_tag, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  input         io_in_bits_metas_3_valid, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  input         io_in_bits_metas_3_dirty, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  input  [63:0] io_in_bits_datas_0_data, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  input  [63:0] io_in_bits_datas_1_data, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  input  [63:0] io_in_bits_datas_2_data, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  input  [63:0] io_in_bits_datas_3_data, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  input         io_in_bits_hit, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  input  [3:0]  io_in_bits_waymask, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  input         io_in_bits_mmio, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  input         io_in_bits_isForwardData, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  input  [63:0] io_in_bits_forwardData_data_data, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  input  [3:0]  io_in_bits_forwardData_waymask, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  input         io_out_ready, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  output        io_out_valid, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  output [3:0]  io_out_bits_cmd, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  output [63:0] io_out_bits_rdata, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  output        io_isFinish, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  input         io_dataReadBus_req_ready, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  output        io_dataReadBus_req_valid, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  output [9:0]  io_dataReadBus_req_bits_setIdx, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  input  [63:0] io_dataReadBus_resp_data_0_data, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  input  [63:0] io_dataReadBus_resp_data_1_data, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  input  [63:0] io_dataReadBus_resp_data_2_data, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  input  [63:0] io_dataReadBus_resp_data_3_data, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  output        io_dataWriteBus_req_valid, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  output [9:0]  io_dataWriteBus_req_bits_setIdx, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  output [63:0] io_dataWriteBus_req_bits_data_data, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  output [3:0]  io_dataWriteBus_req_bits_waymask, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  output        io_metaWriteBus_req_valid, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  output [6:0]  io_metaWriteBus_req_bits_setIdx, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  output [18:0] io_metaWriteBus_req_bits_data_tag, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  output        io_metaWriteBus_req_bits_data_valid, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  output        io_metaWriteBus_req_bits_data_dirty, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  output [3:0]  io_metaWriteBus_req_bits_waymask, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  input         io_mem_req_ready, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  output        io_mem_req_valid, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  output [31:0] io_mem_req_bits_addr, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  output [2:0]  io_mem_req_bits_size, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  output [3:0]  io_mem_req_bits_cmd, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  output [7:0]  io_mem_req_bits_wmask, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  output [63:0] io_mem_req_bits_wdata, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  output        io_mem_resp_ready, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  input         io_mem_resp_valid, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  input  [3:0]  io_mem_resp_bits_cmd, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  input  [63:0] io_mem_resp_bits_rdata, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  input         io_mmio_req_ready, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  output        io_mmio_req_valid, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  output [31:0] io_mmio_req_bits_addr, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  output [2:0]  io_mmio_req_bits_size, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  output [3:0]  io_mmio_req_bits_cmd, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  output [7:0]  io_mmio_req_bits_wmask, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  output [63:0] io_mmio_req_bits_wdata, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  output        io_mmio_resp_ready, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  input         io_mmio_resp_valid, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  input  [63:0] io_mmio_resp_bits_rdata, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  output        io_cohResp_valid, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  output [3:0]  io_cohResp_bits_cmd, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  output [63:0] io_cohResp_bits_rdata, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  output        io_dataReadRespToL1, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  input         DISPLAY_ENABLE,
  output        _WIRE_19
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [63:0] _RAND_14;
  reg [63:0] _RAND_15;
  reg [63:0] _RAND_16;
  reg [63:0] _RAND_17;
  reg [63:0] _RAND_18;
  reg [63:0] _RAND_19;
  reg [63:0] _RAND_20;
  reg [63:0] _RAND_21;
  reg [63:0] _RAND_22;
  reg [63:0] _RAND_23;
  reg [63:0] _RAND_24;
  reg [63:0] _RAND_25;
`endif // RANDOMIZE_REG_INIT
  wire  metaWriteArb_io_in_0_valid; // @[src/main/scala/nutcore/mem/Cache.scala 254:28]
  wire [6:0] metaWriteArb_io_in_0_bits_setIdx; // @[src/main/scala/nutcore/mem/Cache.scala 254:28]
  wire [18:0] metaWriteArb_io_in_0_bits_data_tag; // @[src/main/scala/nutcore/mem/Cache.scala 254:28]
  wire  metaWriteArb_io_in_0_bits_data_dirty; // @[src/main/scala/nutcore/mem/Cache.scala 254:28]
  wire [3:0] metaWriteArb_io_in_0_bits_waymask; // @[src/main/scala/nutcore/mem/Cache.scala 254:28]
  wire  metaWriteArb_io_in_1_valid; // @[src/main/scala/nutcore/mem/Cache.scala 254:28]
  wire [6:0] metaWriteArb_io_in_1_bits_setIdx; // @[src/main/scala/nutcore/mem/Cache.scala 254:28]
  wire [18:0] metaWriteArb_io_in_1_bits_data_tag; // @[src/main/scala/nutcore/mem/Cache.scala 254:28]
  wire  metaWriteArb_io_in_1_bits_data_dirty; // @[src/main/scala/nutcore/mem/Cache.scala 254:28]
  wire [3:0] metaWriteArb_io_in_1_bits_waymask; // @[src/main/scala/nutcore/mem/Cache.scala 254:28]
  wire  metaWriteArb_io_out_valid; // @[src/main/scala/nutcore/mem/Cache.scala 254:28]
  wire [6:0] metaWriteArb_io_out_bits_setIdx; // @[src/main/scala/nutcore/mem/Cache.scala 254:28]
  wire [18:0] metaWriteArb_io_out_bits_data_tag; // @[src/main/scala/nutcore/mem/Cache.scala 254:28]
  wire  metaWriteArb_io_out_bits_data_dirty; // @[src/main/scala/nutcore/mem/Cache.scala 254:28]
  wire [3:0] metaWriteArb_io_out_bits_waymask; // @[src/main/scala/nutcore/mem/Cache.scala 254:28]
  wire  dataWriteArb_io_in_0_valid; // @[src/main/scala/nutcore/mem/Cache.scala 255:28]
  wire [9:0] dataWriteArb_io_in_0_bits_setIdx; // @[src/main/scala/nutcore/mem/Cache.scala 255:28]
  wire [63:0] dataWriteArb_io_in_0_bits_data_data; // @[src/main/scala/nutcore/mem/Cache.scala 255:28]
  wire [3:0] dataWriteArb_io_in_0_bits_waymask; // @[src/main/scala/nutcore/mem/Cache.scala 255:28]
  wire  dataWriteArb_io_in_1_valid; // @[src/main/scala/nutcore/mem/Cache.scala 255:28]
  wire [9:0] dataWriteArb_io_in_1_bits_setIdx; // @[src/main/scala/nutcore/mem/Cache.scala 255:28]
  wire [63:0] dataWriteArb_io_in_1_bits_data_data; // @[src/main/scala/nutcore/mem/Cache.scala 255:28]
  wire [3:0] dataWriteArb_io_in_1_bits_waymask; // @[src/main/scala/nutcore/mem/Cache.scala 255:28]
  wire  dataWriteArb_io_out_valid; // @[src/main/scala/nutcore/mem/Cache.scala 255:28]
  wire [9:0] dataWriteArb_io_out_bits_setIdx; // @[src/main/scala/nutcore/mem/Cache.scala 255:28]
  wire [63:0] dataWriteArb_io_out_bits_data_data; // @[src/main/scala/nutcore/mem/Cache.scala 255:28]
  wire [3:0] dataWriteArb_io_out_bits_waymask; // @[src/main/scala/nutcore/mem/Cache.scala 255:28]
  wire [2:0] addr_wordIndex = io_in_bits_req_addr[5:3]; // @[src/main/scala/nutcore/mem/Cache.scala 258:31]
  wire [6:0] addr_index = io_in_bits_req_addr[12:6]; // @[src/main/scala/nutcore/mem/Cache.scala 258:31]
  wire [18:0] addr_tag = io_in_bits_req_addr[31:13]; // @[src/main/scala/nutcore/mem/Cache.scala 258:31]
  wire  mmio = io_in_valid & io_in_bits_mmio; // @[src/main/scala/nutcore/mem/Cache.scala 259:26]
  wire  hit = io_in_valid & io_in_bits_hit; // @[src/main/scala/nutcore/mem/Cache.scala 260:25]
  wire  miss = io_in_valid & ~io_in_bits_hit; // @[src/main/scala/nutcore/mem/Cache.scala 261:26]
  wire  _probe_T_1 = io_in_bits_req_cmd == 4'h8; // @[src/main/scala/bus/simplebus/SimpleBus.scala 79:23]
  wire  probe = io_in_valid & _probe_T_1; // @[src/main/scala/nutcore/mem/Cache.scala 262:39]
  wire  _hitReadBurst_T = io_in_bits_req_cmd == 4'h2; // @[src/main/scala/bus/simplebus/SimpleBus.scala 76:27]
  wire  hitReadBurst = hit & _hitReadBurst_T; // @[src/main/scala/nutcore/mem/Cache.scala 263:26]
  wire  meta_dirty = io_in_bits_waymask[0] & io_in_bits_metas_0_dirty | io_in_bits_waymask[1] & io_in_bits_metas_1_dirty
     | io_in_bits_waymask[2] & io_in_bits_metas_2_dirty | io_in_bits_waymask[3] & io_in_bits_metas_3_dirty; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [18:0] _meta_T_18 = io_in_bits_waymask[0] ? io_in_bits_metas_0_tag : 19'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [18:0] _meta_T_19 = io_in_bits_waymask[1] ? io_in_bits_metas_1_tag : 19'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [18:0] _meta_T_20 = io_in_bits_waymask[2] ? io_in_bits_metas_2_tag : 19'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [18:0] _meta_T_21 = io_in_bits_waymask[3] ? io_in_bits_metas_3_tag : 19'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [18:0] _meta_T_22 = _meta_T_18 | _meta_T_19; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [18:0] _meta_T_23 = _meta_T_22 | _meta_T_20; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [18:0] meta_tag = _meta_T_23 | _meta_T_21; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _T_3 = ~reset; // @[src/main/scala/nutcore/mem/Cache.scala 265:9]
  wire  useForwardData = io_in_bits_isForwardData & io_in_bits_waymask == io_in_bits_forwardData_waymask; // @[src/main/scala/nutcore/mem/Cache.scala 273:49]
  wire [63:0] _dataReadArray_T_4 = io_in_bits_waymask[0] ? io_in_bits_datas_0_data : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _dataReadArray_T_5 = io_in_bits_waymask[1] ? io_in_bits_datas_1_data : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _dataReadArray_T_6 = io_in_bits_waymask[2] ? io_in_bits_datas_2_data : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _dataReadArray_T_7 = io_in_bits_waymask[3] ? io_in_bits_datas_3_data : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _dataReadArray_T_8 = _dataReadArray_T_4 | _dataReadArray_T_5; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _dataReadArray_T_9 = _dataReadArray_T_8 | _dataReadArray_T_6; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _dataReadArray_T_10 = _dataReadArray_T_9 | _dataReadArray_T_7; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] dataRead = useForwardData ? io_in_bits_forwardData_data_data : _dataReadArray_T_10; // @[src/main/scala/nutcore/mem/Cache.scala 275:21]
  wire [7:0] _wordMask_T_12 = io_in_bits_req_wmask[0] ? 8'hff : 8'h0; // @[src/main/scala/utils/BitUtils.scala 27:45]
  wire [7:0] _wordMask_T_14 = io_in_bits_req_wmask[1] ? 8'hff : 8'h0; // @[src/main/scala/utils/BitUtils.scala 27:45]
  wire [7:0] _wordMask_T_16 = io_in_bits_req_wmask[2] ? 8'hff : 8'h0; // @[src/main/scala/utils/BitUtils.scala 27:45]
  wire [7:0] _wordMask_T_18 = io_in_bits_req_wmask[3] ? 8'hff : 8'h0; // @[src/main/scala/utils/BitUtils.scala 27:45]
  wire [7:0] _wordMask_T_20 = io_in_bits_req_wmask[4] ? 8'hff : 8'h0; // @[src/main/scala/utils/BitUtils.scala 27:45]
  wire [7:0] _wordMask_T_22 = io_in_bits_req_wmask[5] ? 8'hff : 8'h0; // @[src/main/scala/utils/BitUtils.scala 27:45]
  wire [7:0] _wordMask_T_24 = io_in_bits_req_wmask[6] ? 8'hff : 8'h0; // @[src/main/scala/utils/BitUtils.scala 27:45]
  wire [7:0] _wordMask_T_26 = io_in_bits_req_wmask[7] ? 8'hff : 8'h0; // @[src/main/scala/utils/BitUtils.scala 27:45]
  wire [63:0] _wordMask_T_27 = {_wordMask_T_26,_wordMask_T_24,_wordMask_T_22,_wordMask_T_20,_wordMask_T_18,
    _wordMask_T_16,_wordMask_T_14,_wordMask_T_12}; // @[src/main/scala/utils/BitUtils.scala 27:26]
  wire [63:0] wordMask = io_in_bits_req_cmd[0] ? _wordMask_T_27 : 64'h0; // @[src/main/scala/nutcore/mem/Cache.scala 276:21]
  reg [2:0] writeL2BeatCnt_value; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
  wire  _T_5 = io_out_ready & io_out_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  wire  _T_6 = io_in_bits_req_cmd == 4'h3; // @[src/main/scala/nutcore/mem/Cache.scala 279:32]
  wire  _T_7 = io_in_bits_req_cmd == 4'h7; // @[src/main/scala/bus/simplebus/SimpleBus.scala 78:27]
  wire  _T_8 = io_in_bits_req_cmd == 4'h3 | _T_7; // @[src/main/scala/nutcore/mem/Cache.scala 279:60]
  wire [2:0] _value_T_1 = writeL2BeatCnt_value + 3'h1; // @[src/main/scala/chisel3/util/Counter.scala 77:24]
  wire [2:0] _GEN_0 = _T_5 & (io_in_bits_req_cmd == 4'h3 | _T_7) ? _value_T_1 : writeL2BeatCnt_value; // @[src/main/scala/nutcore/mem/Cache.scala 279:83 src/main/scala/chisel3/util/Counter.scala 77:15 61:40]
  wire  hitWrite = hit & io_in_bits_req_cmd[0]; // @[src/main/scala/nutcore/mem/Cache.scala 283:22]
  wire [63:0] _dataHitWriteBus_x1_T = io_in_bits_req_wdata & wordMask; // @[src/main/scala/utils/BitUtils.scala 34:14]
  wire [63:0] _dataHitWriteBus_x1_T_1 = ~wordMask; // @[src/main/scala/utils/BitUtils.scala 34:39]
  wire [63:0] _dataHitWriteBus_x1_T_2 = dataRead & _dataHitWriteBus_x1_T_1; // @[src/main/scala/utils/BitUtils.scala 34:37]
  wire [63:0] dataHitWriteBus_x1_data = _dataHitWriteBus_x1_T | _dataHitWriteBus_x1_T_2; // @[src/main/scala/utils/BitUtils.scala 34:26]
  wire [2:0] _dataHitWriteBus_x3_T_3 = _T_8 ? writeL2BeatCnt_value : addr_wordIndex; // @[src/main/scala/nutcore/mem/Cache.scala 286:51]
  wire [9:0] dataHitWriteBus_x3 = {addr_index,_dataHitWriteBus_x3_T_3}; // @[src/main/scala/nutcore/mem/Cache.scala 286:35]
  wire  metaHitWriteBus_x5 = hitWrite & ~meta_dirty; // @[src/main/scala/nutcore/mem/Cache.scala 289:22]
  reg [3:0] state; // @[src/main/scala/nutcore/mem/Cache.scala 294:22]
  reg [2:0] readBeatCnt_value; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
  reg [2:0] writeBeatCnt_value; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
  reg [1:0] state2; // @[src/main/scala/nutcore/mem/Cache.scala 304:23]
  wire  _T_14 = state == 4'h3; // @[src/main/scala/nutcore/mem/Cache.scala 306:39]
  wire  _T_15 = state == 4'h8; // @[src/main/scala/nutcore/mem/Cache.scala 306:66]
  wire [2:0] _T_20 = _T_15 ? readBeatCnt_value : writeBeatCnt_value; // @[src/main/scala/nutcore/mem/Cache.scala 307:33]
  reg [63:0] dataWay_0_data; // @[src/main/scala/nutcore/mem/Cache.scala 308:26]
  reg [63:0] dataWay_1_data; // @[src/main/scala/nutcore/mem/Cache.scala 308:26]
  reg [63:0] dataWay_2_data; // @[src/main/scala/nutcore/mem/Cache.scala 308:26]
  reg [63:0] dataWay_3_data; // @[src/main/scala/nutcore/mem/Cache.scala 308:26]
  wire [63:0] _dataHitWay_T_4 = io_in_bits_waymask[0] ? dataWay_0_data : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _dataHitWay_T_5 = io_in_bits_waymask[1] ? dataWay_1_data : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _dataHitWay_T_6 = io_in_bits_waymask[2] ? dataWay_2_data : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _dataHitWay_T_7 = io_in_bits_waymask[3] ? dataWay_3_data : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _dataHitWay_T_8 = _dataHitWay_T_4 | _dataHitWay_T_5; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _dataHitWay_T_9 = _dataHitWay_T_8 | _dataHitWay_T_6; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _T_23 = io_dataReadBus_req_ready & io_dataReadBus_req_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  wire  _T_26 = io_mem_req_ready & io_mem_req_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  wire  _T_29 = hitReadBurst & io_out_ready; // @[src/main/scala/nutcore/mem/Cache.scala 314:79]
  wire [1:0] _GEN_8 = _T_26 | io_cohResp_valid | hitReadBurst & io_out_ready ? 2'h0 : state2; // @[src/main/scala/nutcore/mem/Cache.scala 314:105 304:23 314:96]
  wire [31:0] raddr = {io_in_bits_req_addr[31:3],3'h0}; // @[src/main/scala/nutcore/mem/Cache.scala 318:35]
  wire [31:0] waddr = {meta_tag,addr_index,6'h0}; // @[src/main/scala/nutcore/mem/Cache.scala 321:18]
  wire  _cmd_T = state == 4'h1; // @[src/main/scala/nutcore/mem/Cache.scala 322:23]
  wire [2:0] _cmd_T_2 = writeBeatCnt_value == 3'h7 ? 3'h7 : 3'h3; // @[src/main/scala/nutcore/mem/Cache.scala 323:8]
  wire [2:0] cmd = state == 4'h1 ? 3'h2 : _cmd_T_2; // @[src/main/scala/nutcore/mem/Cache.scala 322:16]
  wire  _io_mem_req_valid_T_2 = state2 == 2'h2; // @[src/main/scala/nutcore/mem/Cache.scala 329:89]
  reg  afterFirstRead; // @[src/main/scala/nutcore/mem/Cache.scala 336:31]
  reg  alreadyOutFire; // @[src/main/scala/nutcore/mem/Cache.scala 337:33]
  wire  _GEN_12 = _T_5 | alreadyOutFire; // @[src/main/scala/nutcore/mem/Cache.scala 337:{33,33,33}]
  wire  _readingFirst_T_1 = io_mem_resp_ready & io_mem_resp_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  wire  _readingFirst_T_3 = state == 4'h2; // @[src/main/scala/nutcore/mem/Cache.scala 338:68]
  wire  readingFirst = ~afterFirstRead & _readingFirst_T_1 & state == 4'h2; // @[src/main/scala/nutcore/mem/Cache.scala 338:58]
  wire  _inRdataRegDemand_T_2 = mmio ? state == 4'h6 : readingFirst; // @[src/main/scala/nutcore/mem/Cache.scala 340:39]
  reg [63:0] inRdataRegDemand; // @[src/main/scala/nutcore/mem/Cache.scala 339:35]
  wire  _io_cohResp_valid_T = state == 4'h0; // @[src/main/scala/nutcore/mem/Cache.scala 343:31]
  wire  _io_cohResp_valid_T_4 = _T_15 & _io_mem_req_valid_T_2; // @[src/main/scala/nutcore/mem/Cache.scala 344:46]
  wire  _releaseLast_T_2 = _T_15 & io_cohResp_valid; // @[src/main/scala/nutcore/mem/Cache.scala 346:49]
  reg [2:0] releaseLast_c_value; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
  wire  releaseLast_wrap_wrap = releaseLast_c_value == 3'h7; // @[src/main/scala/chisel3/util/Counter.scala 73:24]
  wire [2:0] _releaseLast_wrap_value_T_1 = releaseLast_c_value + 3'h1; // @[src/main/scala/chisel3/util/Counter.scala 77:24]
  wire  releaseLast = _releaseLast_T_2 & releaseLast_wrap_wrap; // @[src/main/scala/chisel3/util/Counter.scala 118:{16,23} 117:24]
  wire [2:0] _io_cohResp_bits_cmd_T_1 = releaseLast ? 3'h6 : 3'h0; // @[src/main/scala/nutcore/mem/Cache.scala 347:54]
  wire [3:0] _io_cohResp_bits_cmd_T_2 = hit ? 4'hc : 4'h8; // @[src/main/scala/nutcore/mem/Cache.scala 348:8]
  wire  respToL1Fire = _T_29 & _io_mem_req_valid_T_2; // @[src/main/scala/nutcore/mem/Cache.scala 350:51]
  wire  _respToL1Last_T_6 = (_io_cohResp_valid_T | _io_cohResp_valid_T_4) & hitReadBurst & io_out_ready; // @[src/main/scala/nutcore/mem/Cache.scala 351:112]
  reg [2:0] respToL1Last_c_value; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
  wire  respToL1Last_wrap_wrap = respToL1Last_c_value == 3'h7; // @[src/main/scala/chisel3/util/Counter.scala 73:24]
  wire [2:0] _respToL1Last_wrap_value_T_1 = respToL1Last_c_value + 3'h1; // @[src/main/scala/chisel3/util/Counter.scala 77:24]
  wire  respToL1Last = _respToL1Last_T_6 & respToL1Last_wrap_wrap; // @[src/main/scala/chisel3/util/Counter.scala 118:{16,23} 117:24]
  wire [3:0] _state_T = hit ? 4'h8 : 4'h0; // @[src/main/scala/nutcore/mem/Cache.scala 360:23]
  wire [2:0] _value_T_4 = addr_wordIndex + 3'h1; // @[src/main/scala/nutcore/mem/Cache.scala 365:93]
  wire [2:0] _value_T_5 = addr_wordIndex == 3'h7 ? 3'h0 : _value_T_4; // @[src/main/scala/nutcore/mem/Cache.scala 365:33]
  wire [3:0] _state_T_3 = meta_dirty ? 4'h3 : 4'h1; // @[src/main/scala/nutcore/mem/Cache.scala 367:42]
  wire [3:0] _state_T_4 = mmio ? 4'h5 : _state_T_3; // @[src/main/scala/nutcore/mem/Cache.scala 367:21]
  wire [3:0] _GEN_20 = miss | mmio ? _state_T_4 : state; // @[src/main/scala/nutcore/mem/Cache.scala 366:49 367:15 294:22]
  wire  _T_41 = io_mmio_req_ready & io_mmio_req_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  wire  _T_43 = io_mmio_resp_ready & io_mmio_resp_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  wire [3:0] _GEN_26 = _T_43 ? 4'h7 : state; // @[src/main/scala/nutcore/mem/Cache.scala 294:22 372:{48,56}]
  wire [2:0] _value_T_7 = readBeatCnt_value + 3'h1; // @[src/main/scala/chisel3/util/Counter.scala 77:24]
  wire [2:0] _GEN_27 = io_cohResp_valid | respToL1Fire ? _value_T_7 : readBeatCnt_value; // @[src/main/scala/nutcore/mem/Cache.scala 375:46 src/main/scala/chisel3/util/Counter.scala 77:15 61:40]
  wire [3:0] _GEN_28 = probe & io_cohResp_valid & releaseLast | respToL1Fire & respToL1Last ? 4'h0 : state; // @[src/main/scala/nutcore/mem/Cache.scala 294:22 376:{86,94}]
  wire [3:0] _GEN_29 = _T_26 ? 4'h2 : state; // @[src/main/scala/nutcore/mem/Cache.scala 379:48 380:13 294:22]
  wire [2:0] _GEN_30 = _T_26 ? addr_wordIndex : readBeatCnt_value; // @[src/main/scala/nutcore/mem/Cache.scala 379:48 381:25 src/main/scala/chisel3/util/Counter.scala 61:40]
  wire [2:0] _GEN_31 = _T_6 ? 3'h0 : _GEN_0; // @[src/main/scala/nutcore/mem/Cache.scala 388:{52,75}]
  wire  _T_57 = io_mem_resp_bits_cmd == 4'h6; // @[src/main/scala/bus/simplebus/SimpleBus.scala 91:24]
  wire [3:0] _GEN_32 = _T_57 ? 4'h7 : state; // @[src/main/scala/nutcore/mem/Cache.scala 294:22 389:{44,52}]
  wire  _GEN_33 = _readingFirst_T_1 | afterFirstRead; // @[src/main/scala/nutcore/mem/Cache.scala 385:31 386:24 336:31]
  wire [2:0] _GEN_34 = _readingFirst_T_1 ? _value_T_7 : readBeatCnt_value; // @[src/main/scala/nutcore/mem/Cache.scala 385:31 src/main/scala/chisel3/util/Counter.scala 77:15 61:40]
  wire [2:0] _GEN_35 = _readingFirst_T_1 ? _GEN_31 : _GEN_0; // @[src/main/scala/nutcore/mem/Cache.scala 385:31]
  wire [3:0] _GEN_36 = _readingFirst_T_1 ? _GEN_32 : state; // @[src/main/scala/nutcore/mem/Cache.scala 294:22 385:31]
  wire [2:0] _value_T_11 = writeBeatCnt_value + 3'h1; // @[src/main/scala/chisel3/util/Counter.scala 77:24]
  wire [2:0] _GEN_37 = _T_26 ? _value_T_11 : writeBeatCnt_value; // @[src/main/scala/nutcore/mem/Cache.scala 394:30 src/main/scala/chisel3/util/Counter.scala 77:15 61:40]
  wire  _T_60 = io_mem_req_bits_cmd == 4'h7; // @[src/main/scala/bus/simplebus/SimpleBus.scala 78:27]
  wire [3:0] _GEN_38 = _T_60 & _T_26 ? 4'h4 : state; // @[src/main/scala/nutcore/mem/Cache.scala 294:22 395:{63,71}]
  wire [3:0] _GEN_39 = _readingFirst_T_1 ? 4'h1 : state; // @[src/main/scala/nutcore/mem/Cache.scala 294:22 398:{51,59}]
  wire [3:0] _GEN_40 = _GEN_12 ? 4'h0 : state; // @[src/main/scala/nutcore/mem/Cache.scala 294:22 399:{74,82}]
  wire [3:0] _GEN_41 = 4'h7 == state ? _GEN_40 : state; // @[src/main/scala/nutcore/mem/Cache.scala 353:18 294:22]
  wire [3:0] _GEN_42 = 4'h4 == state ? _GEN_39 : _GEN_41; // @[src/main/scala/nutcore/mem/Cache.scala 353:18]
  wire [2:0] _GEN_43 = 4'h3 == state ? _GEN_37 : writeBeatCnt_value; // @[src/main/scala/nutcore/mem/Cache.scala 353:18 src/main/scala/chisel3/util/Counter.scala 61:40]
  wire [3:0] _GEN_44 = 4'h3 == state ? _GEN_38 : _GEN_42; // @[src/main/scala/nutcore/mem/Cache.scala 353:18]
  wire  _GEN_45 = 4'h2 == state ? _GEN_33 : afterFirstRead; // @[src/main/scala/nutcore/mem/Cache.scala 353:18 336:31]
  wire [2:0] _GEN_46 = 4'h2 == state ? _GEN_34 : readBeatCnt_value; // @[src/main/scala/nutcore/mem/Cache.scala 353:18 src/main/scala/chisel3/util/Counter.scala 61:40]
  wire [2:0] _GEN_47 = 4'h2 == state ? _GEN_35 : _GEN_0; // @[src/main/scala/nutcore/mem/Cache.scala 353:18]
  wire [3:0] _GEN_48 = 4'h2 == state ? _GEN_36 : _GEN_44; // @[src/main/scala/nutcore/mem/Cache.scala 353:18]
  wire [2:0] _GEN_49 = 4'h2 == state ? writeBeatCnt_value : _GEN_43; // @[src/main/scala/nutcore/mem/Cache.scala 353:18 src/main/scala/chisel3/util/Counter.scala 61:40]
  wire [3:0] _GEN_50 = 4'h1 == state ? _GEN_29 : _GEN_48; // @[src/main/scala/nutcore/mem/Cache.scala 353:18]
  wire [2:0] _GEN_51 = 4'h1 == state ? _GEN_30 : _GEN_46; // @[src/main/scala/nutcore/mem/Cache.scala 353:18]
  wire  _GEN_52 = 4'h1 == state ? afterFirstRead : _GEN_45; // @[src/main/scala/nutcore/mem/Cache.scala 353:18 336:31]
  wire [2:0] _GEN_53 = 4'h1 == state ? _GEN_0 : _GEN_47; // @[src/main/scala/nutcore/mem/Cache.scala 353:18]
  wire [2:0] _GEN_54 = 4'h1 == state ? writeBeatCnt_value : _GEN_49; // @[src/main/scala/nutcore/mem/Cache.scala 353:18 src/main/scala/chisel3/util/Counter.scala 61:40]
  wire [2:0] _GEN_55 = 4'h8 == state ? _GEN_27 : _GEN_51; // @[src/main/scala/nutcore/mem/Cache.scala 353:18]
  wire [3:0] _GEN_56 = 4'h8 == state ? _GEN_28 : _GEN_50; // @[src/main/scala/nutcore/mem/Cache.scala 353:18]
  wire  _GEN_57 = 4'h8 == state ? afterFirstRead : _GEN_52; // @[src/main/scala/nutcore/mem/Cache.scala 353:18 336:31]
  wire [2:0] _GEN_58 = 4'h8 == state ? _GEN_0 : _GEN_53; // @[src/main/scala/nutcore/mem/Cache.scala 353:18]
  wire [2:0] _GEN_59 = 4'h8 == state ? writeBeatCnt_value : _GEN_54; // @[src/main/scala/nutcore/mem/Cache.scala 353:18 src/main/scala/chisel3/util/Counter.scala 61:40]
  wire [63:0] _dataRefill_T = readingFirst ? wordMask : 64'h0; // @[src/main/scala/nutcore/mem/Cache.scala 402:67]
  wire [63:0] _dataRefill_T_1 = io_in_bits_req_wdata & _dataRefill_T; // @[src/main/scala/utils/BitUtils.scala 34:14]
  wire [63:0] _dataRefill_T_2 = ~_dataRefill_T; // @[src/main/scala/utils/BitUtils.scala 34:39]
  wire [63:0] _dataRefill_T_3 = io_mem_resp_bits_rdata & _dataRefill_T_2; // @[src/main/scala/utils/BitUtils.scala 34:37]
  wire  dataRefillWriteBus_x9 = _readingFirst_T_3 & _readingFirst_T_1; // @[src/main/scala/nutcore/mem/Cache.scala 404:39]
  wire  metaRefillWriteBus_req_valid = dataRefillWriteBus_x9 & _T_57; // @[src/main/scala/nutcore/mem/Cache.scala 412:59]
  wire  _io_out_bits_cmd_T_4 = ~io_in_bits_req_cmd[0] & ~io_in_bits_req_cmd[3]; // @[src/main/scala/bus/simplebus/SimpleBus.scala 73:26]
  wire [2:0] _io_out_bits_cmd_T_6 = io_in_bits_req_cmd[0] ? 3'h5 : 3'h0; // @[src/main/scala/nutcore/mem/Cache.scala 440:79]
  wire [2:0] _io_out_bits_cmd_T_7 = _io_out_bits_cmd_T_4 ? 3'h6 : _io_out_bits_cmd_T_6; // @[src/main/scala/nutcore/mem/Cache.scala 440:27]
  wire  _io_out_valid_T_4 = state == 4'h7; // @[src/main/scala/nutcore/mem/Cache.scala 446:48]
  wire  _io_out_valid_T_23 = io_in_bits_req_cmd[0] | mmio ? _io_out_valid_T_4 : afterFirstRead & ~alreadyOutFire; // @[src/main/scala/nutcore/mem/Cache.scala 447:45]
  wire  _io_out_valid_T_25 = probe ? 1'h0 : hit | _io_out_valid_T_23; // @[src/main/scala/nutcore/mem/Cache.scala 447:8]
  wire  _io_isFinish_T_4 = miss ? _io_cohResp_valid_T : _T_15 & releaseLast; // @[src/main/scala/nutcore/mem/Cache.scala 454:51]
  wire  _io_isFinish_T_13 = hit | io_in_bits_req_cmd[0] ? _T_5 : _io_out_valid_T_4 & _GEN_12; // @[src/main/scala/nutcore/mem/Cache.scala 455:8]
  wire [255:0] _T_89 = {io_in_bits_datas_3_data,io_in_bits_datas_2_data,io_in_bits_datas_1_data,io_in_bits_datas_0_data}
    ; // @[src/main/scala/nutcore/mem/Cache.scala 464:465]
  reg [63:0] c; // @[src/main/scala/utils/GTimer.scala 24:20]
  wire [63:0] _c_T_1 = c + 64'h1; // @[src/main/scala/utils/GTimer.scala 25:12]
  reg [63:0] c_1; // @[src/main/scala/utils/GTimer.scala 24:20]
  wire [63:0] _c_T_3 = c_1 + 64'h1; // @[src/main/scala/utils/GTimer.scala 25:12]
  reg [63:0] c_2; // @[src/main/scala/utils/GTimer.scala 24:20]
  wire [63:0] _c_T_5 = c_2 + 64'h1; // @[src/main/scala/utils/GTimer.scala 25:12]
  wire  _T_96 = io_metaWriteBus_req_valid & DISPLAY_ENABLE; // @[src/main/scala/utils/Debug.scala 55:16]
  reg [63:0] c_3; // @[src/main/scala/utils/GTimer.scala 24:20]
  wire [63:0] _c_T_7 = c_3 + 64'h1; // @[src/main/scala/utils/GTimer.scala 25:12]
  reg [63:0] c_4; // @[src/main/scala/utils/GTimer.scala 24:20]
  wire [63:0] _c_T_9 = c_4 + 64'h1; // @[src/main/scala/utils/GTimer.scala 25:12]
  reg [63:0] c_5; // @[src/main/scala/utils/GTimer.scala 24:20]
  wire [63:0] _c_T_11 = c_5 + 64'h1; // @[src/main/scala/utils/GTimer.scala 25:12]
  reg [63:0] c_6; // @[src/main/scala/utils/GTimer.scala 24:20]
  wire [63:0] _c_T_13 = c_6 + 64'h1; // @[src/main/scala/utils/GTimer.scala 25:12]
  reg [63:0] c_7; // @[src/main/scala/utils/GTimer.scala 24:20]
  wire [63:0] _c_T_15 = c_7 + 64'h1; // @[src/main/scala/utils/GTimer.scala 25:12]
  reg [63:0] c_8; // @[src/main/scala/utils/GTimer.scala 24:20]
  wire [63:0] _c_T_17 = c_8 + 64'h1; // @[src/main/scala/utils/GTimer.scala 25:12]
  wire  _T_128 = io_dataWriteBus_req_valid & DISPLAY_ENABLE; // @[src/main/scala/utils/Debug.scala 55:16]
  wire  _T_135 = _T_14 & _T_26; // @[src/main/scala/nutcore/mem/Cache.scala 473:35]
  reg [63:0] c_9; // @[src/main/scala/utils/GTimer.scala 24:20]
  wire [63:0] _c_T_19 = c_9 + 64'h1; // @[src/main/scala/utils/GTimer.scala 25:12]
  wire  _T_140 = _T_135 & DISPLAY_ENABLE; // @[src/main/scala/utils/Debug.scala 55:16]
  wire  _T_147 = _cmd_T & _T_26; // @[src/main/scala/nutcore/mem/Cache.scala 474:34]
  reg [63:0] c_10; // @[src/main/scala/utils/GTimer.scala 24:20]
  wire [63:0] _c_T_21 = c_10 + 64'h1; // @[src/main/scala/utils/GTimer.scala 25:12]
  wire  _T_152 = _T_147 & DISPLAY_ENABLE; // @[src/main/scala/utils/Debug.scala 55:16]
  reg [63:0] c_11; // @[src/main/scala/utils/GTimer.scala 24:20]
  wire [63:0] _c_T_23 = c_11 + 64'h1; // @[src/main/scala/utils/GTimer.scala 25:12]
  wire  _T_164 = dataRefillWriteBus_x9 & DISPLAY_ENABLE; // @[src/main/scala/utils/Debug.scala 55:16]
  wire  _WIRE = mmio; // @[src/main/scala/nutcore/mem/Cache.scala 259:26]
  Arbiter metaWriteArb ( // @[src/main/scala/nutcore/mem/Cache.scala 254:28]
    .io_in_0_valid(metaWriteArb_io_in_0_valid),
    .io_in_0_bits_setIdx(metaWriteArb_io_in_0_bits_setIdx),
    .io_in_0_bits_data_tag(metaWriteArb_io_in_0_bits_data_tag),
    .io_in_0_bits_data_dirty(metaWriteArb_io_in_0_bits_data_dirty),
    .io_in_0_bits_waymask(metaWriteArb_io_in_0_bits_waymask),
    .io_in_1_valid(metaWriteArb_io_in_1_valid),
    .io_in_1_bits_setIdx(metaWriteArb_io_in_1_bits_setIdx),
    .io_in_1_bits_data_tag(metaWriteArb_io_in_1_bits_data_tag),
    .io_in_1_bits_data_dirty(metaWriteArb_io_in_1_bits_data_dirty),
    .io_in_1_bits_waymask(metaWriteArb_io_in_1_bits_waymask),
    .io_out_valid(metaWriteArb_io_out_valid),
    .io_out_bits_setIdx(metaWriteArb_io_out_bits_setIdx),
    .io_out_bits_data_tag(metaWriteArb_io_out_bits_data_tag),
    .io_out_bits_data_dirty(metaWriteArb_io_out_bits_data_dirty),
    .io_out_bits_waymask(metaWriteArb_io_out_bits_waymask)
  );
  Arbiter_1 dataWriteArb ( // @[src/main/scala/nutcore/mem/Cache.scala 255:28]
    .io_in_0_valid(dataWriteArb_io_in_0_valid),
    .io_in_0_bits_setIdx(dataWriteArb_io_in_0_bits_setIdx),
    .io_in_0_bits_data_data(dataWriteArb_io_in_0_bits_data_data),
    .io_in_0_bits_waymask(dataWriteArb_io_in_0_bits_waymask),
    .io_in_1_valid(dataWriteArb_io_in_1_valid),
    .io_in_1_bits_setIdx(dataWriteArb_io_in_1_bits_setIdx),
    .io_in_1_bits_data_data(dataWriteArb_io_in_1_bits_data_data),
    .io_in_1_bits_waymask(dataWriteArb_io_in_1_bits_waymask),
    .io_out_valid(dataWriteArb_io_out_valid),
    .io_out_bits_setIdx(dataWriteArb_io_out_bits_setIdx),
    .io_out_bits_data_data(dataWriteArb_io_out_bits_data_data),
    .io_out_bits_waymask(dataWriteArb_io_out_bits_waymask)
  );
  assign io_in_ready = io_out_ready & (_io_cohResp_valid_T & ~hitReadBurst) & ~miss & ~probe; // @[src/main/scala/nutcore/mem/Cache.scala 458:79]
  assign io_out_valid = io_in_valid & _io_out_valid_T_25; // @[src/main/scala/nutcore/mem/Cache.scala 445:31]
  assign io_out_bits_cmd = {{1'd0}, _io_out_bits_cmd_T_7}; // @[src/main/scala/nutcore/mem/Cache.scala 440:21]
  assign io_out_bits_rdata = hit ? dataRead : inRdataRegDemand; // @[src/main/scala/nutcore/mem/Cache.scala 439:29]
  assign io_isFinish = probe ? io_cohResp_valid & _io_isFinish_T_4 : _io_isFinish_T_13; // @[src/main/scala/nutcore/mem/Cache.scala 454:21]
  assign io_dataReadBus_req_valid = (state == 4'h3 | state == 4'h8) & state2 == 2'h0; // @[src/main/scala/nutcore/mem/Cache.scala 306:81]
  assign io_dataReadBus_req_bits_setIdx = {addr_index,_T_20}; // @[src/main/scala/nutcore/mem/Cache.scala 307:17]
  assign io_dataWriteBus_req_valid = dataWriteArb_io_out_valid; // @[src/main/scala/nutcore/mem/Cache.scala 409:23]
  assign io_dataWriteBus_req_bits_setIdx = dataWriteArb_io_out_bits_setIdx; // @[src/main/scala/nutcore/mem/Cache.scala 409:23]
  assign io_dataWriteBus_req_bits_data_data = dataWriteArb_io_out_bits_data_data; // @[src/main/scala/nutcore/mem/Cache.scala 409:23]
  assign io_dataWriteBus_req_bits_waymask = dataWriteArb_io_out_bits_waymask; // @[src/main/scala/nutcore/mem/Cache.scala 409:23]
  assign io_metaWriteBus_req_valid = metaWriteArb_io_out_valid; // @[src/main/scala/nutcore/mem/Cache.scala 419:23]
  assign io_metaWriteBus_req_bits_setIdx = metaWriteArb_io_out_bits_setIdx; // @[src/main/scala/nutcore/mem/Cache.scala 419:23]
  assign io_metaWriteBus_req_bits_data_tag = metaWriteArb_io_out_bits_data_tag; // @[src/main/scala/nutcore/mem/Cache.scala 419:23]
  assign io_metaWriteBus_req_bits_data_valid = 1'h1; // @[src/main/scala/nutcore/mem/Cache.scala 419:23]
  assign io_metaWriteBus_req_bits_data_dirty = metaWriteArb_io_out_bits_data_dirty; // @[src/main/scala/nutcore/mem/Cache.scala 419:23]
  assign io_metaWriteBus_req_bits_waymask = metaWriteArb_io_out_bits_waymask; // @[src/main/scala/nutcore/mem/Cache.scala 419:23]
  assign io_mem_req_valid = _cmd_T | _T_14 & state2 == 2'h2; // @[src/main/scala/nutcore/mem/Cache.scala 329:48]
  assign io_mem_req_bits_addr = _cmd_T ? raddr : waddr; // @[src/main/scala/nutcore/mem/Cache.scala 324:35]
  assign io_mem_req_bits_size = 3'h3; // @[src/main/scala/bus/simplebus/SimpleBus.scala 66:15]
  assign io_mem_req_bits_cmd = {{1'd0}, cmd}; // @[src/main/scala/bus/simplebus/SimpleBus.scala 65:14]
  assign io_mem_req_bits_wmask = 8'hff; // @[src/main/scala/nutcore/mem/Cache.scala 326:37]
  assign io_mem_req_bits_wdata = _dataHitWay_T_9 | _dataHitWay_T_7; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign io_mem_resp_ready = 1'h1; // @[src/main/scala/nutcore/mem/Cache.scala 328:21]
  assign io_mmio_req_valid = state == 4'h5; // @[src/main/scala/nutcore/mem/Cache.scala 334:31]
  assign io_mmio_req_bits_addr = io_in_bits_req_addr; // @[src/main/scala/nutcore/mem/Cache.scala 332:20]
  assign io_mmio_req_bits_size = io_in_bits_req_size; // @[src/main/scala/nutcore/mem/Cache.scala 332:20]
  assign io_mmio_req_bits_cmd = io_in_bits_req_cmd; // @[src/main/scala/nutcore/mem/Cache.scala 332:20]
  assign io_mmio_req_bits_wmask = io_in_bits_req_wmask; // @[src/main/scala/nutcore/mem/Cache.scala 332:20]
  assign io_mmio_req_bits_wdata = io_in_bits_req_wdata; // @[src/main/scala/nutcore/mem/Cache.scala 332:20]
  assign io_mmio_resp_ready = 1'h1; // @[src/main/scala/nutcore/mem/Cache.scala 333:22]
  assign io_cohResp_valid = state == 4'h0 & probe | _io_cohResp_valid_T_4; // @[src/main/scala/nutcore/mem/Cache.scala 343:53]
  assign io_cohResp_bits_cmd = _T_15 ? {{1'd0}, _io_cohResp_bits_cmd_T_1} : _io_cohResp_bits_cmd_T_2; // @[src/main/scala/nutcore/mem/Cache.scala 347:29]
  assign io_cohResp_bits_rdata = _dataHitWay_T_9 | _dataHitWay_T_7; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign io_dataReadRespToL1 = hitReadBurst & (_io_cohResp_valid_T & io_out_ready | _io_cohResp_valid_T_4); // @[src/main/scala/nutcore/mem/Cache.scala 459:39]
  assign _WIRE_19 = _WIRE;
  assign metaWriteArb_io_in_0_valid = hitWrite & ~meta_dirty; // @[src/main/scala/nutcore/mem/Cache.scala 289:22]
  assign metaWriteArb_io_in_0_bits_setIdx = io_in_bits_req_addr[12:6]; // @[src/main/scala/nutcore/mem/Cache.scala 77:45]
  assign metaWriteArb_io_in_0_bits_data_tag = _meta_T_23 | _meta_T_21; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign metaWriteArb_io_in_0_bits_data_dirty = 1'h1; // @[src/main/scala/nutcore/mem/Cache.scala 290:16 95:16]
  assign metaWriteArb_io_in_0_bits_waymask = io_in_bits_waymask; // @[src/main/scala/nutcore/mem/Cache.scala 288:29 src/main/scala/utils/SRAMTemplate.scala 38:24]
  assign metaWriteArb_io_in_1_valid = dataRefillWriteBus_x9 & _T_57; // @[src/main/scala/nutcore/mem/Cache.scala 412:59]
  assign metaWriteArb_io_in_1_bits_setIdx = io_in_bits_req_addr[12:6]; // @[src/main/scala/nutcore/mem/Cache.scala 77:45]
  assign metaWriteArb_io_in_1_bits_data_tag = io_in_bits_req_addr[31:13]; // @[src/main/scala/nutcore/mem/Cache.scala 258:31]
  assign metaWriteArb_io_in_1_bits_data_dirty = io_in_bits_req_cmd[0]; // @[src/main/scala/bus/simplebus/SimpleBus.scala 74:22]
  assign metaWriteArb_io_in_1_bits_waymask = io_in_bits_waymask; // @[src/main/scala/nutcore/mem/Cache.scala 411:32 src/main/scala/utils/SRAMTemplate.scala 38:24]
  assign dataWriteArb_io_in_0_valid = hit & io_in_bits_req_cmd[0]; // @[src/main/scala/nutcore/mem/Cache.scala 283:22]
  assign dataWriteArb_io_in_0_bits_setIdx = {addr_index,_dataHitWriteBus_x3_T_3}; // @[src/main/scala/nutcore/mem/Cache.scala 286:35]
  assign dataWriteArb_io_in_0_bits_data_data = _dataHitWriteBus_x1_T | _dataHitWriteBus_x1_T_2; // @[src/main/scala/utils/BitUtils.scala 34:26]
  assign dataWriteArb_io_in_0_bits_waymask = io_in_bits_waymask; // @[src/main/scala/nutcore/mem/Cache.scala 284:29 src/main/scala/utils/SRAMTemplate.scala 38:24]
  assign dataWriteArb_io_in_1_valid = _readingFirst_T_3 & _readingFirst_T_1; // @[src/main/scala/nutcore/mem/Cache.scala 404:39]
  assign dataWriteArb_io_in_1_bits_setIdx = {addr_index,readBeatCnt_value}; // @[src/main/scala/nutcore/mem/Cache.scala 404:72]
  assign dataWriteArb_io_in_1_bits_data_data = _dataRefill_T_1 | _dataRefill_T_3; // @[src/main/scala/utils/BitUtils.scala 34:26]
  assign dataWriteArb_io_in_1_bits_waymask = io_in_bits_waymask; // @[src/main/scala/nutcore/mem/Cache.scala 403:32 src/main/scala/utils/SRAMTemplate.scala 38:24]
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/chisel3/util/Counter.scala 61:40]
      writeL2BeatCnt_value <= 3'h0; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end else if (4'h0 == state) begin // @[src/main/scala/nutcore/mem/Cache.scala 353:18]
      writeL2BeatCnt_value <= _GEN_0;
    end else if (4'h5 == state) begin // @[src/main/scala/nutcore/mem/Cache.scala 353:18]
      writeL2BeatCnt_value <= _GEN_0;
    end else if (4'h6 == state) begin // @[src/main/scala/nutcore/mem/Cache.scala 353:18]
      writeL2BeatCnt_value <= _GEN_0;
    end else begin
      writeL2BeatCnt_value <= _GEN_58;
    end
    if (reset) begin // @[src/main/scala/nutcore/mem/Cache.scala 294:22]
      state <= 4'h0; // @[src/main/scala/nutcore/mem/Cache.scala 294:22]
    end else if (4'h0 == state) begin // @[src/main/scala/nutcore/mem/Cache.scala 353:18]
      if (probe) begin // @[src/main/scala/nutcore/mem/Cache.scala 358:20]
        if (io_cohResp_valid) begin // @[src/main/scala/nutcore/mem/Cache.scala 359:32]
          state <= _state_T; // @[src/main/scala/nutcore/mem/Cache.scala 360:17]
        end
      end else if (_T_29) begin // @[src/main/scala/nutcore/mem/Cache.scala 363:50]
        state <= 4'h8; // @[src/main/scala/nutcore/mem/Cache.scala 364:15]
      end else begin
        state <= _GEN_20;
      end
    end else if (4'h5 == state) begin // @[src/main/scala/nutcore/mem/Cache.scala 353:18]
      if (_T_41) begin // @[src/main/scala/nutcore/mem/Cache.scala 371:46]
        state <= 4'h6; // @[src/main/scala/nutcore/mem/Cache.scala 371:54]
      end
    end else if (4'h6 == state) begin // @[src/main/scala/nutcore/mem/Cache.scala 353:18]
      state <= _GEN_26;
    end else begin
      state <= _GEN_56;
    end
    if (reset) begin // @[src/main/scala/chisel3/util/Counter.scala 61:40]
      readBeatCnt_value <= 3'h0; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end else if (4'h0 == state) begin // @[src/main/scala/nutcore/mem/Cache.scala 353:18]
      if (probe) begin // @[src/main/scala/nutcore/mem/Cache.scala 358:20]
        if (io_cohResp_valid) begin // @[src/main/scala/nutcore/mem/Cache.scala 359:32]
          readBeatCnt_value <= addr_wordIndex; // @[src/main/scala/nutcore/mem/Cache.scala 361:29]
        end
      end else if (_T_29) begin // @[src/main/scala/nutcore/mem/Cache.scala 363:50]
        readBeatCnt_value <= _value_T_5; // @[src/main/scala/nutcore/mem/Cache.scala 365:27]
      end
    end else if (!(4'h5 == state)) begin // @[src/main/scala/nutcore/mem/Cache.scala 353:18]
      if (!(4'h6 == state)) begin // @[src/main/scala/nutcore/mem/Cache.scala 353:18]
        readBeatCnt_value <= _GEN_55;
      end
    end
    if (reset) begin // @[src/main/scala/chisel3/util/Counter.scala 61:40]
      writeBeatCnt_value <= 3'h0; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end else if (!(4'h0 == state)) begin // @[src/main/scala/nutcore/mem/Cache.scala 353:18]
      if (!(4'h5 == state)) begin // @[src/main/scala/nutcore/mem/Cache.scala 353:18]
        if (!(4'h6 == state)) begin // @[src/main/scala/nutcore/mem/Cache.scala 353:18]
          writeBeatCnt_value <= _GEN_59;
        end
      end
    end
    if (reset) begin // @[src/main/scala/nutcore/mem/Cache.scala 304:23]
      state2 <= 2'h0; // @[src/main/scala/nutcore/mem/Cache.scala 304:23]
    end else if (2'h0 == state2) begin // @[src/main/scala/nutcore/mem/Cache.scala 311:19]
      if (_T_23) begin // @[src/main/scala/nutcore/mem/Cache.scala 312:51]
        state2 <= 2'h1; // @[src/main/scala/nutcore/mem/Cache.scala 312:60]
      end
    end else if (2'h1 == state2) begin // @[src/main/scala/nutcore/mem/Cache.scala 311:19]
      state2 <= 2'h2; // @[src/main/scala/nutcore/mem/Cache.scala 313:35]
    end else if (2'h2 == state2) begin // @[src/main/scala/nutcore/mem/Cache.scala 311:19]
      state2 <= _GEN_8;
    end
    if (state2 == 2'h1) begin // @[src/main/scala/nutcore/mem/Cache.scala 308:26]
      dataWay_0_data <= io_dataReadBus_resp_data_0_data; // @[src/main/scala/nutcore/mem/Cache.scala 308:26]
    end
    if (state2 == 2'h1) begin // @[src/main/scala/nutcore/mem/Cache.scala 308:26]
      dataWay_1_data <= io_dataReadBus_resp_data_1_data; // @[src/main/scala/nutcore/mem/Cache.scala 308:26]
    end
    if (state2 == 2'h1) begin // @[src/main/scala/nutcore/mem/Cache.scala 308:26]
      dataWay_2_data <= io_dataReadBus_resp_data_2_data; // @[src/main/scala/nutcore/mem/Cache.scala 308:26]
    end
    if (state2 == 2'h1) begin // @[src/main/scala/nutcore/mem/Cache.scala 308:26]
      dataWay_3_data <= io_dataReadBus_resp_data_3_data; // @[src/main/scala/nutcore/mem/Cache.scala 308:26]
    end
    if (reset) begin // @[src/main/scala/nutcore/mem/Cache.scala 336:31]
      afterFirstRead <= 1'h0; // @[src/main/scala/nutcore/mem/Cache.scala 336:31]
    end else if (4'h0 == state) begin // @[src/main/scala/nutcore/mem/Cache.scala 353:18]
      afterFirstRead <= 1'h0; // @[src/main/scala/nutcore/mem/Cache.scala 355:22]
    end else if (!(4'h5 == state)) begin // @[src/main/scala/nutcore/mem/Cache.scala 353:18]
      if (!(4'h6 == state)) begin // @[src/main/scala/nutcore/mem/Cache.scala 353:18]
        afterFirstRead <= _GEN_57;
      end
    end
    if (reset) begin // @[src/main/scala/nutcore/mem/Cache.scala 337:33]
      alreadyOutFire <= 1'h0; // @[src/main/scala/nutcore/mem/Cache.scala 337:33]
    end else if (4'h0 == state) begin // @[src/main/scala/nutcore/mem/Cache.scala 353:18]
      alreadyOutFire <= 1'h0; // @[src/main/scala/nutcore/mem/Cache.scala 356:22]
    end else begin
      alreadyOutFire <= _GEN_12;
    end
    if (_inRdataRegDemand_T_2) begin // @[src/main/scala/nutcore/mem/Cache.scala 339:35]
      if (mmio) begin // @[src/main/scala/nutcore/mem/Cache.scala 339:39]
        inRdataRegDemand <= io_mmio_resp_bits_rdata;
      end else begin
        inRdataRegDemand <= io_mem_resp_bits_rdata;
      end
    end
    if (reset) begin // @[src/main/scala/chisel3/util/Counter.scala 61:40]
      releaseLast_c_value <= 3'h0; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end else if (_releaseLast_T_2) begin // @[src/main/scala/chisel3/util/Counter.scala 118:16]
      releaseLast_c_value <= _releaseLast_wrap_value_T_1; // @[src/main/scala/chisel3/util/Counter.scala 77:15]
    end
    if (reset) begin // @[src/main/scala/chisel3/util/Counter.scala 61:40]
      respToL1Last_c_value <= 3'h0; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end else if (_respToL1Last_T_6) begin // @[src/main/scala/chisel3/util/Counter.scala 118:16]
      respToL1Last_c_value <= _respToL1Last_wrap_value_T_1; // @[src/main/scala/chisel3/util/Counter.scala 77:15]
    end
    if (reset) begin // @[src/main/scala/utils/GTimer.scala 24:20]
      c <= 64'h0; // @[src/main/scala/utils/GTimer.scala 24:20]
    end else begin
      c <= _c_T_1; // @[src/main/scala/utils/GTimer.scala 25:7]
    end
    if (reset) begin // @[src/main/scala/utils/GTimer.scala 24:20]
      c_1 <= 64'h0; // @[src/main/scala/utils/GTimer.scala 24:20]
    end else begin
      c_1 <= _c_T_3; // @[src/main/scala/utils/GTimer.scala 25:7]
    end
    if (reset) begin // @[src/main/scala/utils/GTimer.scala 24:20]
      c_2 <= 64'h0; // @[src/main/scala/utils/GTimer.scala 24:20]
    end else begin
      c_2 <= _c_T_5; // @[src/main/scala/utils/GTimer.scala 25:7]
    end
    if (reset) begin // @[src/main/scala/utils/GTimer.scala 24:20]
      c_3 <= 64'h0; // @[src/main/scala/utils/GTimer.scala 24:20]
    end else begin
      c_3 <= _c_T_7; // @[src/main/scala/utils/GTimer.scala 25:7]
    end
    if (reset) begin // @[src/main/scala/utils/GTimer.scala 24:20]
      c_4 <= 64'h0; // @[src/main/scala/utils/GTimer.scala 24:20]
    end else begin
      c_4 <= _c_T_9; // @[src/main/scala/utils/GTimer.scala 25:7]
    end
    if (reset) begin // @[src/main/scala/utils/GTimer.scala 24:20]
      c_5 <= 64'h0; // @[src/main/scala/utils/GTimer.scala 24:20]
    end else begin
      c_5 <= _c_T_11; // @[src/main/scala/utils/GTimer.scala 25:7]
    end
    if (reset) begin // @[src/main/scala/utils/GTimer.scala 24:20]
      c_6 <= 64'h0; // @[src/main/scala/utils/GTimer.scala 24:20]
    end else begin
      c_6 <= _c_T_13; // @[src/main/scala/utils/GTimer.scala 25:7]
    end
    if (reset) begin // @[src/main/scala/utils/GTimer.scala 24:20]
      c_7 <= 64'h0; // @[src/main/scala/utils/GTimer.scala 24:20]
    end else begin
      c_7 <= _c_T_15; // @[src/main/scala/utils/GTimer.scala 25:7]
    end
    if (reset) begin // @[src/main/scala/utils/GTimer.scala 24:20]
      c_8 <= 64'h0; // @[src/main/scala/utils/GTimer.scala 24:20]
    end else begin
      c_8 <= _c_T_17; // @[src/main/scala/utils/GTimer.scala 25:7]
    end
    if (reset) begin // @[src/main/scala/utils/GTimer.scala 24:20]
      c_9 <= 64'h0; // @[src/main/scala/utils/GTimer.scala 24:20]
    end else begin
      c_9 <= _c_T_19; // @[src/main/scala/utils/GTimer.scala 25:7]
    end
    if (reset) begin // @[src/main/scala/utils/GTimer.scala 24:20]
      c_10 <= 64'h0; // @[src/main/scala/utils/GTimer.scala 24:20]
    end else begin
      c_10 <= _c_T_21; // @[src/main/scala/utils/GTimer.scala 25:7]
    end
    if (reset) begin // @[src/main/scala/utils/GTimer.scala 24:20]
      c_11 <= 64'h0; // @[src/main/scala/utils/GTimer.scala 24:20]
    end else begin
      c_11 <= _c_T_23; // @[src/main/scala/utils/GTimer.scala 25:7]
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~(mmio & hit))) begin
          $fwrite(32'h80000002,
            "Assertion failed: MMIO request should not hit in cache\n    at Cache.scala:265 assert(!(mmio && hit), \"MMIO request should not hit in cache\")\n"
            ); // @[src/main/scala/nutcore/mem/Cache.scala 265:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~(mmio & hit)) & ~reset) begin
          $fatal; // @[src/main/scala/nutcore/mem/Cache.scala 265:9]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3 & ~(~(metaHitWriteBus_x5 & metaRefillWriteBus_req_valid))) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Cache.scala:461 assert(!(metaHitWriteBus.req.valid && metaRefillWriteBus.req.valid))\n"
            ); // @[src/main/scala/nutcore/mem/Cache.scala 461:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~(metaHitWriteBus_x5 & metaRefillWriteBus_req_valid)) & _T_3) begin
          $fatal; // @[src/main/scala/nutcore/mem/Cache.scala 461:9]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3 & ~(~(hitWrite & dataRefillWriteBus_x9))) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Cache.scala:462 assert(!(dataHitWriteBus.req.valid && dataRefillWriteBus.req.valid))\n"
            ); // @[src/main/scala/nutcore/mem/Cache.scala 462:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~(hitWrite & dataRefillWriteBus_x9)) & _T_3) begin
          $fatal; // @[src/main/scala/nutcore/mem/Cache.scala 462:9]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_3) begin
          $fwrite(32'h80000002,"[%d] CacheStage3_1: ",c); // @[src/main/scala/utils/Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_3) begin
          $fwrite(32'h80000002," metaread idx %x waymask %b metas %x%x:%x %x%x:%x %x%x:%x %x%x:%x %x\n",addr_index,
            io_in_bits_waymask,io_in_bits_metas_0_valid,io_in_bits_metas_0_dirty,io_in_bits_metas_0_tag,
            io_in_bits_metas_1_valid,io_in_bits_metas_1_dirty,io_in_bits_metas_1_tag,io_in_bits_metas_2_valid,
            io_in_bits_metas_2_dirty,io_in_bits_metas_2_tag,io_in_bits_metas_3_valid,io_in_bits_metas_3_dirty,
            io_in_bits_metas_3_tag,_T_89); // @[src/main/scala/utils/Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_96 & _T_3) begin
          $fwrite(32'h80000002,"[%d] CacheStage3_1: ",c_2); // @[src/main/scala/utils/Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_96 & _T_3) begin
          $fwrite(32'h80000002,"%d: [dcache S3]: metawrite idx %x wmask %b meta %x%x:%x\n",c_1,
            io_metaWriteBus_req_bits_setIdx,io_metaWriteBus_req_bits_waymask,io_metaWriteBus_req_bits_data_valid,
            io_metaWriteBus_req_bits_data_dirty,io_metaWriteBus_req_bits_data_tag); // @[src/main/scala/utils/Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_3) begin
          $fwrite(32'h80000002,"[%d] CacheStage3_1: ",c_3); // @[src/main/scala/utils/Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_3) begin
          $fwrite(32'h80000002,
            " in.ready = %d, in.valid = %d, hit = %x, state = %d, addr = %x cmd:%d probe:%d isFinish:%d\n",io_in_ready,
            io_in_valid,hit,state,io_in_bits_req_addr,io_in_bits_req_cmd,probe,io_isFinish); // @[src/main/scala/utils/Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_3) begin
          $fwrite(32'h80000002,"[%d] CacheStage3_1: ",c_4); // @[src/main/scala/utils/Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_3) begin
          $fwrite(32'h80000002," out.valid:%d rdata:%x cmd:%d user:%x id:%x \n",io_out_valid,io_out_bits_rdata,
            io_out_bits_cmd,1'h0,1'h0); // @[src/main/scala/utils/Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_3) begin
          $fwrite(32'h80000002,"[%d] CacheStage3_1: ",c_5); // @[src/main/scala/utils/Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_3) begin
          $fwrite(32'h80000002," DHW: (%d, %d), data:%x setIdx:%x MHW:(%d, %d)\n",hitWrite,1'h1,dataHitWriteBus_x1_data,
            dataHitWriteBus_x3,metaHitWriteBus_x5,1'h1); // @[src/main/scala/utils/Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_3) begin
          $fwrite(32'h80000002,"[%d] CacheStage3_1: ",c_6); // @[src/main/scala/utils/Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_3) begin
          $fwrite(32'h80000002," DreadCache: %x \n",_T_89); // @[src/main/scala/utils/Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_3) begin
          $fwrite(32'h80000002,"[%d] CacheStage3_1: ",c_7); // @[src/main/scala/utils/Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_3) begin
          $fwrite(32'h80000002," useFD:%d isFD:%d FD:%x DreadArray:%x dataRead:%x inwaymask:%x FDwaymask:%x \n",
            useForwardData,io_in_bits_isForwardData,io_in_bits_forwardData_data_data,_dataReadArray_T_10,dataRead,
            io_in_bits_waymask,io_in_bits_forwardData_waymask); // @[src/main/scala/utils/Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_128 & _T_3) begin
          $fwrite(32'h80000002,"[%d] CacheStage3_1: ",c_8); // @[src/main/scala/utils/Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_128 & _T_3) begin
          $fwrite(32'h80000002,"[WB] waymask: %b data:%x setIdx:%x\n",io_dataWriteBus_req_bits_waymask,
            io_dataWriteBus_req_bits_data_data,io_dataWriteBus_req_bits_setIdx); // @[src/main/scala/utils/Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_140 & _T_3) begin
          $fwrite(32'h80000002,"[%d] CacheStage3_1: ",c_9); // @[src/main/scala/utils/Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_140 & _T_3) begin
          $fwrite(32'h80000002,"[COUTW] cnt %x addr %x data %x cmd %x size %x wmask %x tag %x idx %x waymask %b \n",
            writeBeatCnt_value,io_mem_req_bits_addr,io_mem_req_bits_wdata,io_mem_req_bits_cmd,io_mem_req_bits_size,
            io_mem_req_bits_wmask,addr_tag,addr_index,io_in_bits_waymask); // @[src/main/scala/utils/Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_152 & _T_3) begin
          $fwrite(32'h80000002,"[%d] CacheStage3_1: ",c_10); // @[src/main/scala/utils/Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_152 & _T_3) begin
          $fwrite(32'h80000002,"[COUTR] addr %x tag %x idx %x waymask %b \n",io_mem_req_bits_addr,addr_tag,addr_index,
            io_in_bits_waymask); // @[src/main/scala/utils/Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_164 & _T_3) begin
          $fwrite(32'h80000002,"[%d] CacheStage3_1: ",c_11); // @[src/main/scala/utils/Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_164 & _T_3) begin
          $fwrite(32'h80000002,"[COUTR] cnt %x data %x tag %x idx %x waymask %b \n",readBeatCnt_value,
            io_mem_resp_bits_rdata,addr_tag,addr_index,io_in_bits_waymask); // @[src/main/scala/utils/Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  writeL2BeatCnt_value = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  state = _RAND_1[3:0];
  _RAND_2 = {1{`RANDOM}};
  readBeatCnt_value = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  writeBeatCnt_value = _RAND_3[2:0];
  _RAND_4 = {1{`RANDOM}};
  state2 = _RAND_4[1:0];
  _RAND_5 = {2{`RANDOM}};
  dataWay_0_data = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  dataWay_1_data = _RAND_6[63:0];
  _RAND_7 = {2{`RANDOM}};
  dataWay_2_data = _RAND_7[63:0];
  _RAND_8 = {2{`RANDOM}};
  dataWay_3_data = _RAND_8[63:0];
  _RAND_9 = {1{`RANDOM}};
  afterFirstRead = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  alreadyOutFire = _RAND_10[0:0];
  _RAND_11 = {2{`RANDOM}};
  inRdataRegDemand = _RAND_11[63:0];
  _RAND_12 = {1{`RANDOM}};
  releaseLast_c_value = _RAND_12[2:0];
  _RAND_13 = {1{`RANDOM}};
  respToL1Last_c_value = _RAND_13[2:0];
  _RAND_14 = {2{`RANDOM}};
  c = _RAND_14[63:0];
  _RAND_15 = {2{`RANDOM}};
  c_1 = _RAND_15[63:0];
  _RAND_16 = {2{`RANDOM}};
  c_2 = _RAND_16[63:0];
  _RAND_17 = {2{`RANDOM}};
  c_3 = _RAND_17[63:0];
  _RAND_18 = {2{`RANDOM}};
  c_4 = _RAND_18[63:0];
  _RAND_19 = {2{`RANDOM}};
  c_5 = _RAND_19[63:0];
  _RAND_20 = {2{`RANDOM}};
  c_6 = _RAND_20[63:0];
  _RAND_21 = {2{`RANDOM}};
  c_7 = _RAND_21[63:0];
  _RAND_22 = {2{`RANDOM}};
  c_8 = _RAND_22[63:0];
  _RAND_23 = {2{`RANDOM}};
  c_9 = _RAND_23[63:0];
  _RAND_24 = {2{`RANDOM}};
  c_10 = _RAND_24[63:0];
  _RAND_25 = {2{`RANDOM}};
  c_11 = _RAND_25[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Arbiter_9(
  output        io_in_0_ready, // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
  input         io_in_0_valid, // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
  input  [31:0] io_in_0_bits_addr, // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
  input  [2:0]  io_in_0_bits_size, // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
  input  [3:0]  io_in_0_bits_cmd, // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
  input  [7:0]  io_in_0_bits_wmask, // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
  input  [63:0] io_in_0_bits_wdata, // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
  output        io_in_1_ready, // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
  input         io_in_1_valid, // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
  input  [31:0] io_in_1_bits_addr, // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
  input  [2:0]  io_in_1_bits_size, // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
  input  [3:0]  io_in_1_bits_cmd, // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
  input  [7:0]  io_in_1_bits_wmask, // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
  input  [63:0] io_in_1_bits_wdata, // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
  input         io_out_ready, // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
  output        io_out_valid, // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
  output [31:0] io_out_bits_addr, // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
  output [2:0]  io_out_bits_size, // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
  output [3:0]  io_out_bits_cmd, // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
  output [7:0]  io_out_bits_wmask, // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
  output [63:0] io_out_bits_wdata // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
);
  wire  grant_1 = ~io_in_0_valid; // @[src/main/scala/chisel3/util/Arbiter.scala 45:78]
  assign io_in_0_ready = io_out_ready; // @[src/main/scala/chisel3/util/Arbiter.scala 147:19]
  assign io_in_1_ready = grant_1 & io_out_ready; // @[src/main/scala/chisel3/util/Arbiter.scala 147:19]
  assign io_out_valid = ~grant_1 | io_in_1_valid; // @[src/main/scala/chisel3/util/Arbiter.scala 148:31]
  assign io_out_bits_addr = io_in_0_valid ? io_in_0_bits_addr : io_in_1_bits_addr; // @[src/main/scala/chisel3/util/Arbiter.scala 137:15 139:26 141:19]
  assign io_out_bits_size = io_in_0_valid ? io_in_0_bits_size : io_in_1_bits_size; // @[src/main/scala/chisel3/util/Arbiter.scala 137:15 139:26 141:19]
  assign io_out_bits_cmd = io_in_0_valid ? io_in_0_bits_cmd : io_in_1_bits_cmd; // @[src/main/scala/chisel3/util/Arbiter.scala 137:15 139:26 141:19]
  assign io_out_bits_wmask = io_in_0_valid ? io_in_0_bits_wmask : io_in_1_bits_wmask; // @[src/main/scala/chisel3/util/Arbiter.scala 137:15 139:26 141:19]
  assign io_out_bits_wdata = io_in_0_valid ? io_in_0_bits_wdata : io_in_1_bits_wdata; // @[src/main/scala/chisel3/util/Arbiter.scala 137:15 139:26 141:19]
endmodule
module Cache_1(
  input         clock,
  input         reset,
  output        io_in_req_ready, // @[src/main/scala/nutcore/mem/Cache.scala 122:14]
  input         io_in_req_valid, // @[src/main/scala/nutcore/mem/Cache.scala 122:14]
  input  [31:0] io_in_req_bits_addr, // @[src/main/scala/nutcore/mem/Cache.scala 122:14]
  input  [2:0]  io_in_req_bits_size, // @[src/main/scala/nutcore/mem/Cache.scala 122:14]
  input  [3:0]  io_in_req_bits_cmd, // @[src/main/scala/nutcore/mem/Cache.scala 122:14]
  input  [7:0]  io_in_req_bits_wmask, // @[src/main/scala/nutcore/mem/Cache.scala 122:14]
  input  [63:0] io_in_req_bits_wdata, // @[src/main/scala/nutcore/mem/Cache.scala 122:14]
  input         io_in_resp_ready, // @[src/main/scala/nutcore/mem/Cache.scala 122:14]
  output        io_in_resp_valid, // @[src/main/scala/nutcore/mem/Cache.scala 122:14]
  output [3:0]  io_in_resp_bits_cmd, // @[src/main/scala/nutcore/mem/Cache.scala 122:14]
  output [63:0] io_in_resp_bits_rdata, // @[src/main/scala/nutcore/mem/Cache.scala 122:14]
  input         io_out_mem_req_ready, // @[src/main/scala/nutcore/mem/Cache.scala 122:14]
  output        io_out_mem_req_valid, // @[src/main/scala/nutcore/mem/Cache.scala 122:14]
  output [31:0] io_out_mem_req_bits_addr, // @[src/main/scala/nutcore/mem/Cache.scala 122:14]
  output [3:0]  io_out_mem_req_bits_cmd, // @[src/main/scala/nutcore/mem/Cache.scala 122:14]
  output [63:0] io_out_mem_req_bits_wdata, // @[src/main/scala/nutcore/mem/Cache.scala 122:14]
  input         io_out_mem_resp_valid, // @[src/main/scala/nutcore/mem/Cache.scala 122:14]
  input  [3:0]  io_out_mem_resp_bits_cmd, // @[src/main/scala/nutcore/mem/Cache.scala 122:14]
  input  [63:0] io_out_mem_resp_bits_rdata, // @[src/main/scala/nutcore/mem/Cache.scala 122:14]
  output        io_out_coh_req_ready, // @[src/main/scala/nutcore/mem/Cache.scala 122:14]
  input         io_out_coh_req_valid, // @[src/main/scala/nutcore/mem/Cache.scala 122:14]
  input  [31:0] io_out_coh_req_bits_addr, // @[src/main/scala/nutcore/mem/Cache.scala 122:14]
  input  [63:0] io_out_coh_req_bits_wdata, // @[src/main/scala/nutcore/mem/Cache.scala 122:14]
  output        io_out_coh_resp_valid, // @[src/main/scala/nutcore/mem/Cache.scala 122:14]
  output [3:0]  io_out_coh_resp_bits_cmd, // @[src/main/scala/nutcore/mem/Cache.scala 122:14]
  output [63:0] io_out_coh_resp_bits_rdata, // @[src/main/scala/nutcore/mem/Cache.scala 122:14]
  input         io_mmio_req_ready, // @[src/main/scala/nutcore/mem/Cache.scala 122:14]
  output        io_mmio_req_valid, // @[src/main/scala/nutcore/mem/Cache.scala 122:14]
  output [31:0] io_mmio_req_bits_addr, // @[src/main/scala/nutcore/mem/Cache.scala 122:14]
  output [2:0]  io_mmio_req_bits_size, // @[src/main/scala/nutcore/mem/Cache.scala 122:14]
  output [3:0]  io_mmio_req_bits_cmd, // @[src/main/scala/nutcore/mem/Cache.scala 122:14]
  output [7:0]  io_mmio_req_bits_wmask, // @[src/main/scala/nutcore/mem/Cache.scala 122:14]
  output [63:0] io_mmio_req_bits_wdata, // @[src/main/scala/nutcore/mem/Cache.scala 122:14]
  input         io_mmio_resp_valid, // @[src/main/scala/nutcore/mem/Cache.scala 122:14]
  input  [63:0] io_mmio_resp_bits_rdata, // @[src/main/scala/nutcore/mem/Cache.scala 122:14]
  output        io_empty, // @[src/main/scala/nutcore/mem/Cache.scala 122:14]
  input         DISPLAY_ENABLE,
  output        _WIRE_17
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [63:0] _RAND_24;
  reg [63:0] _RAND_25;
  reg [63:0] _RAND_26;
  reg [63:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [63:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [63:0] _RAND_34;
  reg [63:0] _RAND_35;
  reg [63:0] _RAND_36;
  reg [63:0] _RAND_37;
  reg [63:0] _RAND_38;
`endif // RANDOMIZE_REG_INIT
  wire  s1_clock; // @[src/main/scala/nutcore/mem/Cache.scala 480:18]
  wire  s1_reset; // @[src/main/scala/nutcore/mem/Cache.scala 480:18]
  wire  s1_io_in_ready; // @[src/main/scala/nutcore/mem/Cache.scala 480:18]
  wire  s1_io_in_valid; // @[src/main/scala/nutcore/mem/Cache.scala 480:18]
  wire [31:0] s1_io_in_bits_addr; // @[src/main/scala/nutcore/mem/Cache.scala 480:18]
  wire [2:0] s1_io_in_bits_size; // @[src/main/scala/nutcore/mem/Cache.scala 480:18]
  wire [3:0] s1_io_in_bits_cmd; // @[src/main/scala/nutcore/mem/Cache.scala 480:18]
  wire [7:0] s1_io_in_bits_wmask; // @[src/main/scala/nutcore/mem/Cache.scala 480:18]
  wire [63:0] s1_io_in_bits_wdata; // @[src/main/scala/nutcore/mem/Cache.scala 480:18]
  wire  s1_io_out_ready; // @[src/main/scala/nutcore/mem/Cache.scala 480:18]
  wire  s1_io_out_valid; // @[src/main/scala/nutcore/mem/Cache.scala 480:18]
  wire [31:0] s1_io_out_bits_req_addr; // @[src/main/scala/nutcore/mem/Cache.scala 480:18]
  wire [2:0] s1_io_out_bits_req_size; // @[src/main/scala/nutcore/mem/Cache.scala 480:18]
  wire [3:0] s1_io_out_bits_req_cmd; // @[src/main/scala/nutcore/mem/Cache.scala 480:18]
  wire [7:0] s1_io_out_bits_req_wmask; // @[src/main/scala/nutcore/mem/Cache.scala 480:18]
  wire [63:0] s1_io_out_bits_req_wdata; // @[src/main/scala/nutcore/mem/Cache.scala 480:18]
  wire  s1_io_metaReadBus_req_ready; // @[src/main/scala/nutcore/mem/Cache.scala 480:18]
  wire  s1_io_metaReadBus_req_valid; // @[src/main/scala/nutcore/mem/Cache.scala 480:18]
  wire [6:0] s1_io_metaReadBus_req_bits_setIdx; // @[src/main/scala/nutcore/mem/Cache.scala 480:18]
  wire [18:0] s1_io_metaReadBus_resp_data_0_tag; // @[src/main/scala/nutcore/mem/Cache.scala 480:18]
  wire  s1_io_metaReadBus_resp_data_0_valid; // @[src/main/scala/nutcore/mem/Cache.scala 480:18]
  wire  s1_io_metaReadBus_resp_data_0_dirty; // @[src/main/scala/nutcore/mem/Cache.scala 480:18]
  wire [18:0] s1_io_metaReadBus_resp_data_1_tag; // @[src/main/scala/nutcore/mem/Cache.scala 480:18]
  wire  s1_io_metaReadBus_resp_data_1_valid; // @[src/main/scala/nutcore/mem/Cache.scala 480:18]
  wire  s1_io_metaReadBus_resp_data_1_dirty; // @[src/main/scala/nutcore/mem/Cache.scala 480:18]
  wire [18:0] s1_io_metaReadBus_resp_data_2_tag; // @[src/main/scala/nutcore/mem/Cache.scala 480:18]
  wire  s1_io_metaReadBus_resp_data_2_valid; // @[src/main/scala/nutcore/mem/Cache.scala 480:18]
  wire  s1_io_metaReadBus_resp_data_2_dirty; // @[src/main/scala/nutcore/mem/Cache.scala 480:18]
  wire [18:0] s1_io_metaReadBus_resp_data_3_tag; // @[src/main/scala/nutcore/mem/Cache.scala 480:18]
  wire  s1_io_metaReadBus_resp_data_3_valid; // @[src/main/scala/nutcore/mem/Cache.scala 480:18]
  wire  s1_io_metaReadBus_resp_data_3_dirty; // @[src/main/scala/nutcore/mem/Cache.scala 480:18]
  wire  s1_io_dataReadBus_req_ready; // @[src/main/scala/nutcore/mem/Cache.scala 480:18]
  wire  s1_io_dataReadBus_req_valid; // @[src/main/scala/nutcore/mem/Cache.scala 480:18]
  wire [9:0] s1_io_dataReadBus_req_bits_setIdx; // @[src/main/scala/nutcore/mem/Cache.scala 480:18]
  wire [63:0] s1_io_dataReadBus_resp_data_0_data; // @[src/main/scala/nutcore/mem/Cache.scala 480:18]
  wire [63:0] s1_io_dataReadBus_resp_data_1_data; // @[src/main/scala/nutcore/mem/Cache.scala 480:18]
  wire [63:0] s1_io_dataReadBus_resp_data_2_data; // @[src/main/scala/nutcore/mem/Cache.scala 480:18]
  wire [63:0] s1_io_dataReadBus_resp_data_3_data; // @[src/main/scala/nutcore/mem/Cache.scala 480:18]
  wire  s1_DISPLAY_ENABLE; // @[src/main/scala/nutcore/mem/Cache.scala 480:18]
  wire  s2_clock; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire  s2_reset; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire  s2_io_in_ready; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire  s2_io_in_valid; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire [31:0] s2_io_in_bits_req_addr; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire [2:0] s2_io_in_bits_req_size; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire [3:0] s2_io_in_bits_req_cmd; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire [7:0] s2_io_in_bits_req_wmask; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire [63:0] s2_io_in_bits_req_wdata; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire  s2_io_out_ready; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire  s2_io_out_valid; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire [31:0] s2_io_out_bits_req_addr; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire [2:0] s2_io_out_bits_req_size; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire [3:0] s2_io_out_bits_req_cmd; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire [7:0] s2_io_out_bits_req_wmask; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire [63:0] s2_io_out_bits_req_wdata; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire [18:0] s2_io_out_bits_metas_0_tag; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire  s2_io_out_bits_metas_0_valid; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire  s2_io_out_bits_metas_0_dirty; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire [18:0] s2_io_out_bits_metas_1_tag; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire  s2_io_out_bits_metas_1_valid; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire  s2_io_out_bits_metas_1_dirty; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire [18:0] s2_io_out_bits_metas_2_tag; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire  s2_io_out_bits_metas_2_valid; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire  s2_io_out_bits_metas_2_dirty; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire [18:0] s2_io_out_bits_metas_3_tag; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire  s2_io_out_bits_metas_3_valid; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire  s2_io_out_bits_metas_3_dirty; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire [63:0] s2_io_out_bits_datas_0_data; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire [63:0] s2_io_out_bits_datas_1_data; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire [63:0] s2_io_out_bits_datas_2_data; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire [63:0] s2_io_out_bits_datas_3_data; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire  s2_io_out_bits_hit; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire [3:0] s2_io_out_bits_waymask; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire  s2_io_out_bits_mmio; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire  s2_io_out_bits_isForwardData; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire [63:0] s2_io_out_bits_forwardData_data_data; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire [3:0] s2_io_out_bits_forwardData_waymask; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire [18:0] s2_io_metaReadResp_0_tag; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire  s2_io_metaReadResp_0_valid; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire  s2_io_metaReadResp_0_dirty; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire [18:0] s2_io_metaReadResp_1_tag; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire  s2_io_metaReadResp_1_valid; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire  s2_io_metaReadResp_1_dirty; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire [18:0] s2_io_metaReadResp_2_tag; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire  s2_io_metaReadResp_2_valid; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire  s2_io_metaReadResp_2_dirty; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire [18:0] s2_io_metaReadResp_3_tag; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire  s2_io_metaReadResp_3_valid; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire  s2_io_metaReadResp_3_dirty; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire [63:0] s2_io_dataReadResp_0_data; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire [63:0] s2_io_dataReadResp_1_data; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire [63:0] s2_io_dataReadResp_2_data; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire [63:0] s2_io_dataReadResp_3_data; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire  s2_io_metaWriteBus_req_valid; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire [6:0] s2_io_metaWriteBus_req_bits_setIdx; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire [18:0] s2_io_metaWriteBus_req_bits_data_tag; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire  s2_io_metaWriteBus_req_bits_data_dirty; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire [3:0] s2_io_metaWriteBus_req_bits_waymask; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire  s2_io_dataWriteBus_req_valid; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire [9:0] s2_io_dataWriteBus_req_bits_setIdx; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire [63:0] s2_io_dataWriteBus_req_bits_data_data; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire [3:0] s2_io_dataWriteBus_req_bits_waymask; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire  s2_DISPLAY_ENABLE; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire  s3_clock; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire  s3_reset; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire  s3_io_in_ready; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire  s3_io_in_valid; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire [31:0] s3_io_in_bits_req_addr; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire [2:0] s3_io_in_bits_req_size; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire [3:0] s3_io_in_bits_req_cmd; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire [7:0] s3_io_in_bits_req_wmask; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire [63:0] s3_io_in_bits_req_wdata; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire [18:0] s3_io_in_bits_metas_0_tag; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire  s3_io_in_bits_metas_0_valid; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire  s3_io_in_bits_metas_0_dirty; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire [18:0] s3_io_in_bits_metas_1_tag; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire  s3_io_in_bits_metas_1_valid; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire  s3_io_in_bits_metas_1_dirty; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire [18:0] s3_io_in_bits_metas_2_tag; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire  s3_io_in_bits_metas_2_valid; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire  s3_io_in_bits_metas_2_dirty; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire [18:0] s3_io_in_bits_metas_3_tag; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire  s3_io_in_bits_metas_3_valid; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire  s3_io_in_bits_metas_3_dirty; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire [63:0] s3_io_in_bits_datas_0_data; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire [63:0] s3_io_in_bits_datas_1_data; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire [63:0] s3_io_in_bits_datas_2_data; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire [63:0] s3_io_in_bits_datas_3_data; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire  s3_io_in_bits_hit; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire [3:0] s3_io_in_bits_waymask; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire  s3_io_in_bits_mmio; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire  s3_io_in_bits_isForwardData; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire [63:0] s3_io_in_bits_forwardData_data_data; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire [3:0] s3_io_in_bits_forwardData_waymask; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire  s3_io_out_ready; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire  s3_io_out_valid; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire [3:0] s3_io_out_bits_cmd; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire [63:0] s3_io_out_bits_rdata; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire  s3_io_isFinish; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire  s3_io_dataReadBus_req_ready; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire  s3_io_dataReadBus_req_valid; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire [9:0] s3_io_dataReadBus_req_bits_setIdx; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire [63:0] s3_io_dataReadBus_resp_data_0_data; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire [63:0] s3_io_dataReadBus_resp_data_1_data; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire [63:0] s3_io_dataReadBus_resp_data_2_data; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire [63:0] s3_io_dataReadBus_resp_data_3_data; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire  s3_io_dataWriteBus_req_valid; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire [9:0] s3_io_dataWriteBus_req_bits_setIdx; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire [63:0] s3_io_dataWriteBus_req_bits_data_data; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire [3:0] s3_io_dataWriteBus_req_bits_waymask; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire  s3_io_metaWriteBus_req_valid; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire [6:0] s3_io_metaWriteBus_req_bits_setIdx; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire [18:0] s3_io_metaWriteBus_req_bits_data_tag; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire  s3_io_metaWriteBus_req_bits_data_valid; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire  s3_io_metaWriteBus_req_bits_data_dirty; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire [3:0] s3_io_metaWriteBus_req_bits_waymask; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire  s3_io_mem_req_ready; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire  s3_io_mem_req_valid; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire [31:0] s3_io_mem_req_bits_addr; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire [2:0] s3_io_mem_req_bits_size; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire [3:0] s3_io_mem_req_bits_cmd; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire [7:0] s3_io_mem_req_bits_wmask; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire [63:0] s3_io_mem_req_bits_wdata; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire  s3_io_mem_resp_ready; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire  s3_io_mem_resp_valid; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire [3:0] s3_io_mem_resp_bits_cmd; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire [63:0] s3_io_mem_resp_bits_rdata; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire  s3_io_mmio_req_ready; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire  s3_io_mmio_req_valid; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire [31:0] s3_io_mmio_req_bits_addr; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire [2:0] s3_io_mmio_req_bits_size; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire [3:0] s3_io_mmio_req_bits_cmd; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire [7:0] s3_io_mmio_req_bits_wmask; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire [63:0] s3_io_mmio_req_bits_wdata; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire  s3_io_mmio_resp_ready; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire  s3_io_mmio_resp_valid; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire [63:0] s3_io_mmio_resp_bits_rdata; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire  s3_io_cohResp_valid; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire [3:0] s3_io_cohResp_bits_cmd; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire [63:0] s3_io_cohResp_bits_rdata; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire  s3_io_dataReadRespToL1; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire  s3_DISPLAY_ENABLE; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire  s3__WIRE_19; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire  metaArray_clock; // @[src/main/scala/nutcore/mem/Cache.scala 483:25]
  wire  metaArray_reset; // @[src/main/scala/nutcore/mem/Cache.scala 483:25]
  wire  metaArray_io_r_0_req_ready; // @[src/main/scala/nutcore/mem/Cache.scala 483:25]
  wire  metaArray_io_r_0_req_valid; // @[src/main/scala/nutcore/mem/Cache.scala 483:25]
  wire [6:0] metaArray_io_r_0_req_bits_setIdx; // @[src/main/scala/nutcore/mem/Cache.scala 483:25]
  wire [18:0] metaArray_io_r_0_resp_data_0_tag; // @[src/main/scala/nutcore/mem/Cache.scala 483:25]
  wire  metaArray_io_r_0_resp_data_0_valid; // @[src/main/scala/nutcore/mem/Cache.scala 483:25]
  wire  metaArray_io_r_0_resp_data_0_dirty; // @[src/main/scala/nutcore/mem/Cache.scala 483:25]
  wire [18:0] metaArray_io_r_0_resp_data_1_tag; // @[src/main/scala/nutcore/mem/Cache.scala 483:25]
  wire  metaArray_io_r_0_resp_data_1_valid; // @[src/main/scala/nutcore/mem/Cache.scala 483:25]
  wire  metaArray_io_r_0_resp_data_1_dirty; // @[src/main/scala/nutcore/mem/Cache.scala 483:25]
  wire [18:0] metaArray_io_r_0_resp_data_2_tag; // @[src/main/scala/nutcore/mem/Cache.scala 483:25]
  wire  metaArray_io_r_0_resp_data_2_valid; // @[src/main/scala/nutcore/mem/Cache.scala 483:25]
  wire  metaArray_io_r_0_resp_data_2_dirty; // @[src/main/scala/nutcore/mem/Cache.scala 483:25]
  wire [18:0] metaArray_io_r_0_resp_data_3_tag; // @[src/main/scala/nutcore/mem/Cache.scala 483:25]
  wire  metaArray_io_r_0_resp_data_3_valid; // @[src/main/scala/nutcore/mem/Cache.scala 483:25]
  wire  metaArray_io_r_0_resp_data_3_dirty; // @[src/main/scala/nutcore/mem/Cache.scala 483:25]
  wire  metaArray_io_w_req_valid; // @[src/main/scala/nutcore/mem/Cache.scala 483:25]
  wire [6:0] metaArray_io_w_req_bits_setIdx; // @[src/main/scala/nutcore/mem/Cache.scala 483:25]
  wire [18:0] metaArray_io_w_req_bits_data_tag; // @[src/main/scala/nutcore/mem/Cache.scala 483:25]
  wire  metaArray_io_w_req_bits_data_dirty; // @[src/main/scala/nutcore/mem/Cache.scala 483:25]
  wire [3:0] metaArray_io_w_req_bits_waymask; // @[src/main/scala/nutcore/mem/Cache.scala 483:25]
  wire  dataArray_clock; // @[src/main/scala/nutcore/mem/Cache.scala 484:25]
  wire  dataArray_reset; // @[src/main/scala/nutcore/mem/Cache.scala 484:25]
  wire  dataArray_io_r_0_req_ready; // @[src/main/scala/nutcore/mem/Cache.scala 484:25]
  wire  dataArray_io_r_0_req_valid; // @[src/main/scala/nutcore/mem/Cache.scala 484:25]
  wire [9:0] dataArray_io_r_0_req_bits_setIdx; // @[src/main/scala/nutcore/mem/Cache.scala 484:25]
  wire [63:0] dataArray_io_r_0_resp_data_0_data; // @[src/main/scala/nutcore/mem/Cache.scala 484:25]
  wire [63:0] dataArray_io_r_0_resp_data_1_data; // @[src/main/scala/nutcore/mem/Cache.scala 484:25]
  wire [63:0] dataArray_io_r_0_resp_data_2_data; // @[src/main/scala/nutcore/mem/Cache.scala 484:25]
  wire [63:0] dataArray_io_r_0_resp_data_3_data; // @[src/main/scala/nutcore/mem/Cache.scala 484:25]
  wire  dataArray_io_r_1_req_ready; // @[src/main/scala/nutcore/mem/Cache.scala 484:25]
  wire  dataArray_io_r_1_req_valid; // @[src/main/scala/nutcore/mem/Cache.scala 484:25]
  wire [9:0] dataArray_io_r_1_req_bits_setIdx; // @[src/main/scala/nutcore/mem/Cache.scala 484:25]
  wire [63:0] dataArray_io_r_1_resp_data_0_data; // @[src/main/scala/nutcore/mem/Cache.scala 484:25]
  wire [63:0] dataArray_io_r_1_resp_data_1_data; // @[src/main/scala/nutcore/mem/Cache.scala 484:25]
  wire [63:0] dataArray_io_r_1_resp_data_2_data; // @[src/main/scala/nutcore/mem/Cache.scala 484:25]
  wire [63:0] dataArray_io_r_1_resp_data_3_data; // @[src/main/scala/nutcore/mem/Cache.scala 484:25]
  wire  dataArray_io_w_req_valid; // @[src/main/scala/nutcore/mem/Cache.scala 484:25]
  wire [9:0] dataArray_io_w_req_bits_setIdx; // @[src/main/scala/nutcore/mem/Cache.scala 484:25]
  wire [63:0] dataArray_io_w_req_bits_data_data; // @[src/main/scala/nutcore/mem/Cache.scala 484:25]
  wire [3:0] dataArray_io_w_req_bits_waymask; // @[src/main/scala/nutcore/mem/Cache.scala 484:25]
  wire  arb_io_in_0_ready; // @[src/main/scala/nutcore/mem/Cache.scala 493:19]
  wire  arb_io_in_0_valid; // @[src/main/scala/nutcore/mem/Cache.scala 493:19]
  wire [31:0] arb_io_in_0_bits_addr; // @[src/main/scala/nutcore/mem/Cache.scala 493:19]
  wire [2:0] arb_io_in_0_bits_size; // @[src/main/scala/nutcore/mem/Cache.scala 493:19]
  wire [3:0] arb_io_in_0_bits_cmd; // @[src/main/scala/nutcore/mem/Cache.scala 493:19]
  wire [7:0] arb_io_in_0_bits_wmask; // @[src/main/scala/nutcore/mem/Cache.scala 493:19]
  wire [63:0] arb_io_in_0_bits_wdata; // @[src/main/scala/nutcore/mem/Cache.scala 493:19]
  wire  arb_io_in_1_ready; // @[src/main/scala/nutcore/mem/Cache.scala 493:19]
  wire  arb_io_in_1_valid; // @[src/main/scala/nutcore/mem/Cache.scala 493:19]
  wire [31:0] arb_io_in_1_bits_addr; // @[src/main/scala/nutcore/mem/Cache.scala 493:19]
  wire [2:0] arb_io_in_1_bits_size; // @[src/main/scala/nutcore/mem/Cache.scala 493:19]
  wire [3:0] arb_io_in_1_bits_cmd; // @[src/main/scala/nutcore/mem/Cache.scala 493:19]
  wire [7:0] arb_io_in_1_bits_wmask; // @[src/main/scala/nutcore/mem/Cache.scala 493:19]
  wire [63:0] arb_io_in_1_bits_wdata; // @[src/main/scala/nutcore/mem/Cache.scala 493:19]
  wire  arb_io_out_ready; // @[src/main/scala/nutcore/mem/Cache.scala 493:19]
  wire  arb_io_out_valid; // @[src/main/scala/nutcore/mem/Cache.scala 493:19]
  wire [31:0] arb_io_out_bits_addr; // @[src/main/scala/nutcore/mem/Cache.scala 493:19]
  wire [2:0] arb_io_out_bits_size; // @[src/main/scala/nutcore/mem/Cache.scala 493:19]
  wire [3:0] arb_io_out_bits_cmd; // @[src/main/scala/nutcore/mem/Cache.scala 493:19]
  wire [7:0] arb_io_out_bits_wmask; // @[src/main/scala/nutcore/mem/Cache.scala 493:19]
  wire [63:0] arb_io_out_bits_wdata; // @[src/main/scala/nutcore/mem/Cache.scala 493:19]
  wire  _T = s2_io_out_ready & s2_io_out_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  reg  valid; // @[src/main/scala/utils/Pipeline.scala 24:24]
  wire  _GEN_0 = _T ? 1'h0 : valid; // @[src/main/scala/utils/Pipeline.scala 24:24 25:{25,33}]
  wire  _T_2 = s1_io_out_valid & s2_io_in_ready; // @[src/main/scala/utils/Pipeline.scala 26:22]
  wire  _GEN_1 = s1_io_out_valid & s2_io_in_ready | _GEN_0; // @[src/main/scala/utils/Pipeline.scala 26:{38,46}]
  reg [31:0] s2_io_in_bits_r_req_addr; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg [2:0] s2_io_in_bits_r_req_size; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg [3:0] s2_io_in_bits_r_req_cmd; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg [7:0] s2_io_in_bits_r_req_wmask; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg [63:0] s2_io_in_bits_r_req_wdata; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg  valid_1; // @[src/main/scala/utils/Pipeline.scala 24:24]
  wire  _GEN_8 = s3_io_isFinish ? 1'h0 : valid_1; // @[src/main/scala/utils/Pipeline.scala 24:24 25:{25,33}]
  wire  _T_4 = s2_io_out_valid & s3_io_in_ready; // @[src/main/scala/utils/Pipeline.scala 26:22]
  wire  _GEN_9 = s2_io_out_valid & s3_io_in_ready | _GEN_8; // @[src/main/scala/utils/Pipeline.scala 26:{38,46}]
  reg [31:0] s3_io_in_bits_r_req_addr; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg [2:0] s3_io_in_bits_r_req_size; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg [3:0] s3_io_in_bits_r_req_cmd; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg [7:0] s3_io_in_bits_r_req_wmask; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg [63:0] s3_io_in_bits_r_req_wdata; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg [18:0] s3_io_in_bits_r_metas_0_tag; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg  s3_io_in_bits_r_metas_0_valid; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg  s3_io_in_bits_r_metas_0_dirty; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg [18:0] s3_io_in_bits_r_metas_1_tag; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg  s3_io_in_bits_r_metas_1_valid; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg  s3_io_in_bits_r_metas_1_dirty; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg [18:0] s3_io_in_bits_r_metas_2_tag; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg  s3_io_in_bits_r_metas_2_valid; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg  s3_io_in_bits_r_metas_2_dirty; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg [18:0] s3_io_in_bits_r_metas_3_tag; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg  s3_io_in_bits_r_metas_3_valid; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg  s3_io_in_bits_r_metas_3_dirty; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg [63:0] s3_io_in_bits_r_datas_0_data; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg [63:0] s3_io_in_bits_r_datas_1_data; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg [63:0] s3_io_in_bits_r_datas_2_data; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg [63:0] s3_io_in_bits_r_datas_3_data; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg  s3_io_in_bits_r_hit; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg [3:0] s3_io_in_bits_r_waymask; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg  s3_io_in_bits_r_mmio; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg  s3_io_in_bits_r_isForwardData; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg [63:0] s3_io_in_bits_r_forwardData_data_data; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg [3:0] s3_io_in_bits_r_forwardData_waymask; // @[src/main/scala/utils/Pipeline.scala 30:28]
  wire  _io_in_resp_valid_T = s3_io_out_bits_cmd == 4'h4; // @[src/main/scala/bus/simplebus/SimpleBus.scala 95:24]
  reg [63:0] c; // @[src/main/scala/utils/GTimer.scala 24:20]
  wire [63:0] _c_T_1 = c + 64'h1; // @[src/main/scala/utils/GTimer.scala 25:12]
  wire  _T_7 = ~reset; // @[src/main/scala/utils/Debug.scala 56:24]
  reg [63:0] c_1; // @[src/main/scala/utils/GTimer.scala 24:20]
  wire [63:0] _c_T_3 = c_1 + 64'h1; // @[src/main/scala/utils/GTimer.scala 25:12]
  reg [63:0] c_2; // @[src/main/scala/utils/GTimer.scala 24:20]
  wire [63:0] _c_T_5 = c_2 + 64'h1; // @[src/main/scala/utils/GTimer.scala 25:12]
  reg [63:0] c_3; // @[src/main/scala/utils/GTimer.scala 24:20]
  wire [63:0] _c_T_7 = c_3 + 64'h1; // @[src/main/scala/utils/GTimer.scala 25:12]
  reg [63:0] c_4; // @[src/main/scala/utils/GTimer.scala 24:20]
  wire [63:0] _c_T_9 = c_4 + 64'h1; // @[src/main/scala/utils/GTimer.scala 25:12]
  wire  _GEN_39 = s1_io_in_valid & DISPLAY_ENABLE; // @[src/main/scala/utils/Debug.scala 56:24]
  wire  _GEN_41 = s2_io_in_valid & DISPLAY_ENABLE; // @[src/main/scala/utils/Debug.scala 56:24]
  wire  _GEN_43 = s3_io_in_valid & DISPLAY_ENABLE; // @[src/main/scala/utils/Debug.scala 56:24]
  CacheStage1_1 s1 ( // @[src/main/scala/nutcore/mem/Cache.scala 480:18]
    .clock(s1_clock),
    .reset(s1_reset),
    .io_in_ready(s1_io_in_ready),
    .io_in_valid(s1_io_in_valid),
    .io_in_bits_addr(s1_io_in_bits_addr),
    .io_in_bits_size(s1_io_in_bits_size),
    .io_in_bits_cmd(s1_io_in_bits_cmd),
    .io_in_bits_wmask(s1_io_in_bits_wmask),
    .io_in_bits_wdata(s1_io_in_bits_wdata),
    .io_out_ready(s1_io_out_ready),
    .io_out_valid(s1_io_out_valid),
    .io_out_bits_req_addr(s1_io_out_bits_req_addr),
    .io_out_bits_req_size(s1_io_out_bits_req_size),
    .io_out_bits_req_cmd(s1_io_out_bits_req_cmd),
    .io_out_bits_req_wmask(s1_io_out_bits_req_wmask),
    .io_out_bits_req_wdata(s1_io_out_bits_req_wdata),
    .io_metaReadBus_req_ready(s1_io_metaReadBus_req_ready),
    .io_metaReadBus_req_valid(s1_io_metaReadBus_req_valid),
    .io_metaReadBus_req_bits_setIdx(s1_io_metaReadBus_req_bits_setIdx),
    .io_metaReadBus_resp_data_0_tag(s1_io_metaReadBus_resp_data_0_tag),
    .io_metaReadBus_resp_data_0_valid(s1_io_metaReadBus_resp_data_0_valid),
    .io_metaReadBus_resp_data_0_dirty(s1_io_metaReadBus_resp_data_0_dirty),
    .io_metaReadBus_resp_data_1_tag(s1_io_metaReadBus_resp_data_1_tag),
    .io_metaReadBus_resp_data_1_valid(s1_io_metaReadBus_resp_data_1_valid),
    .io_metaReadBus_resp_data_1_dirty(s1_io_metaReadBus_resp_data_1_dirty),
    .io_metaReadBus_resp_data_2_tag(s1_io_metaReadBus_resp_data_2_tag),
    .io_metaReadBus_resp_data_2_valid(s1_io_metaReadBus_resp_data_2_valid),
    .io_metaReadBus_resp_data_2_dirty(s1_io_metaReadBus_resp_data_2_dirty),
    .io_metaReadBus_resp_data_3_tag(s1_io_metaReadBus_resp_data_3_tag),
    .io_metaReadBus_resp_data_3_valid(s1_io_metaReadBus_resp_data_3_valid),
    .io_metaReadBus_resp_data_3_dirty(s1_io_metaReadBus_resp_data_3_dirty),
    .io_dataReadBus_req_ready(s1_io_dataReadBus_req_ready),
    .io_dataReadBus_req_valid(s1_io_dataReadBus_req_valid),
    .io_dataReadBus_req_bits_setIdx(s1_io_dataReadBus_req_bits_setIdx),
    .io_dataReadBus_resp_data_0_data(s1_io_dataReadBus_resp_data_0_data),
    .io_dataReadBus_resp_data_1_data(s1_io_dataReadBus_resp_data_1_data),
    .io_dataReadBus_resp_data_2_data(s1_io_dataReadBus_resp_data_2_data),
    .io_dataReadBus_resp_data_3_data(s1_io_dataReadBus_resp_data_3_data),
    .DISPLAY_ENABLE(s1_DISPLAY_ENABLE)
  );
  CacheStage2_1 s2 ( // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
    .clock(s2_clock),
    .reset(s2_reset),
    .io_in_ready(s2_io_in_ready),
    .io_in_valid(s2_io_in_valid),
    .io_in_bits_req_addr(s2_io_in_bits_req_addr),
    .io_in_bits_req_size(s2_io_in_bits_req_size),
    .io_in_bits_req_cmd(s2_io_in_bits_req_cmd),
    .io_in_bits_req_wmask(s2_io_in_bits_req_wmask),
    .io_in_bits_req_wdata(s2_io_in_bits_req_wdata),
    .io_out_ready(s2_io_out_ready),
    .io_out_valid(s2_io_out_valid),
    .io_out_bits_req_addr(s2_io_out_bits_req_addr),
    .io_out_bits_req_size(s2_io_out_bits_req_size),
    .io_out_bits_req_cmd(s2_io_out_bits_req_cmd),
    .io_out_bits_req_wmask(s2_io_out_bits_req_wmask),
    .io_out_bits_req_wdata(s2_io_out_bits_req_wdata),
    .io_out_bits_metas_0_tag(s2_io_out_bits_metas_0_tag),
    .io_out_bits_metas_0_valid(s2_io_out_bits_metas_0_valid),
    .io_out_bits_metas_0_dirty(s2_io_out_bits_metas_0_dirty),
    .io_out_bits_metas_1_tag(s2_io_out_bits_metas_1_tag),
    .io_out_bits_metas_1_valid(s2_io_out_bits_metas_1_valid),
    .io_out_bits_metas_1_dirty(s2_io_out_bits_metas_1_dirty),
    .io_out_bits_metas_2_tag(s2_io_out_bits_metas_2_tag),
    .io_out_bits_metas_2_valid(s2_io_out_bits_metas_2_valid),
    .io_out_bits_metas_2_dirty(s2_io_out_bits_metas_2_dirty),
    .io_out_bits_metas_3_tag(s2_io_out_bits_metas_3_tag),
    .io_out_bits_metas_3_valid(s2_io_out_bits_metas_3_valid),
    .io_out_bits_metas_3_dirty(s2_io_out_bits_metas_3_dirty),
    .io_out_bits_datas_0_data(s2_io_out_bits_datas_0_data),
    .io_out_bits_datas_1_data(s2_io_out_bits_datas_1_data),
    .io_out_bits_datas_2_data(s2_io_out_bits_datas_2_data),
    .io_out_bits_datas_3_data(s2_io_out_bits_datas_3_data),
    .io_out_bits_hit(s2_io_out_bits_hit),
    .io_out_bits_waymask(s2_io_out_bits_waymask),
    .io_out_bits_mmio(s2_io_out_bits_mmio),
    .io_out_bits_isForwardData(s2_io_out_bits_isForwardData),
    .io_out_bits_forwardData_data_data(s2_io_out_bits_forwardData_data_data),
    .io_out_bits_forwardData_waymask(s2_io_out_bits_forwardData_waymask),
    .io_metaReadResp_0_tag(s2_io_metaReadResp_0_tag),
    .io_metaReadResp_0_valid(s2_io_metaReadResp_0_valid),
    .io_metaReadResp_0_dirty(s2_io_metaReadResp_0_dirty),
    .io_metaReadResp_1_tag(s2_io_metaReadResp_1_tag),
    .io_metaReadResp_1_valid(s2_io_metaReadResp_1_valid),
    .io_metaReadResp_1_dirty(s2_io_metaReadResp_1_dirty),
    .io_metaReadResp_2_tag(s2_io_metaReadResp_2_tag),
    .io_metaReadResp_2_valid(s2_io_metaReadResp_2_valid),
    .io_metaReadResp_2_dirty(s2_io_metaReadResp_2_dirty),
    .io_metaReadResp_3_tag(s2_io_metaReadResp_3_tag),
    .io_metaReadResp_3_valid(s2_io_metaReadResp_3_valid),
    .io_metaReadResp_3_dirty(s2_io_metaReadResp_3_dirty),
    .io_dataReadResp_0_data(s2_io_dataReadResp_0_data),
    .io_dataReadResp_1_data(s2_io_dataReadResp_1_data),
    .io_dataReadResp_2_data(s2_io_dataReadResp_2_data),
    .io_dataReadResp_3_data(s2_io_dataReadResp_3_data),
    .io_metaWriteBus_req_valid(s2_io_metaWriteBus_req_valid),
    .io_metaWriteBus_req_bits_setIdx(s2_io_metaWriteBus_req_bits_setIdx),
    .io_metaWriteBus_req_bits_data_tag(s2_io_metaWriteBus_req_bits_data_tag),
    .io_metaWriteBus_req_bits_data_dirty(s2_io_metaWriteBus_req_bits_data_dirty),
    .io_metaWriteBus_req_bits_waymask(s2_io_metaWriteBus_req_bits_waymask),
    .io_dataWriteBus_req_valid(s2_io_dataWriteBus_req_valid),
    .io_dataWriteBus_req_bits_setIdx(s2_io_dataWriteBus_req_bits_setIdx),
    .io_dataWriteBus_req_bits_data_data(s2_io_dataWriteBus_req_bits_data_data),
    .io_dataWriteBus_req_bits_waymask(s2_io_dataWriteBus_req_bits_waymask),
    .DISPLAY_ENABLE(s2_DISPLAY_ENABLE)
  );
  CacheStage3_1 s3 ( // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
    .clock(s3_clock),
    .reset(s3_reset),
    .io_in_ready(s3_io_in_ready),
    .io_in_valid(s3_io_in_valid),
    .io_in_bits_req_addr(s3_io_in_bits_req_addr),
    .io_in_bits_req_size(s3_io_in_bits_req_size),
    .io_in_bits_req_cmd(s3_io_in_bits_req_cmd),
    .io_in_bits_req_wmask(s3_io_in_bits_req_wmask),
    .io_in_bits_req_wdata(s3_io_in_bits_req_wdata),
    .io_in_bits_metas_0_tag(s3_io_in_bits_metas_0_tag),
    .io_in_bits_metas_0_valid(s3_io_in_bits_metas_0_valid),
    .io_in_bits_metas_0_dirty(s3_io_in_bits_metas_0_dirty),
    .io_in_bits_metas_1_tag(s3_io_in_bits_metas_1_tag),
    .io_in_bits_metas_1_valid(s3_io_in_bits_metas_1_valid),
    .io_in_bits_metas_1_dirty(s3_io_in_bits_metas_1_dirty),
    .io_in_bits_metas_2_tag(s3_io_in_bits_metas_2_tag),
    .io_in_bits_metas_2_valid(s3_io_in_bits_metas_2_valid),
    .io_in_bits_metas_2_dirty(s3_io_in_bits_metas_2_dirty),
    .io_in_bits_metas_3_tag(s3_io_in_bits_metas_3_tag),
    .io_in_bits_metas_3_valid(s3_io_in_bits_metas_3_valid),
    .io_in_bits_metas_3_dirty(s3_io_in_bits_metas_3_dirty),
    .io_in_bits_datas_0_data(s3_io_in_bits_datas_0_data),
    .io_in_bits_datas_1_data(s3_io_in_bits_datas_1_data),
    .io_in_bits_datas_2_data(s3_io_in_bits_datas_2_data),
    .io_in_bits_datas_3_data(s3_io_in_bits_datas_3_data),
    .io_in_bits_hit(s3_io_in_bits_hit),
    .io_in_bits_waymask(s3_io_in_bits_waymask),
    .io_in_bits_mmio(s3_io_in_bits_mmio),
    .io_in_bits_isForwardData(s3_io_in_bits_isForwardData),
    .io_in_bits_forwardData_data_data(s3_io_in_bits_forwardData_data_data),
    .io_in_bits_forwardData_waymask(s3_io_in_bits_forwardData_waymask),
    .io_out_ready(s3_io_out_ready),
    .io_out_valid(s3_io_out_valid),
    .io_out_bits_cmd(s3_io_out_bits_cmd),
    .io_out_bits_rdata(s3_io_out_bits_rdata),
    .io_isFinish(s3_io_isFinish),
    .io_dataReadBus_req_ready(s3_io_dataReadBus_req_ready),
    .io_dataReadBus_req_valid(s3_io_dataReadBus_req_valid),
    .io_dataReadBus_req_bits_setIdx(s3_io_dataReadBus_req_bits_setIdx),
    .io_dataReadBus_resp_data_0_data(s3_io_dataReadBus_resp_data_0_data),
    .io_dataReadBus_resp_data_1_data(s3_io_dataReadBus_resp_data_1_data),
    .io_dataReadBus_resp_data_2_data(s3_io_dataReadBus_resp_data_2_data),
    .io_dataReadBus_resp_data_3_data(s3_io_dataReadBus_resp_data_3_data),
    .io_dataWriteBus_req_valid(s3_io_dataWriteBus_req_valid),
    .io_dataWriteBus_req_bits_setIdx(s3_io_dataWriteBus_req_bits_setIdx),
    .io_dataWriteBus_req_bits_data_data(s3_io_dataWriteBus_req_bits_data_data),
    .io_dataWriteBus_req_bits_waymask(s3_io_dataWriteBus_req_bits_waymask),
    .io_metaWriteBus_req_valid(s3_io_metaWriteBus_req_valid),
    .io_metaWriteBus_req_bits_setIdx(s3_io_metaWriteBus_req_bits_setIdx),
    .io_metaWriteBus_req_bits_data_tag(s3_io_metaWriteBus_req_bits_data_tag),
    .io_metaWriteBus_req_bits_data_valid(s3_io_metaWriteBus_req_bits_data_valid),
    .io_metaWriteBus_req_bits_data_dirty(s3_io_metaWriteBus_req_bits_data_dirty),
    .io_metaWriteBus_req_bits_waymask(s3_io_metaWriteBus_req_bits_waymask),
    .io_mem_req_ready(s3_io_mem_req_ready),
    .io_mem_req_valid(s3_io_mem_req_valid),
    .io_mem_req_bits_addr(s3_io_mem_req_bits_addr),
    .io_mem_req_bits_size(s3_io_mem_req_bits_size),
    .io_mem_req_bits_cmd(s3_io_mem_req_bits_cmd),
    .io_mem_req_bits_wmask(s3_io_mem_req_bits_wmask),
    .io_mem_req_bits_wdata(s3_io_mem_req_bits_wdata),
    .io_mem_resp_ready(s3_io_mem_resp_ready),
    .io_mem_resp_valid(s3_io_mem_resp_valid),
    .io_mem_resp_bits_cmd(s3_io_mem_resp_bits_cmd),
    .io_mem_resp_bits_rdata(s3_io_mem_resp_bits_rdata),
    .io_mmio_req_ready(s3_io_mmio_req_ready),
    .io_mmio_req_valid(s3_io_mmio_req_valid),
    .io_mmio_req_bits_addr(s3_io_mmio_req_bits_addr),
    .io_mmio_req_bits_size(s3_io_mmio_req_bits_size),
    .io_mmio_req_bits_cmd(s3_io_mmio_req_bits_cmd),
    .io_mmio_req_bits_wmask(s3_io_mmio_req_bits_wmask),
    .io_mmio_req_bits_wdata(s3_io_mmio_req_bits_wdata),
    .io_mmio_resp_ready(s3_io_mmio_resp_ready),
    .io_mmio_resp_valid(s3_io_mmio_resp_valid),
    .io_mmio_resp_bits_rdata(s3_io_mmio_resp_bits_rdata),
    .io_cohResp_valid(s3_io_cohResp_valid),
    .io_cohResp_bits_cmd(s3_io_cohResp_bits_cmd),
    .io_cohResp_bits_rdata(s3_io_cohResp_bits_rdata),
    .io_dataReadRespToL1(s3_io_dataReadRespToL1),
    .DISPLAY_ENABLE(s3_DISPLAY_ENABLE),
    ._WIRE_19(s3__WIRE_19)
  );
  SRAMTemplateWithArbiter metaArray ( // @[src/main/scala/nutcore/mem/Cache.scala 483:25]
    .clock(metaArray_clock),
    .reset(metaArray_reset),
    .io_r_0_req_ready(metaArray_io_r_0_req_ready),
    .io_r_0_req_valid(metaArray_io_r_0_req_valid),
    .io_r_0_req_bits_setIdx(metaArray_io_r_0_req_bits_setIdx),
    .io_r_0_resp_data_0_tag(metaArray_io_r_0_resp_data_0_tag),
    .io_r_0_resp_data_0_valid(metaArray_io_r_0_resp_data_0_valid),
    .io_r_0_resp_data_0_dirty(metaArray_io_r_0_resp_data_0_dirty),
    .io_r_0_resp_data_1_tag(metaArray_io_r_0_resp_data_1_tag),
    .io_r_0_resp_data_1_valid(metaArray_io_r_0_resp_data_1_valid),
    .io_r_0_resp_data_1_dirty(metaArray_io_r_0_resp_data_1_dirty),
    .io_r_0_resp_data_2_tag(metaArray_io_r_0_resp_data_2_tag),
    .io_r_0_resp_data_2_valid(metaArray_io_r_0_resp_data_2_valid),
    .io_r_0_resp_data_2_dirty(metaArray_io_r_0_resp_data_2_dirty),
    .io_r_0_resp_data_3_tag(metaArray_io_r_0_resp_data_3_tag),
    .io_r_0_resp_data_3_valid(metaArray_io_r_0_resp_data_3_valid),
    .io_r_0_resp_data_3_dirty(metaArray_io_r_0_resp_data_3_dirty),
    .io_w_req_valid(metaArray_io_w_req_valid),
    .io_w_req_bits_setIdx(metaArray_io_w_req_bits_setIdx),
    .io_w_req_bits_data_tag(metaArray_io_w_req_bits_data_tag),
    .io_w_req_bits_data_dirty(metaArray_io_w_req_bits_data_dirty),
    .io_w_req_bits_waymask(metaArray_io_w_req_bits_waymask)
  );
  SRAMTemplateWithArbiter_1 dataArray ( // @[src/main/scala/nutcore/mem/Cache.scala 484:25]
    .clock(dataArray_clock),
    .reset(dataArray_reset),
    .io_r_0_req_ready(dataArray_io_r_0_req_ready),
    .io_r_0_req_valid(dataArray_io_r_0_req_valid),
    .io_r_0_req_bits_setIdx(dataArray_io_r_0_req_bits_setIdx),
    .io_r_0_resp_data_0_data(dataArray_io_r_0_resp_data_0_data),
    .io_r_0_resp_data_1_data(dataArray_io_r_0_resp_data_1_data),
    .io_r_0_resp_data_2_data(dataArray_io_r_0_resp_data_2_data),
    .io_r_0_resp_data_3_data(dataArray_io_r_0_resp_data_3_data),
    .io_r_1_req_ready(dataArray_io_r_1_req_ready),
    .io_r_1_req_valid(dataArray_io_r_1_req_valid),
    .io_r_1_req_bits_setIdx(dataArray_io_r_1_req_bits_setIdx),
    .io_r_1_resp_data_0_data(dataArray_io_r_1_resp_data_0_data),
    .io_r_1_resp_data_1_data(dataArray_io_r_1_resp_data_1_data),
    .io_r_1_resp_data_2_data(dataArray_io_r_1_resp_data_2_data),
    .io_r_1_resp_data_3_data(dataArray_io_r_1_resp_data_3_data),
    .io_w_req_valid(dataArray_io_w_req_valid),
    .io_w_req_bits_setIdx(dataArray_io_w_req_bits_setIdx),
    .io_w_req_bits_data_data(dataArray_io_w_req_bits_data_data),
    .io_w_req_bits_waymask(dataArray_io_w_req_bits_waymask)
  );
  Arbiter_9 arb ( // @[src/main/scala/nutcore/mem/Cache.scala 493:19]
    .io_in_0_ready(arb_io_in_0_ready),
    .io_in_0_valid(arb_io_in_0_valid),
    .io_in_0_bits_addr(arb_io_in_0_bits_addr),
    .io_in_0_bits_size(arb_io_in_0_bits_size),
    .io_in_0_bits_cmd(arb_io_in_0_bits_cmd),
    .io_in_0_bits_wmask(arb_io_in_0_bits_wmask),
    .io_in_0_bits_wdata(arb_io_in_0_bits_wdata),
    .io_in_1_ready(arb_io_in_1_ready),
    .io_in_1_valid(arb_io_in_1_valid),
    .io_in_1_bits_addr(arb_io_in_1_bits_addr),
    .io_in_1_bits_size(arb_io_in_1_bits_size),
    .io_in_1_bits_cmd(arb_io_in_1_bits_cmd),
    .io_in_1_bits_wmask(arb_io_in_1_bits_wmask),
    .io_in_1_bits_wdata(arb_io_in_1_bits_wdata),
    .io_out_ready(arb_io_out_ready),
    .io_out_valid(arb_io_out_valid),
    .io_out_bits_addr(arb_io_out_bits_addr),
    .io_out_bits_size(arb_io_out_bits_size),
    .io_out_bits_cmd(arb_io_out_bits_cmd),
    .io_out_bits_wmask(arb_io_out_bits_wmask),
    .io_out_bits_wdata(arb_io_out_bits_wdata)
  );
  assign io_in_req_ready = arb_io_in_1_ready; // @[src/main/scala/nutcore/mem/Cache.scala 494:28]
  assign io_in_resp_valid = s3_io_out_valid & _io_in_resp_valid_T ? 1'h0 : s3_io_out_valid | s3_io_dataReadRespToL1; // @[src/main/scala/nutcore/mem/Cache.scala 510:26]
  assign io_in_resp_bits_cmd = s3_io_out_bits_cmd; // @[src/main/scala/nutcore/mem/Cache.scala 504:14]
  assign io_in_resp_bits_rdata = s3_io_out_bits_rdata; // @[src/main/scala/nutcore/mem/Cache.scala 504:14]
  assign io_out_mem_req_valid = s3_io_mem_req_valid; // @[src/main/scala/nutcore/mem/Cache.scala 506:14]
  assign io_out_mem_req_bits_addr = s3_io_mem_req_bits_addr; // @[src/main/scala/nutcore/mem/Cache.scala 506:14]
  assign io_out_mem_req_bits_cmd = s3_io_mem_req_bits_cmd; // @[src/main/scala/nutcore/mem/Cache.scala 506:14]
  assign io_out_mem_req_bits_wdata = s3_io_mem_req_bits_wdata; // @[src/main/scala/nutcore/mem/Cache.scala 506:14]
  assign io_out_coh_req_ready = arb_io_in_0_ready; // @[src/main/scala/nutcore/mem/Cache.scala 519:26]
  assign io_out_coh_resp_valid = s3_io_cohResp_valid; // @[src/main/scala/nutcore/mem/Cache.scala 520:21]
  assign io_out_coh_resp_bits_cmd = s3_io_cohResp_bits_cmd; // @[src/main/scala/nutcore/mem/Cache.scala 520:21]
  assign io_out_coh_resp_bits_rdata = s3_io_cohResp_bits_rdata; // @[src/main/scala/nutcore/mem/Cache.scala 520:21]
  assign io_mmio_req_valid = s3_io_mmio_req_valid; // @[src/main/scala/nutcore/mem/Cache.scala 507:11]
  assign io_mmio_req_bits_addr = s3_io_mmio_req_bits_addr; // @[src/main/scala/nutcore/mem/Cache.scala 507:11]
  assign io_mmio_req_bits_size = s3_io_mmio_req_bits_size; // @[src/main/scala/nutcore/mem/Cache.scala 507:11]
  assign io_mmio_req_bits_cmd = s3_io_mmio_req_bits_cmd; // @[src/main/scala/nutcore/mem/Cache.scala 507:11]
  assign io_mmio_req_bits_wmask = s3_io_mmio_req_bits_wmask; // @[src/main/scala/nutcore/mem/Cache.scala 507:11]
  assign io_mmio_req_bits_wdata = s3_io_mmio_req_bits_wdata; // @[src/main/scala/nutcore/mem/Cache.scala 507:11]
  assign io_empty = ~s2_io_in_valid & ~s3_io_in_valid; // @[src/main/scala/nutcore/mem/Cache.scala 508:31]
  assign _WIRE_17 = s3__WIRE_19;
  assign s1_clock = clock;
  assign s1_reset = reset;
  assign s1_io_in_valid = arb_io_out_valid; // @[src/main/scala/nutcore/mem/Cache.scala 496:12]
  assign s1_io_in_bits_addr = arb_io_out_bits_addr; // @[src/main/scala/nutcore/mem/Cache.scala 496:12]
  assign s1_io_in_bits_size = arb_io_out_bits_size; // @[src/main/scala/nutcore/mem/Cache.scala 496:12]
  assign s1_io_in_bits_cmd = arb_io_out_bits_cmd; // @[src/main/scala/nutcore/mem/Cache.scala 496:12]
  assign s1_io_in_bits_wmask = arb_io_out_bits_wmask; // @[src/main/scala/nutcore/mem/Cache.scala 496:12]
  assign s1_io_in_bits_wdata = arb_io_out_bits_wdata; // @[src/main/scala/nutcore/mem/Cache.scala 496:12]
  assign s1_io_out_ready = s2_io_in_ready; // @[src/main/scala/utils/Pipeline.scala 29:16]
  assign s1_io_metaReadBus_req_ready = metaArray_io_r_0_req_ready; // @[src/main/scala/nutcore/mem/Cache.scala 528:21]
  assign s1_io_metaReadBus_resp_data_0_tag = metaArray_io_r_0_resp_data_0_tag; // @[src/main/scala/nutcore/mem/Cache.scala 528:21]
  assign s1_io_metaReadBus_resp_data_0_valid = metaArray_io_r_0_resp_data_0_valid; // @[src/main/scala/nutcore/mem/Cache.scala 528:21]
  assign s1_io_metaReadBus_resp_data_0_dirty = metaArray_io_r_0_resp_data_0_dirty; // @[src/main/scala/nutcore/mem/Cache.scala 528:21]
  assign s1_io_metaReadBus_resp_data_1_tag = metaArray_io_r_0_resp_data_1_tag; // @[src/main/scala/nutcore/mem/Cache.scala 528:21]
  assign s1_io_metaReadBus_resp_data_1_valid = metaArray_io_r_0_resp_data_1_valid; // @[src/main/scala/nutcore/mem/Cache.scala 528:21]
  assign s1_io_metaReadBus_resp_data_1_dirty = metaArray_io_r_0_resp_data_1_dirty; // @[src/main/scala/nutcore/mem/Cache.scala 528:21]
  assign s1_io_metaReadBus_resp_data_2_tag = metaArray_io_r_0_resp_data_2_tag; // @[src/main/scala/nutcore/mem/Cache.scala 528:21]
  assign s1_io_metaReadBus_resp_data_2_valid = metaArray_io_r_0_resp_data_2_valid; // @[src/main/scala/nutcore/mem/Cache.scala 528:21]
  assign s1_io_metaReadBus_resp_data_2_dirty = metaArray_io_r_0_resp_data_2_dirty; // @[src/main/scala/nutcore/mem/Cache.scala 528:21]
  assign s1_io_metaReadBus_resp_data_3_tag = metaArray_io_r_0_resp_data_3_tag; // @[src/main/scala/nutcore/mem/Cache.scala 528:21]
  assign s1_io_metaReadBus_resp_data_3_valid = metaArray_io_r_0_resp_data_3_valid; // @[src/main/scala/nutcore/mem/Cache.scala 528:21]
  assign s1_io_metaReadBus_resp_data_3_dirty = metaArray_io_r_0_resp_data_3_dirty; // @[src/main/scala/nutcore/mem/Cache.scala 528:21]
  assign s1_io_dataReadBus_req_ready = dataArray_io_r_0_req_ready; // @[src/main/scala/nutcore/mem/Cache.scala 529:21]
  assign s1_io_dataReadBus_resp_data_0_data = dataArray_io_r_0_resp_data_0_data; // @[src/main/scala/nutcore/mem/Cache.scala 529:21]
  assign s1_io_dataReadBus_resp_data_1_data = dataArray_io_r_0_resp_data_1_data; // @[src/main/scala/nutcore/mem/Cache.scala 529:21]
  assign s1_io_dataReadBus_resp_data_2_data = dataArray_io_r_0_resp_data_2_data; // @[src/main/scala/nutcore/mem/Cache.scala 529:21]
  assign s1_io_dataReadBus_resp_data_3_data = dataArray_io_r_0_resp_data_3_data; // @[src/main/scala/nutcore/mem/Cache.scala 529:21]
  assign s1_DISPLAY_ENABLE = DISPLAY_ENABLE;
  assign s2_clock = clock;
  assign s2_reset = reset;
  assign s2_io_in_valid = valid; // @[src/main/scala/utils/Pipeline.scala 31:17]
  assign s2_io_in_bits_req_addr = s2_io_in_bits_r_req_addr; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign s2_io_in_bits_req_size = s2_io_in_bits_r_req_size; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign s2_io_in_bits_req_cmd = s2_io_in_bits_r_req_cmd; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign s2_io_in_bits_req_wmask = s2_io_in_bits_r_req_wmask; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign s2_io_in_bits_req_wdata = s2_io_in_bits_r_req_wdata; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign s2_io_out_ready = s3_io_in_ready; // @[src/main/scala/utils/Pipeline.scala 29:16]
  assign s2_io_metaReadResp_0_tag = s1_io_metaReadBus_resp_data_0_tag; // @[src/main/scala/nutcore/mem/Cache.scala 535:22]
  assign s2_io_metaReadResp_0_valid = s1_io_metaReadBus_resp_data_0_valid; // @[src/main/scala/nutcore/mem/Cache.scala 535:22]
  assign s2_io_metaReadResp_0_dirty = s1_io_metaReadBus_resp_data_0_dirty; // @[src/main/scala/nutcore/mem/Cache.scala 535:22]
  assign s2_io_metaReadResp_1_tag = s1_io_metaReadBus_resp_data_1_tag; // @[src/main/scala/nutcore/mem/Cache.scala 535:22]
  assign s2_io_metaReadResp_1_valid = s1_io_metaReadBus_resp_data_1_valid; // @[src/main/scala/nutcore/mem/Cache.scala 535:22]
  assign s2_io_metaReadResp_1_dirty = s1_io_metaReadBus_resp_data_1_dirty; // @[src/main/scala/nutcore/mem/Cache.scala 535:22]
  assign s2_io_metaReadResp_2_tag = s1_io_metaReadBus_resp_data_2_tag; // @[src/main/scala/nutcore/mem/Cache.scala 535:22]
  assign s2_io_metaReadResp_2_valid = s1_io_metaReadBus_resp_data_2_valid; // @[src/main/scala/nutcore/mem/Cache.scala 535:22]
  assign s2_io_metaReadResp_2_dirty = s1_io_metaReadBus_resp_data_2_dirty; // @[src/main/scala/nutcore/mem/Cache.scala 535:22]
  assign s2_io_metaReadResp_3_tag = s1_io_metaReadBus_resp_data_3_tag; // @[src/main/scala/nutcore/mem/Cache.scala 535:22]
  assign s2_io_metaReadResp_3_valid = s1_io_metaReadBus_resp_data_3_valid; // @[src/main/scala/nutcore/mem/Cache.scala 535:22]
  assign s2_io_metaReadResp_3_dirty = s1_io_metaReadBus_resp_data_3_dirty; // @[src/main/scala/nutcore/mem/Cache.scala 535:22]
  assign s2_io_dataReadResp_0_data = s1_io_dataReadBus_resp_data_0_data; // @[src/main/scala/nutcore/mem/Cache.scala 536:22]
  assign s2_io_dataReadResp_1_data = s1_io_dataReadBus_resp_data_1_data; // @[src/main/scala/nutcore/mem/Cache.scala 536:22]
  assign s2_io_dataReadResp_2_data = s1_io_dataReadBus_resp_data_2_data; // @[src/main/scala/nutcore/mem/Cache.scala 536:22]
  assign s2_io_dataReadResp_3_data = s1_io_dataReadBus_resp_data_3_data; // @[src/main/scala/nutcore/mem/Cache.scala 536:22]
  assign s2_io_metaWriteBus_req_valid = s3_io_metaWriteBus_req_valid; // @[src/main/scala/nutcore/mem/Cache.scala 538:22]
  assign s2_io_metaWriteBus_req_bits_setIdx = s3_io_metaWriteBus_req_bits_setIdx; // @[src/main/scala/nutcore/mem/Cache.scala 538:22]
  assign s2_io_metaWriteBus_req_bits_data_tag = s3_io_metaWriteBus_req_bits_data_tag; // @[src/main/scala/nutcore/mem/Cache.scala 538:22]
  assign s2_io_metaWriteBus_req_bits_data_dirty = s3_io_metaWriteBus_req_bits_data_dirty; // @[src/main/scala/nutcore/mem/Cache.scala 538:22]
  assign s2_io_metaWriteBus_req_bits_waymask = s3_io_metaWriteBus_req_bits_waymask; // @[src/main/scala/nutcore/mem/Cache.scala 538:22]
  assign s2_io_dataWriteBus_req_valid = s3_io_dataWriteBus_req_valid; // @[src/main/scala/nutcore/mem/Cache.scala 537:22]
  assign s2_io_dataWriteBus_req_bits_setIdx = s3_io_dataWriteBus_req_bits_setIdx; // @[src/main/scala/nutcore/mem/Cache.scala 537:22]
  assign s2_io_dataWriteBus_req_bits_data_data = s3_io_dataWriteBus_req_bits_data_data; // @[src/main/scala/nutcore/mem/Cache.scala 537:22]
  assign s2_io_dataWriteBus_req_bits_waymask = s3_io_dataWriteBus_req_bits_waymask; // @[src/main/scala/nutcore/mem/Cache.scala 537:22]
  assign s2_DISPLAY_ENABLE = DISPLAY_ENABLE;
  assign s3_clock = clock;
  assign s3_reset = reset;
  assign s3_io_in_valid = valid_1; // @[src/main/scala/utils/Pipeline.scala 31:17]
  assign s3_io_in_bits_req_addr = s3_io_in_bits_r_req_addr; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign s3_io_in_bits_req_size = s3_io_in_bits_r_req_size; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign s3_io_in_bits_req_cmd = s3_io_in_bits_r_req_cmd; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign s3_io_in_bits_req_wmask = s3_io_in_bits_r_req_wmask; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign s3_io_in_bits_req_wdata = s3_io_in_bits_r_req_wdata; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign s3_io_in_bits_metas_0_tag = s3_io_in_bits_r_metas_0_tag; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign s3_io_in_bits_metas_0_valid = s3_io_in_bits_r_metas_0_valid; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign s3_io_in_bits_metas_0_dirty = s3_io_in_bits_r_metas_0_dirty; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign s3_io_in_bits_metas_1_tag = s3_io_in_bits_r_metas_1_tag; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign s3_io_in_bits_metas_1_valid = s3_io_in_bits_r_metas_1_valid; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign s3_io_in_bits_metas_1_dirty = s3_io_in_bits_r_metas_1_dirty; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign s3_io_in_bits_metas_2_tag = s3_io_in_bits_r_metas_2_tag; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign s3_io_in_bits_metas_2_valid = s3_io_in_bits_r_metas_2_valid; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign s3_io_in_bits_metas_2_dirty = s3_io_in_bits_r_metas_2_dirty; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign s3_io_in_bits_metas_3_tag = s3_io_in_bits_r_metas_3_tag; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign s3_io_in_bits_metas_3_valid = s3_io_in_bits_r_metas_3_valid; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign s3_io_in_bits_metas_3_dirty = s3_io_in_bits_r_metas_3_dirty; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign s3_io_in_bits_datas_0_data = s3_io_in_bits_r_datas_0_data; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign s3_io_in_bits_datas_1_data = s3_io_in_bits_r_datas_1_data; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign s3_io_in_bits_datas_2_data = s3_io_in_bits_r_datas_2_data; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign s3_io_in_bits_datas_3_data = s3_io_in_bits_r_datas_3_data; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign s3_io_in_bits_hit = s3_io_in_bits_r_hit; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign s3_io_in_bits_waymask = s3_io_in_bits_r_waymask; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign s3_io_in_bits_mmio = s3_io_in_bits_r_mmio; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign s3_io_in_bits_isForwardData = s3_io_in_bits_r_isForwardData; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign s3_io_in_bits_forwardData_data_data = s3_io_in_bits_r_forwardData_data_data; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign s3_io_in_bits_forwardData_waymask = s3_io_in_bits_r_forwardData_waymask; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign s3_io_out_ready = io_in_resp_ready; // @[src/main/scala/nutcore/mem/Cache.scala 504:14]
  assign s3_io_dataReadBus_req_ready = dataArray_io_r_1_req_ready; // @[src/main/scala/nutcore/mem/Cache.scala 530:21]
  assign s3_io_dataReadBus_resp_data_0_data = dataArray_io_r_1_resp_data_0_data; // @[src/main/scala/nutcore/mem/Cache.scala 530:21]
  assign s3_io_dataReadBus_resp_data_1_data = dataArray_io_r_1_resp_data_1_data; // @[src/main/scala/nutcore/mem/Cache.scala 530:21]
  assign s3_io_dataReadBus_resp_data_2_data = dataArray_io_r_1_resp_data_2_data; // @[src/main/scala/nutcore/mem/Cache.scala 530:21]
  assign s3_io_dataReadBus_resp_data_3_data = dataArray_io_r_1_resp_data_3_data; // @[src/main/scala/nutcore/mem/Cache.scala 530:21]
  assign s3_io_mem_req_ready = io_out_mem_req_ready; // @[src/main/scala/nutcore/mem/Cache.scala 506:14]
  assign s3_io_mem_resp_valid = io_out_mem_resp_valid; // @[src/main/scala/nutcore/mem/Cache.scala 506:14]
  assign s3_io_mem_resp_bits_cmd = io_out_mem_resp_bits_cmd; // @[src/main/scala/nutcore/mem/Cache.scala 506:14]
  assign s3_io_mem_resp_bits_rdata = io_out_mem_resp_bits_rdata; // @[src/main/scala/nutcore/mem/Cache.scala 506:14]
  assign s3_io_mmio_req_ready = io_mmio_req_ready; // @[src/main/scala/nutcore/mem/Cache.scala 507:11]
  assign s3_io_mmio_resp_valid = io_mmio_resp_valid; // @[src/main/scala/nutcore/mem/Cache.scala 507:11]
  assign s3_io_mmio_resp_bits_rdata = io_mmio_resp_bits_rdata; // @[src/main/scala/nutcore/mem/Cache.scala 507:11]
  assign s3_DISPLAY_ENABLE = DISPLAY_ENABLE;
  assign metaArray_clock = clock;
  assign metaArray_reset = reset;
  assign metaArray_io_r_0_req_valid = s1_io_metaReadBus_req_valid; // @[src/main/scala/nutcore/mem/Cache.scala 528:21]
  assign metaArray_io_r_0_req_bits_setIdx = s1_io_metaReadBus_req_bits_setIdx; // @[src/main/scala/nutcore/mem/Cache.scala 528:21]
  assign metaArray_io_w_req_valid = s3_io_metaWriteBus_req_valid; // @[src/main/scala/nutcore/mem/Cache.scala 532:18]
  assign metaArray_io_w_req_bits_setIdx = s3_io_metaWriteBus_req_bits_setIdx; // @[src/main/scala/nutcore/mem/Cache.scala 532:18]
  assign metaArray_io_w_req_bits_data_tag = s3_io_metaWriteBus_req_bits_data_tag; // @[src/main/scala/nutcore/mem/Cache.scala 532:18]
  assign metaArray_io_w_req_bits_data_dirty = s3_io_metaWriteBus_req_bits_data_dirty; // @[src/main/scala/nutcore/mem/Cache.scala 532:18]
  assign metaArray_io_w_req_bits_waymask = s3_io_metaWriteBus_req_bits_waymask; // @[src/main/scala/nutcore/mem/Cache.scala 532:18]
  assign dataArray_clock = clock;
  assign dataArray_reset = reset;
  assign dataArray_io_r_0_req_valid = s1_io_dataReadBus_req_valid; // @[src/main/scala/nutcore/mem/Cache.scala 529:21]
  assign dataArray_io_r_0_req_bits_setIdx = s1_io_dataReadBus_req_bits_setIdx; // @[src/main/scala/nutcore/mem/Cache.scala 529:21]
  assign dataArray_io_r_1_req_valid = s3_io_dataReadBus_req_valid; // @[src/main/scala/nutcore/mem/Cache.scala 530:21]
  assign dataArray_io_r_1_req_bits_setIdx = s3_io_dataReadBus_req_bits_setIdx; // @[src/main/scala/nutcore/mem/Cache.scala 530:21]
  assign dataArray_io_w_req_valid = s3_io_dataWriteBus_req_valid; // @[src/main/scala/nutcore/mem/Cache.scala 533:18]
  assign dataArray_io_w_req_bits_setIdx = s3_io_dataWriteBus_req_bits_setIdx; // @[src/main/scala/nutcore/mem/Cache.scala 533:18]
  assign dataArray_io_w_req_bits_data_data = s3_io_dataWriteBus_req_bits_data_data; // @[src/main/scala/nutcore/mem/Cache.scala 533:18]
  assign dataArray_io_w_req_bits_waymask = s3_io_dataWriteBus_req_bits_waymask; // @[src/main/scala/nutcore/mem/Cache.scala 533:18]
  assign arb_io_in_0_valid = io_out_coh_req_valid; // @[src/main/scala/nutcore/mem/Cache.scala 518:24]
  assign arb_io_in_0_bits_addr = io_out_coh_req_bits_addr; // @[src/main/scala/nutcore/mem/Cache.scala 515:19 src/main/scala/bus/simplebus/SimpleBus.scala 64:15]
  assign arb_io_in_0_bits_size = 3'h3; // @[src/main/scala/nutcore/mem/Cache.scala 515:19 src/main/scala/bus/simplebus/SimpleBus.scala 66:15]
  assign arb_io_in_0_bits_cmd = 4'h8; // @[src/main/scala/nutcore/mem/Cache.scala 515:19 src/main/scala/bus/simplebus/SimpleBus.scala 65:14]
  assign arb_io_in_0_bits_wmask = 8'hff; // @[src/main/scala/nutcore/mem/Cache.scala 515:19 src/main/scala/bus/simplebus/SimpleBus.scala 68:16]
  assign arb_io_in_0_bits_wdata = io_out_coh_req_bits_wdata; // @[src/main/scala/nutcore/mem/Cache.scala 515:19 src/main/scala/bus/simplebus/SimpleBus.scala 67:16]
  assign arb_io_in_1_valid = io_in_req_valid; // @[src/main/scala/nutcore/mem/Cache.scala 494:28]
  assign arb_io_in_1_bits_addr = io_in_req_bits_addr; // @[src/main/scala/nutcore/mem/Cache.scala 494:28]
  assign arb_io_in_1_bits_size = io_in_req_bits_size; // @[src/main/scala/nutcore/mem/Cache.scala 494:28]
  assign arb_io_in_1_bits_cmd = io_in_req_bits_cmd; // @[src/main/scala/nutcore/mem/Cache.scala 494:28]
  assign arb_io_in_1_bits_wmask = io_in_req_bits_wmask; // @[src/main/scala/nutcore/mem/Cache.scala 494:28]
  assign arb_io_in_1_bits_wdata = io_in_req_bits_wdata; // @[src/main/scala/nutcore/mem/Cache.scala 494:28]
  assign arb_io_out_ready = s1_io_in_ready; // @[src/main/scala/nutcore/mem/Cache.scala 496:12]
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/utils/Pipeline.scala 24:24]
      valid <= 1'h0; // @[src/main/scala/utils/Pipeline.scala 24:24]
    end else begin
      valid <= _GEN_1;
    end
    if (_T_2) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      s2_io_in_bits_r_req_addr <= s1_io_out_bits_req_addr; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_2) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      s2_io_in_bits_r_req_size <= s1_io_out_bits_req_size; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_2) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      s2_io_in_bits_r_req_cmd <= s1_io_out_bits_req_cmd; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_2) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      s2_io_in_bits_r_req_wmask <= s1_io_out_bits_req_wmask; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_2) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      s2_io_in_bits_r_req_wdata <= s1_io_out_bits_req_wdata; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (reset) begin // @[src/main/scala/utils/Pipeline.scala 24:24]
      valid_1 <= 1'h0; // @[src/main/scala/utils/Pipeline.scala 24:24]
    end else begin
      valid_1 <= _GEN_9;
    end
    if (_T_4) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      s3_io_in_bits_r_req_addr <= s2_io_out_bits_req_addr; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_4) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      s3_io_in_bits_r_req_size <= s2_io_out_bits_req_size; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_4) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      s3_io_in_bits_r_req_cmd <= s2_io_out_bits_req_cmd; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_4) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      s3_io_in_bits_r_req_wmask <= s2_io_out_bits_req_wmask; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_4) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      s3_io_in_bits_r_req_wdata <= s2_io_out_bits_req_wdata; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_4) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      s3_io_in_bits_r_metas_0_tag <= s2_io_out_bits_metas_0_tag; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_4) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      s3_io_in_bits_r_metas_0_valid <= s2_io_out_bits_metas_0_valid; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_4) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      s3_io_in_bits_r_metas_0_dirty <= s2_io_out_bits_metas_0_dirty; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_4) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      s3_io_in_bits_r_metas_1_tag <= s2_io_out_bits_metas_1_tag; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_4) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      s3_io_in_bits_r_metas_1_valid <= s2_io_out_bits_metas_1_valid; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_4) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      s3_io_in_bits_r_metas_1_dirty <= s2_io_out_bits_metas_1_dirty; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_4) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      s3_io_in_bits_r_metas_2_tag <= s2_io_out_bits_metas_2_tag; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_4) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      s3_io_in_bits_r_metas_2_valid <= s2_io_out_bits_metas_2_valid; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_4) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      s3_io_in_bits_r_metas_2_dirty <= s2_io_out_bits_metas_2_dirty; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_4) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      s3_io_in_bits_r_metas_3_tag <= s2_io_out_bits_metas_3_tag; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_4) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      s3_io_in_bits_r_metas_3_valid <= s2_io_out_bits_metas_3_valid; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_4) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      s3_io_in_bits_r_metas_3_dirty <= s2_io_out_bits_metas_3_dirty; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_4) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      s3_io_in_bits_r_datas_0_data <= s2_io_out_bits_datas_0_data; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_4) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      s3_io_in_bits_r_datas_1_data <= s2_io_out_bits_datas_1_data; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_4) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      s3_io_in_bits_r_datas_2_data <= s2_io_out_bits_datas_2_data; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_4) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      s3_io_in_bits_r_datas_3_data <= s2_io_out_bits_datas_3_data; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_4) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      s3_io_in_bits_r_hit <= s2_io_out_bits_hit; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_4) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      s3_io_in_bits_r_waymask <= s2_io_out_bits_waymask; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_4) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      s3_io_in_bits_r_mmio <= s2_io_out_bits_mmio; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_4) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      s3_io_in_bits_r_isForwardData <= s2_io_out_bits_isForwardData; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_4) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      s3_io_in_bits_r_forwardData_data_data <= s2_io_out_bits_forwardData_data_data; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_4) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      s3_io_in_bits_r_forwardData_waymask <= s2_io_out_bits_forwardData_waymask; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (reset) begin // @[src/main/scala/utils/GTimer.scala 24:20]
      c <= 64'h0; // @[src/main/scala/utils/GTimer.scala 24:20]
    end else begin
      c <= _c_T_1; // @[src/main/scala/utils/GTimer.scala 25:7]
    end
    if (reset) begin // @[src/main/scala/utils/GTimer.scala 24:20]
      c_1 <= 64'h0; // @[src/main/scala/utils/GTimer.scala 24:20]
    end else begin
      c_1 <= _c_T_3; // @[src/main/scala/utils/GTimer.scala 25:7]
    end
    if (reset) begin // @[src/main/scala/utils/GTimer.scala 24:20]
      c_2 <= 64'h0; // @[src/main/scala/utils/GTimer.scala 24:20]
    end else begin
      c_2 <= _c_T_5; // @[src/main/scala/utils/GTimer.scala 25:7]
    end
    if (reset) begin // @[src/main/scala/utils/GTimer.scala 24:20]
      c_3 <= 64'h0; // @[src/main/scala/utils/GTimer.scala 24:20]
    end else begin
      c_3 <= _c_T_7; // @[src/main/scala/utils/GTimer.scala 25:7]
    end
    if (reset) begin // @[src/main/scala/utils/GTimer.scala 24:20]
      c_4 <= 64'h0; // @[src/main/scala/utils/GTimer.scala 24:20]
    end else begin
      c_4 <= _c_T_9; // @[src/main/scala/utils/GTimer.scala 25:7]
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & ~reset) begin
          $fwrite(32'h80000002,"[%d] Cache_1: ",c); // @[src/main/scala/utils/Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_7) begin
          $fwrite(32'h80000002,"InReq(%d, %d) InResp(%d, %d) \n",io_in_req_valid,io_in_req_ready,io_in_resp_valid,
            io_in_resp_ready); // @[src/main/scala/utils/Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & ~reset) begin
          $fwrite(32'h80000002,"[%d] Cache_1: ",c_1); // @[src/main/scala/utils/Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_7) begin
          $fwrite(32'h80000002,"{IN s1:(%d,%d), s2:(%d,%d), s3:(%d,%d)} {OUT s1:(%d,%d), s2:(%d,%d), s3:(%d,%d)}\n",
            s1_io_in_valid,s1_io_in_ready,s2_io_in_valid,s2_io_in_ready,s3_io_in_valid,s3_io_in_ready,s1_io_out_valid,
            s1_io_out_ready,s2_io_out_valid,s2_io_out_ready,s3_io_out_valid,s3_io_out_ready); // @[src/main/scala/utils/Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (s1_io_in_valid & DISPLAY_ENABLE & ~reset) begin
          $fwrite(32'h80000002,"[%d] Cache_1: ",c_2); // @[src/main/scala/utils/Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_39 & _T_7) begin
          $fwrite(32'h80000002,"[dcache.S1]: addr = 0x%x, cmd = %d, size = %d, wmask = 0x%x, wdata = 0x%x\n",
            s1_io_in_bits_addr,s1_io_in_bits_cmd,s1_io_in_bits_size,s1_io_in_bits_wmask,s1_io_in_bits_wdata); // @[src/main/scala/utils/Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (s2_io_in_valid & DISPLAY_ENABLE & ~reset) begin
          $fwrite(32'h80000002,"[%d] Cache_1: ",c_3); // @[src/main/scala/utils/Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_41 & _T_7) begin
          $fwrite(32'h80000002,"[dcache.S2]: addr = 0x%x, cmd = %d, size = %d, wmask = 0x%x, wdata = 0x%x\n",
            s2_io_in_bits_req_addr,s2_io_in_bits_req_cmd,s2_io_in_bits_req_size,s2_io_in_bits_req_wmask,
            s2_io_in_bits_req_wdata); // @[src/main/scala/utils/Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (s3_io_in_valid & DISPLAY_ENABLE & ~reset) begin
          $fwrite(32'h80000002,"[%d] Cache_1: ",c_4); // @[src/main/scala/utils/Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_43 & _T_7) begin
          $fwrite(32'h80000002,"[dcache.S3]: addr = 0x%x, cmd = %d, size = %d, wmask = 0x%x, wdata = 0x%x\n",
            s3_io_in_bits_req_addr,s3_io_in_bits_req_cmd,s3_io_in_bits_req_size,s3_io_in_bits_req_wmask,
            s3_io_in_bits_req_wdata); // @[src/main/scala/utils/Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  valid = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  s2_io_in_bits_r_req_addr = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  s2_io_in_bits_r_req_size = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  s2_io_in_bits_r_req_cmd = _RAND_3[3:0];
  _RAND_4 = {1{`RANDOM}};
  s2_io_in_bits_r_req_wmask = _RAND_4[7:0];
  _RAND_5 = {2{`RANDOM}};
  s2_io_in_bits_r_req_wdata = _RAND_5[63:0];
  _RAND_6 = {1{`RANDOM}};
  valid_1 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  s3_io_in_bits_r_req_addr = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  s3_io_in_bits_r_req_size = _RAND_8[2:0];
  _RAND_9 = {1{`RANDOM}};
  s3_io_in_bits_r_req_cmd = _RAND_9[3:0];
  _RAND_10 = {1{`RANDOM}};
  s3_io_in_bits_r_req_wmask = _RAND_10[7:0];
  _RAND_11 = {2{`RANDOM}};
  s3_io_in_bits_r_req_wdata = _RAND_11[63:0];
  _RAND_12 = {1{`RANDOM}};
  s3_io_in_bits_r_metas_0_tag = _RAND_12[18:0];
  _RAND_13 = {1{`RANDOM}};
  s3_io_in_bits_r_metas_0_valid = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  s3_io_in_bits_r_metas_0_dirty = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  s3_io_in_bits_r_metas_1_tag = _RAND_15[18:0];
  _RAND_16 = {1{`RANDOM}};
  s3_io_in_bits_r_metas_1_valid = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  s3_io_in_bits_r_metas_1_dirty = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  s3_io_in_bits_r_metas_2_tag = _RAND_18[18:0];
  _RAND_19 = {1{`RANDOM}};
  s3_io_in_bits_r_metas_2_valid = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  s3_io_in_bits_r_metas_2_dirty = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  s3_io_in_bits_r_metas_3_tag = _RAND_21[18:0];
  _RAND_22 = {1{`RANDOM}};
  s3_io_in_bits_r_metas_3_valid = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  s3_io_in_bits_r_metas_3_dirty = _RAND_23[0:0];
  _RAND_24 = {2{`RANDOM}};
  s3_io_in_bits_r_datas_0_data = _RAND_24[63:0];
  _RAND_25 = {2{`RANDOM}};
  s3_io_in_bits_r_datas_1_data = _RAND_25[63:0];
  _RAND_26 = {2{`RANDOM}};
  s3_io_in_bits_r_datas_2_data = _RAND_26[63:0];
  _RAND_27 = {2{`RANDOM}};
  s3_io_in_bits_r_datas_3_data = _RAND_27[63:0];
  _RAND_28 = {1{`RANDOM}};
  s3_io_in_bits_r_hit = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  s3_io_in_bits_r_waymask = _RAND_29[3:0];
  _RAND_30 = {1{`RANDOM}};
  s3_io_in_bits_r_mmio = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  s3_io_in_bits_r_isForwardData = _RAND_31[0:0];
  _RAND_32 = {2{`RANDOM}};
  s3_io_in_bits_r_forwardData_data_data = _RAND_32[63:0];
  _RAND_33 = {1{`RANDOM}};
  s3_io_in_bits_r_forwardData_waymask = _RAND_33[3:0];
  _RAND_34 = {2{`RANDOM}};
  c = _RAND_34[63:0];
  _RAND_35 = {2{`RANDOM}};
  c_1 = _RAND_35[63:0];
  _RAND_36 = {2{`RANDOM}};
  c_2 = _RAND_36[63:0];
  _RAND_37 = {2{`RANDOM}};
  c_3 = _RAND_37[63:0];
  _RAND_38 = {2{`RANDOM}};
  c_4 = _RAND_38[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module NutCore(
  input         clock,
  input         reset,
  input         io_imem_mem_req_ready, // @[src/main/scala/nutcore/NutCore.scala 98:14]
  output        io_imem_mem_req_valid, // @[src/main/scala/nutcore/NutCore.scala 98:14]
  output [31:0] io_imem_mem_req_bits_addr, // @[src/main/scala/nutcore/NutCore.scala 98:14]
  output [3:0]  io_imem_mem_req_bits_cmd, // @[src/main/scala/nutcore/NutCore.scala 98:14]
  output [63:0] io_imem_mem_req_bits_wdata, // @[src/main/scala/nutcore/NutCore.scala 98:14]
  input         io_imem_mem_resp_valid, // @[src/main/scala/nutcore/NutCore.scala 98:14]
  input  [3:0]  io_imem_mem_resp_bits_cmd, // @[src/main/scala/nutcore/NutCore.scala 98:14]
  input  [63:0] io_imem_mem_resp_bits_rdata, // @[src/main/scala/nutcore/NutCore.scala 98:14]
  input         io_dmem_mem_req_ready, // @[src/main/scala/nutcore/NutCore.scala 98:14]
  output        io_dmem_mem_req_valid, // @[src/main/scala/nutcore/NutCore.scala 98:14]
  output [31:0] io_dmem_mem_req_bits_addr, // @[src/main/scala/nutcore/NutCore.scala 98:14]
  output [3:0]  io_dmem_mem_req_bits_cmd, // @[src/main/scala/nutcore/NutCore.scala 98:14]
  output [63:0] io_dmem_mem_req_bits_wdata, // @[src/main/scala/nutcore/NutCore.scala 98:14]
  input         io_dmem_mem_resp_valid, // @[src/main/scala/nutcore/NutCore.scala 98:14]
  input  [3:0]  io_dmem_mem_resp_bits_cmd, // @[src/main/scala/nutcore/NutCore.scala 98:14]
  input  [63:0] io_dmem_mem_resp_bits_rdata, // @[src/main/scala/nutcore/NutCore.scala 98:14]
  output        io_dmem_coh_req_ready, // @[src/main/scala/nutcore/NutCore.scala 98:14]
  input         io_dmem_coh_req_valid, // @[src/main/scala/nutcore/NutCore.scala 98:14]
  input  [31:0] io_dmem_coh_req_bits_addr, // @[src/main/scala/nutcore/NutCore.scala 98:14]
  input  [63:0] io_dmem_coh_req_bits_wdata, // @[src/main/scala/nutcore/NutCore.scala 98:14]
  output        io_dmem_coh_resp_valid, // @[src/main/scala/nutcore/NutCore.scala 98:14]
  output [3:0]  io_dmem_coh_resp_bits_cmd, // @[src/main/scala/nutcore/NutCore.scala 98:14]
  output [63:0] io_dmem_coh_resp_bits_rdata, // @[src/main/scala/nutcore/NutCore.scala 98:14]
  input         io_mmio_req_ready, // @[src/main/scala/nutcore/NutCore.scala 98:14]
  output        io_mmio_req_valid, // @[src/main/scala/nutcore/NutCore.scala 98:14]
  output [31:0] io_mmio_req_bits_addr, // @[src/main/scala/nutcore/NutCore.scala 98:14]
  output [2:0]  io_mmio_req_bits_size, // @[src/main/scala/nutcore/NutCore.scala 98:14]
  output [3:0]  io_mmio_req_bits_cmd, // @[src/main/scala/nutcore/NutCore.scala 98:14]
  output [7:0]  io_mmio_req_bits_wmask, // @[src/main/scala/nutcore/NutCore.scala 98:14]
  output [63:0] io_mmio_req_bits_wdata, // @[src/main/scala/nutcore/NutCore.scala 98:14]
  input         io_mmio_resp_valid, // @[src/main/scala/nutcore/NutCore.scala 98:14]
  input  [3:0]  io_mmio_resp_bits_cmd, // @[src/main/scala/nutcore/NutCore.scala 98:14]
  input  [63:0] io_mmio_resp_bits_rdata, // @[src/main/scala/nutcore/NutCore.scala 98:14]
  output        io_frontend_req_ready, // @[src/main/scala/nutcore/NutCore.scala 98:14]
  input         io_frontend_req_valid, // @[src/main/scala/nutcore/NutCore.scala 98:14]
  input  [31:0] io_frontend_req_bits_addr, // @[src/main/scala/nutcore/NutCore.scala 98:14]
  input  [2:0]  io_frontend_req_bits_size, // @[src/main/scala/nutcore/NutCore.scala 98:14]
  input  [3:0]  io_frontend_req_bits_cmd, // @[src/main/scala/nutcore/NutCore.scala 98:14]
  input  [7:0]  io_frontend_req_bits_wmask, // @[src/main/scala/nutcore/NutCore.scala 98:14]
  input  [63:0] io_frontend_req_bits_wdata, // @[src/main/scala/nutcore/NutCore.scala 98:14]
  input         io_frontend_resp_ready, // @[src/main/scala/nutcore/NutCore.scala 98:14]
  output        io_frontend_resp_valid, // @[src/main/scala/nutcore/NutCore.scala 98:14]
  output [3:0]  io_frontend_resp_bits_cmd, // @[src/main/scala/nutcore/NutCore.scala 98:14]
  output [63:0] io_frontend_resp_bits_rdata, // @[src/main/scala/nutcore/NutCore.scala 98:14]
  input         io_extra_meip_0,
  output        _WIRE_0,
  input         DISPLAY_ENABLE,
  input         io_extra_mtip,
  input         io_extra_msip
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [63:0] _RAND_29;
  reg [63:0] _RAND_30;
  reg [63:0] _RAND_31;
  reg [63:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [63:0] _RAND_59;
  reg [63:0] _RAND_60;
  reg [63:0] _RAND_61;
  reg [63:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [63:0] _RAND_89;
  reg [63:0] _RAND_90;
  reg [63:0] _RAND_91;
  reg [63:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [63:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [63:0] _RAND_122;
`endif // RANDOMIZE_REG_INIT
  wire  frontend_clock; // @[src/main/scala/nutcore/NutCore.scala 104:34]
  wire  frontend_reset; // @[src/main/scala/nutcore/NutCore.scala 104:34]
  wire  frontend_io_imem_req_ready; // @[src/main/scala/nutcore/NutCore.scala 104:34]
  wire  frontend_io_imem_req_valid; // @[src/main/scala/nutcore/NutCore.scala 104:34]
  wire [38:0] frontend_io_imem_req_bits_addr; // @[src/main/scala/nutcore/NutCore.scala 104:34]
  wire [86:0] frontend_io_imem_req_bits_user; // @[src/main/scala/nutcore/NutCore.scala 104:34]
  wire  frontend_io_imem_resp_ready; // @[src/main/scala/nutcore/NutCore.scala 104:34]
  wire  frontend_io_imem_resp_valid; // @[src/main/scala/nutcore/NutCore.scala 104:34]
  wire [63:0] frontend_io_imem_resp_bits_rdata; // @[src/main/scala/nutcore/NutCore.scala 104:34]
  wire [86:0] frontend_io_imem_resp_bits_user; // @[src/main/scala/nutcore/NutCore.scala 104:34]
  wire  frontend_io_out_0_ready; // @[src/main/scala/nutcore/NutCore.scala 104:34]
  wire  frontend_io_out_0_valid; // @[src/main/scala/nutcore/NutCore.scala 104:34]
  wire [63:0] frontend_io_out_0_bits_cf_instr; // @[src/main/scala/nutcore/NutCore.scala 104:34]
  wire [38:0] frontend_io_out_0_bits_cf_pc; // @[src/main/scala/nutcore/NutCore.scala 104:34]
  wire [38:0] frontend_io_out_0_bits_cf_pnpc; // @[src/main/scala/nutcore/NutCore.scala 104:34]
  wire  frontend_io_out_0_bits_cf_exceptionVec_1; // @[src/main/scala/nutcore/NutCore.scala 104:34]
  wire  frontend_io_out_0_bits_cf_exceptionVec_2; // @[src/main/scala/nutcore/NutCore.scala 104:34]
  wire  frontend_io_out_0_bits_cf_exceptionVec_12; // @[src/main/scala/nutcore/NutCore.scala 104:34]
  wire  frontend_io_out_0_bits_cf_intrVec_0; // @[src/main/scala/nutcore/NutCore.scala 104:34]
  wire  frontend_io_out_0_bits_cf_intrVec_1; // @[src/main/scala/nutcore/NutCore.scala 104:34]
  wire  frontend_io_out_0_bits_cf_intrVec_2; // @[src/main/scala/nutcore/NutCore.scala 104:34]
  wire  frontend_io_out_0_bits_cf_intrVec_3; // @[src/main/scala/nutcore/NutCore.scala 104:34]
  wire  frontend_io_out_0_bits_cf_intrVec_4; // @[src/main/scala/nutcore/NutCore.scala 104:34]
  wire  frontend_io_out_0_bits_cf_intrVec_5; // @[src/main/scala/nutcore/NutCore.scala 104:34]
  wire  frontend_io_out_0_bits_cf_intrVec_6; // @[src/main/scala/nutcore/NutCore.scala 104:34]
  wire  frontend_io_out_0_bits_cf_intrVec_7; // @[src/main/scala/nutcore/NutCore.scala 104:34]
  wire  frontend_io_out_0_bits_cf_intrVec_8; // @[src/main/scala/nutcore/NutCore.scala 104:34]
  wire  frontend_io_out_0_bits_cf_intrVec_9; // @[src/main/scala/nutcore/NutCore.scala 104:34]
  wire  frontend_io_out_0_bits_cf_intrVec_10; // @[src/main/scala/nutcore/NutCore.scala 104:34]
  wire  frontend_io_out_0_bits_cf_intrVec_11; // @[src/main/scala/nutcore/NutCore.scala 104:34]
  wire [3:0] frontend_io_out_0_bits_cf_brIdx; // @[src/main/scala/nutcore/NutCore.scala 104:34]
  wire  frontend_io_out_0_bits_cf_crossPageIPFFix; // @[src/main/scala/nutcore/NutCore.scala 104:34]
  wire  frontend_io_out_0_bits_ctrl_src1Type; // @[src/main/scala/nutcore/NutCore.scala 104:34]
  wire  frontend_io_out_0_bits_ctrl_src2Type; // @[src/main/scala/nutcore/NutCore.scala 104:34]
  wire [2:0] frontend_io_out_0_bits_ctrl_fuType; // @[src/main/scala/nutcore/NutCore.scala 104:34]
  wire [6:0] frontend_io_out_0_bits_ctrl_fuOpType; // @[src/main/scala/nutcore/NutCore.scala 104:34]
  wire [4:0] frontend_io_out_0_bits_ctrl_rfSrc1; // @[src/main/scala/nutcore/NutCore.scala 104:34]
  wire [4:0] frontend_io_out_0_bits_ctrl_rfSrc2; // @[src/main/scala/nutcore/NutCore.scala 104:34]
  wire  frontend_io_out_0_bits_ctrl_rfWen; // @[src/main/scala/nutcore/NutCore.scala 104:34]
  wire [4:0] frontend_io_out_0_bits_ctrl_rfDest; // @[src/main/scala/nutcore/NutCore.scala 104:34]
  wire  frontend_io_out_0_bits_ctrl_isNutCoreTrap; // @[src/main/scala/nutcore/NutCore.scala 104:34]
  wire [63:0] frontend_io_out_0_bits_data_imm; // @[src/main/scala/nutcore/NutCore.scala 104:34]
  wire  frontend_io_out_1_bits_cf_intrVec_0; // @[src/main/scala/nutcore/NutCore.scala 104:34]
  wire  frontend_io_out_1_bits_cf_intrVec_1; // @[src/main/scala/nutcore/NutCore.scala 104:34]
  wire  frontend_io_out_1_bits_cf_intrVec_2; // @[src/main/scala/nutcore/NutCore.scala 104:34]
  wire  frontend_io_out_1_bits_cf_intrVec_3; // @[src/main/scala/nutcore/NutCore.scala 104:34]
  wire  frontend_io_out_1_bits_cf_intrVec_4; // @[src/main/scala/nutcore/NutCore.scala 104:34]
  wire  frontend_io_out_1_bits_cf_intrVec_5; // @[src/main/scala/nutcore/NutCore.scala 104:34]
  wire  frontend_io_out_1_bits_cf_intrVec_6; // @[src/main/scala/nutcore/NutCore.scala 104:34]
  wire  frontend_io_out_1_bits_cf_intrVec_7; // @[src/main/scala/nutcore/NutCore.scala 104:34]
  wire  frontend_io_out_1_bits_cf_intrVec_8; // @[src/main/scala/nutcore/NutCore.scala 104:34]
  wire  frontend_io_out_1_bits_cf_intrVec_9; // @[src/main/scala/nutcore/NutCore.scala 104:34]
  wire  frontend_io_out_1_bits_cf_intrVec_10; // @[src/main/scala/nutcore/NutCore.scala 104:34]
  wire  frontend_io_out_1_bits_cf_intrVec_11; // @[src/main/scala/nutcore/NutCore.scala 104:34]
  wire [3:0] frontend_io_flushVec; // @[src/main/scala/nutcore/NutCore.scala 104:34]
  wire [38:0] frontend_io_redirect_target; // @[src/main/scala/nutcore/NutCore.scala 104:34]
  wire  frontend_io_redirect_valid; // @[src/main/scala/nutcore/NutCore.scala 104:34]
  wire  frontend_io_ipf; // @[src/main/scala/nutcore/NutCore.scala 104:34]
  wire  frontend_REG_valid; // @[src/main/scala/nutcore/NutCore.scala 104:34]
  wire [38:0] frontend_REG_pc; // @[src/main/scala/nutcore/NutCore.scala 104:34]
  wire  frontend_REG_isMissPredict; // @[src/main/scala/nutcore/NutCore.scala 104:34]
  wire [38:0] frontend_REG_actualTarget; // @[src/main/scala/nutcore/NutCore.scala 104:34]
  wire  frontend_REG_actualTaken; // @[src/main/scala/nutcore/NutCore.scala 104:34]
  wire [6:0] frontend_REG_fuOpType; // @[src/main/scala/nutcore/NutCore.scala 104:34]
  wire [1:0] frontend_REG_btbType; // @[src/main/scala/nutcore/NutCore.scala 104:34]
  wire  frontend_REG_isRVC; // @[src/main/scala/nutcore/NutCore.scala 104:34]
  wire  frontend__WIRE_0; // @[src/main/scala/nutcore/NutCore.scala 104:34]
  wire  frontend_DISPLAY_ENABLE; // @[src/main/scala/nutcore/NutCore.scala 104:34]
  wire  frontend__WIRE_7; // @[src/main/scala/nutcore/NutCore.scala 104:34]
  wire  frontend__WIRE_11; // @[src/main/scala/nutcore/NutCore.scala 104:34]
  wire  frontend__WIRE_1_4; // @[src/main/scala/nutcore/NutCore.scala 104:34]
  wire [11:0] frontend__WIRE_14; // @[src/main/scala/nutcore/NutCore.scala 104:34]
  wire  frontend__WIRE_2_2; // @[src/main/scala/nutcore/NutCore.scala 104:34]
  wire  frontend_r_0; // @[src/main/scala/nutcore/NutCore.scala 104:34]
  wire  backend_clock; // @[src/main/scala/nutcore/NutCore.scala 147:25]
  wire  backend_reset; // @[src/main/scala/nutcore/NutCore.scala 147:25]
  wire  backend_io_in_0_ready; // @[src/main/scala/nutcore/NutCore.scala 147:25]
  wire  backend_io_in_0_valid; // @[src/main/scala/nutcore/NutCore.scala 147:25]
  wire [63:0] backend_io_in_0_bits_cf_instr; // @[src/main/scala/nutcore/NutCore.scala 147:25]
  wire [38:0] backend_io_in_0_bits_cf_pc; // @[src/main/scala/nutcore/NutCore.scala 147:25]
  wire [38:0] backend_io_in_0_bits_cf_pnpc; // @[src/main/scala/nutcore/NutCore.scala 147:25]
  wire  backend_io_in_0_bits_cf_exceptionVec_1; // @[src/main/scala/nutcore/NutCore.scala 147:25]
  wire  backend_io_in_0_bits_cf_exceptionVec_2; // @[src/main/scala/nutcore/NutCore.scala 147:25]
  wire  backend_io_in_0_bits_cf_exceptionVec_12; // @[src/main/scala/nutcore/NutCore.scala 147:25]
  wire  backend_io_in_0_bits_cf_intrVec_0; // @[src/main/scala/nutcore/NutCore.scala 147:25]
  wire  backend_io_in_0_bits_cf_intrVec_1; // @[src/main/scala/nutcore/NutCore.scala 147:25]
  wire  backend_io_in_0_bits_cf_intrVec_2; // @[src/main/scala/nutcore/NutCore.scala 147:25]
  wire  backend_io_in_0_bits_cf_intrVec_3; // @[src/main/scala/nutcore/NutCore.scala 147:25]
  wire  backend_io_in_0_bits_cf_intrVec_4; // @[src/main/scala/nutcore/NutCore.scala 147:25]
  wire  backend_io_in_0_bits_cf_intrVec_5; // @[src/main/scala/nutcore/NutCore.scala 147:25]
  wire  backend_io_in_0_bits_cf_intrVec_6; // @[src/main/scala/nutcore/NutCore.scala 147:25]
  wire  backend_io_in_0_bits_cf_intrVec_7; // @[src/main/scala/nutcore/NutCore.scala 147:25]
  wire  backend_io_in_0_bits_cf_intrVec_8; // @[src/main/scala/nutcore/NutCore.scala 147:25]
  wire  backend_io_in_0_bits_cf_intrVec_9; // @[src/main/scala/nutcore/NutCore.scala 147:25]
  wire  backend_io_in_0_bits_cf_intrVec_10; // @[src/main/scala/nutcore/NutCore.scala 147:25]
  wire  backend_io_in_0_bits_cf_intrVec_11; // @[src/main/scala/nutcore/NutCore.scala 147:25]
  wire [3:0] backend_io_in_0_bits_cf_brIdx; // @[src/main/scala/nutcore/NutCore.scala 147:25]
  wire  backend_io_in_0_bits_cf_crossPageIPFFix; // @[src/main/scala/nutcore/NutCore.scala 147:25]
  wire  backend_io_in_0_bits_ctrl_src1Type; // @[src/main/scala/nutcore/NutCore.scala 147:25]
  wire  backend_io_in_0_bits_ctrl_src2Type; // @[src/main/scala/nutcore/NutCore.scala 147:25]
  wire [2:0] backend_io_in_0_bits_ctrl_fuType; // @[src/main/scala/nutcore/NutCore.scala 147:25]
  wire [6:0] backend_io_in_0_bits_ctrl_fuOpType; // @[src/main/scala/nutcore/NutCore.scala 147:25]
  wire [4:0] backend_io_in_0_bits_ctrl_rfSrc1; // @[src/main/scala/nutcore/NutCore.scala 147:25]
  wire [4:0] backend_io_in_0_bits_ctrl_rfSrc2; // @[src/main/scala/nutcore/NutCore.scala 147:25]
  wire  backend_io_in_0_bits_ctrl_rfWen; // @[src/main/scala/nutcore/NutCore.scala 147:25]
  wire [4:0] backend_io_in_0_bits_ctrl_rfDest; // @[src/main/scala/nutcore/NutCore.scala 147:25]
  wire  backend_io_in_0_bits_ctrl_isNutCoreTrap; // @[src/main/scala/nutcore/NutCore.scala 147:25]
  wire [63:0] backend_io_in_0_bits_data_imm; // @[src/main/scala/nutcore/NutCore.scala 147:25]
  wire [1:0] backend_io_flush; // @[src/main/scala/nutcore/NutCore.scala 147:25]
  wire  backend_io_dmem_req_ready; // @[src/main/scala/nutcore/NutCore.scala 147:25]
  wire  backend_io_dmem_req_valid; // @[src/main/scala/nutcore/NutCore.scala 147:25]
  wire [38:0] backend_io_dmem_req_bits_addr; // @[src/main/scala/nutcore/NutCore.scala 147:25]
  wire [2:0] backend_io_dmem_req_bits_size; // @[src/main/scala/nutcore/NutCore.scala 147:25]
  wire [3:0] backend_io_dmem_req_bits_cmd; // @[src/main/scala/nutcore/NutCore.scala 147:25]
  wire [7:0] backend_io_dmem_req_bits_wmask; // @[src/main/scala/nutcore/NutCore.scala 147:25]
  wire [63:0] backend_io_dmem_req_bits_wdata; // @[src/main/scala/nutcore/NutCore.scala 147:25]
  wire  backend_io_dmem_resp_valid; // @[src/main/scala/nutcore/NutCore.scala 147:25]
  wire [63:0] backend_io_dmem_resp_bits_rdata; // @[src/main/scala/nutcore/NutCore.scala 147:25]
  wire [1:0] backend_io_memMMU_imem_priviledgeMode; // @[src/main/scala/nutcore/NutCore.scala 147:25]
  wire [1:0] backend_io_memMMU_dmem_priviledgeMode; // @[src/main/scala/nutcore/NutCore.scala 147:25]
  wire  backend_io_memMMU_dmem_status_sum; // @[src/main/scala/nutcore/NutCore.scala 147:25]
  wire  backend_io_memMMU_dmem_status_mxr; // @[src/main/scala/nutcore/NutCore.scala 147:25]
  wire  backend_io_memMMU_dmem_loadPF; // @[src/main/scala/nutcore/NutCore.scala 147:25]
  wire  backend_io_memMMU_dmem_storePF; // @[src/main/scala/nutcore/NutCore.scala 147:25]
  wire [38:0] backend_io_memMMU_dmem_addr; // @[src/main/scala/nutcore/NutCore.scala 147:25]
  wire [38:0] backend_io_redirect_target; // @[src/main/scala/nutcore/NutCore.scala 147:25]
  wire  backend_io_redirect_valid; // @[src/main/scala/nutcore/NutCore.scala 147:25]
  wire  backend_io_extra_meip_0; // @[src/main/scala/nutcore/NutCore.scala 147:25]
  wire  backend_REG_valid; // @[src/main/scala/nutcore/NutCore.scala 147:25]
  wire [38:0] backend_REG_pc; // @[src/main/scala/nutcore/NutCore.scala 147:25]
  wire  backend_REG_isMissPredict; // @[src/main/scala/nutcore/NutCore.scala 147:25]
  wire [38:0] backend_REG_actualTarget; // @[src/main/scala/nutcore/NutCore.scala 147:25]
  wire  backend_REG_actualTaken; // @[src/main/scala/nutcore/NutCore.scala 147:25]
  wire [6:0] backend_REG_fuOpType; // @[src/main/scala/nutcore/NutCore.scala 147:25]
  wire [1:0] backend_REG_btbType; // @[src/main/scala/nutcore/NutCore.scala 147:25]
  wire  backend_REG_isRVC; // @[src/main/scala/nutcore/NutCore.scala 147:25]
  wire  backend__WIRE_1; // @[src/main/scala/nutcore/NutCore.scala 147:25]
  wire [63:0] backend_satp; // @[src/main/scala/nutcore/NutCore.scala 147:25]
  wire  backend__WIRE_4; // @[src/main/scala/nutcore/NutCore.scala 147:25]
  wire  backend__WIRE_1_1; // @[src/main/scala/nutcore/NutCore.scala 147:25]
  wire  backend__WIRE_7; // @[src/main/scala/nutcore/NutCore.scala 147:25]
  wire  backend_io_extra_mtip; // @[src/main/scala/nutcore/NutCore.scala 147:25]
  wire  backend__WIRE_11; // @[src/main/scala/nutcore/NutCore.scala 147:25]
  wire  backend__WIRE_1_4; // @[src/main/scala/nutcore/NutCore.scala 147:25]
  wire [11:0] backend__WIRE_14; // @[src/main/scala/nutcore/NutCore.scala 147:25]
  wire  backend__WIRE_2_2; // @[src/main/scala/nutcore/NutCore.scala 147:25]
  wire  backend__WIRE_16; // @[src/main/scala/nutcore/NutCore.scala 147:25]
  wire  backend__WIRE_17; // @[src/main/scala/nutcore/NutCore.scala 147:25]
  wire  backend_r_0; // @[src/main/scala/nutcore/NutCore.scala 147:25]
  wire  backend_io_extra_msip; // @[src/main/scala/nutcore/NutCore.scala 147:25]
  wire  mmioXbar_clock; // @[src/main/scala/nutcore/NutCore.scala 151:26]
  wire  mmioXbar_reset; // @[src/main/scala/nutcore/NutCore.scala 151:26]
  wire  mmioXbar_io_in_0_req_ready; // @[src/main/scala/nutcore/NutCore.scala 151:26]
  wire  mmioXbar_io_in_0_req_valid; // @[src/main/scala/nutcore/NutCore.scala 151:26]
  wire [31:0] mmioXbar_io_in_0_req_bits_addr; // @[src/main/scala/nutcore/NutCore.scala 151:26]
  wire [3:0] mmioXbar_io_in_0_req_bits_cmd; // @[src/main/scala/nutcore/NutCore.scala 151:26]
  wire [7:0] mmioXbar_io_in_0_req_bits_wmask; // @[src/main/scala/nutcore/NutCore.scala 151:26]
  wire [63:0] mmioXbar_io_in_0_req_bits_wdata; // @[src/main/scala/nutcore/NutCore.scala 151:26]
  wire  mmioXbar_io_in_0_resp_valid; // @[src/main/scala/nutcore/NutCore.scala 151:26]
  wire [3:0] mmioXbar_io_in_0_resp_bits_cmd; // @[src/main/scala/nutcore/NutCore.scala 151:26]
  wire [63:0] mmioXbar_io_in_0_resp_bits_rdata; // @[src/main/scala/nutcore/NutCore.scala 151:26]
  wire  mmioXbar_io_in_1_req_ready; // @[src/main/scala/nutcore/NutCore.scala 151:26]
  wire  mmioXbar_io_in_1_req_valid; // @[src/main/scala/nutcore/NutCore.scala 151:26]
  wire [31:0] mmioXbar_io_in_1_req_bits_addr; // @[src/main/scala/nutcore/NutCore.scala 151:26]
  wire [2:0] mmioXbar_io_in_1_req_bits_size; // @[src/main/scala/nutcore/NutCore.scala 151:26]
  wire [3:0] mmioXbar_io_in_1_req_bits_cmd; // @[src/main/scala/nutcore/NutCore.scala 151:26]
  wire [7:0] mmioXbar_io_in_1_req_bits_wmask; // @[src/main/scala/nutcore/NutCore.scala 151:26]
  wire [63:0] mmioXbar_io_in_1_req_bits_wdata; // @[src/main/scala/nutcore/NutCore.scala 151:26]
  wire  mmioXbar_io_in_1_resp_valid; // @[src/main/scala/nutcore/NutCore.scala 151:26]
  wire [3:0] mmioXbar_io_in_1_resp_bits_cmd; // @[src/main/scala/nutcore/NutCore.scala 151:26]
  wire [63:0] mmioXbar_io_in_1_resp_bits_rdata; // @[src/main/scala/nutcore/NutCore.scala 151:26]
  wire  mmioXbar_io_out_req_ready; // @[src/main/scala/nutcore/NutCore.scala 151:26]
  wire  mmioXbar_io_out_req_valid; // @[src/main/scala/nutcore/NutCore.scala 151:26]
  wire [31:0] mmioXbar_io_out_req_bits_addr; // @[src/main/scala/nutcore/NutCore.scala 151:26]
  wire [2:0] mmioXbar_io_out_req_bits_size; // @[src/main/scala/nutcore/NutCore.scala 151:26]
  wire [3:0] mmioXbar_io_out_req_bits_cmd; // @[src/main/scala/nutcore/NutCore.scala 151:26]
  wire [7:0] mmioXbar_io_out_req_bits_wmask; // @[src/main/scala/nutcore/NutCore.scala 151:26]
  wire [63:0] mmioXbar_io_out_req_bits_wdata; // @[src/main/scala/nutcore/NutCore.scala 151:26]
  wire  mmioXbar_io_out_resp_ready; // @[src/main/scala/nutcore/NutCore.scala 151:26]
  wire  mmioXbar_io_out_resp_valid; // @[src/main/scala/nutcore/NutCore.scala 151:26]
  wire [3:0] mmioXbar_io_out_resp_bits_cmd; // @[src/main/scala/nutcore/NutCore.scala 151:26]
  wire [63:0] mmioXbar_io_out_resp_bits_rdata; // @[src/main/scala/nutcore/NutCore.scala 151:26]
  wire  dmemXbar_clock; // @[src/main/scala/nutcore/NutCore.scala 152:26]
  wire  dmemXbar_reset; // @[src/main/scala/nutcore/NutCore.scala 152:26]
  wire  dmemXbar_io_in_0_req_ready; // @[src/main/scala/nutcore/NutCore.scala 152:26]
  wire  dmemXbar_io_in_0_req_valid; // @[src/main/scala/nutcore/NutCore.scala 152:26]
  wire [31:0] dmemXbar_io_in_0_req_bits_addr; // @[src/main/scala/nutcore/NutCore.scala 152:26]
  wire [2:0] dmemXbar_io_in_0_req_bits_size; // @[src/main/scala/nutcore/NutCore.scala 152:26]
  wire [3:0] dmemXbar_io_in_0_req_bits_cmd; // @[src/main/scala/nutcore/NutCore.scala 152:26]
  wire [7:0] dmemXbar_io_in_0_req_bits_wmask; // @[src/main/scala/nutcore/NutCore.scala 152:26]
  wire [63:0] dmemXbar_io_in_0_req_bits_wdata; // @[src/main/scala/nutcore/NutCore.scala 152:26]
  wire  dmemXbar_io_in_0_resp_valid; // @[src/main/scala/nutcore/NutCore.scala 152:26]
  wire [3:0] dmemXbar_io_in_0_resp_bits_cmd; // @[src/main/scala/nutcore/NutCore.scala 152:26]
  wire [63:0] dmemXbar_io_in_0_resp_bits_rdata; // @[src/main/scala/nutcore/NutCore.scala 152:26]
  wire  dmemXbar_io_in_1_req_ready; // @[src/main/scala/nutcore/NutCore.scala 152:26]
  wire  dmemXbar_io_in_1_req_valid; // @[src/main/scala/nutcore/NutCore.scala 152:26]
  wire [31:0] dmemXbar_io_in_1_req_bits_addr; // @[src/main/scala/nutcore/NutCore.scala 152:26]
  wire [3:0] dmemXbar_io_in_1_req_bits_cmd; // @[src/main/scala/nutcore/NutCore.scala 152:26]
  wire [63:0] dmemXbar_io_in_1_req_bits_wdata; // @[src/main/scala/nutcore/NutCore.scala 152:26]
  wire  dmemXbar_io_in_1_resp_valid; // @[src/main/scala/nutcore/NutCore.scala 152:26]
  wire [3:0] dmemXbar_io_in_1_resp_bits_cmd; // @[src/main/scala/nutcore/NutCore.scala 152:26]
  wire [63:0] dmemXbar_io_in_1_resp_bits_rdata; // @[src/main/scala/nutcore/NutCore.scala 152:26]
  wire  dmemXbar_io_in_2_req_ready; // @[src/main/scala/nutcore/NutCore.scala 152:26]
  wire  dmemXbar_io_in_2_req_valid; // @[src/main/scala/nutcore/NutCore.scala 152:26]
  wire [31:0] dmemXbar_io_in_2_req_bits_addr; // @[src/main/scala/nutcore/NutCore.scala 152:26]
  wire [3:0] dmemXbar_io_in_2_req_bits_cmd; // @[src/main/scala/nutcore/NutCore.scala 152:26]
  wire [63:0] dmemXbar_io_in_2_req_bits_wdata; // @[src/main/scala/nutcore/NutCore.scala 152:26]
  wire  dmemXbar_io_in_2_resp_valid; // @[src/main/scala/nutcore/NutCore.scala 152:26]
  wire [3:0] dmemXbar_io_in_2_resp_bits_cmd; // @[src/main/scala/nutcore/NutCore.scala 152:26]
  wire [63:0] dmemXbar_io_in_2_resp_bits_rdata; // @[src/main/scala/nutcore/NutCore.scala 152:26]
  wire  dmemXbar_io_in_3_req_ready; // @[src/main/scala/nutcore/NutCore.scala 152:26]
  wire  dmemXbar_io_in_3_req_valid; // @[src/main/scala/nutcore/NutCore.scala 152:26]
  wire [31:0] dmemXbar_io_in_3_req_bits_addr; // @[src/main/scala/nutcore/NutCore.scala 152:26]
  wire [2:0] dmemXbar_io_in_3_req_bits_size; // @[src/main/scala/nutcore/NutCore.scala 152:26]
  wire [3:0] dmemXbar_io_in_3_req_bits_cmd; // @[src/main/scala/nutcore/NutCore.scala 152:26]
  wire [7:0] dmemXbar_io_in_3_req_bits_wmask; // @[src/main/scala/nutcore/NutCore.scala 152:26]
  wire [63:0] dmemXbar_io_in_3_req_bits_wdata; // @[src/main/scala/nutcore/NutCore.scala 152:26]
  wire  dmemXbar_io_in_3_resp_ready; // @[src/main/scala/nutcore/NutCore.scala 152:26]
  wire  dmemXbar_io_in_3_resp_valid; // @[src/main/scala/nutcore/NutCore.scala 152:26]
  wire [3:0] dmemXbar_io_in_3_resp_bits_cmd; // @[src/main/scala/nutcore/NutCore.scala 152:26]
  wire [63:0] dmemXbar_io_in_3_resp_bits_rdata; // @[src/main/scala/nutcore/NutCore.scala 152:26]
  wire  dmemXbar_io_out_req_ready; // @[src/main/scala/nutcore/NutCore.scala 152:26]
  wire  dmemXbar_io_out_req_valid; // @[src/main/scala/nutcore/NutCore.scala 152:26]
  wire [31:0] dmemXbar_io_out_req_bits_addr; // @[src/main/scala/nutcore/NutCore.scala 152:26]
  wire [2:0] dmemXbar_io_out_req_bits_size; // @[src/main/scala/nutcore/NutCore.scala 152:26]
  wire [3:0] dmemXbar_io_out_req_bits_cmd; // @[src/main/scala/nutcore/NutCore.scala 152:26]
  wire [7:0] dmemXbar_io_out_req_bits_wmask; // @[src/main/scala/nutcore/NutCore.scala 152:26]
  wire [63:0] dmemXbar_io_out_req_bits_wdata; // @[src/main/scala/nutcore/NutCore.scala 152:26]
  wire  dmemXbar_io_out_resp_ready; // @[src/main/scala/nutcore/NutCore.scala 152:26]
  wire  dmemXbar_io_out_resp_valid; // @[src/main/scala/nutcore/NutCore.scala 152:26]
  wire [3:0] dmemXbar_io_out_resp_bits_cmd; // @[src/main/scala/nutcore/NutCore.scala 152:26]
  wire [63:0] dmemXbar_io_out_resp_bits_rdata; // @[src/main/scala/nutcore/NutCore.scala 152:26]
  wire  itlb_clock; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 426:13]
  wire  itlb_reset; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 426:13]
  wire  itlb_io_in_req_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 426:13]
  wire  itlb_io_in_req_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 426:13]
  wire [38:0] itlb_io_in_req_bits_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 426:13]
  wire [86:0] itlb_io_in_req_bits_user; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 426:13]
  wire  itlb_io_in_resp_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 426:13]
  wire  itlb_io_in_resp_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 426:13]
  wire [3:0] itlb_io_in_resp_bits_cmd; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 426:13]
  wire [63:0] itlb_io_in_resp_bits_rdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 426:13]
  wire [86:0] itlb_io_in_resp_bits_user; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 426:13]
  wire  itlb_io_out_req_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 426:13]
  wire  itlb_io_out_req_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 426:13]
  wire [31:0] itlb_io_out_req_bits_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 426:13]
  wire [3:0] itlb_io_out_req_bits_cmd; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 426:13]
  wire [63:0] itlb_io_out_req_bits_wdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 426:13]
  wire [86:0] itlb_io_out_req_bits_user; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 426:13]
  wire  itlb_io_out_resp_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 426:13]
  wire  itlb_io_out_resp_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 426:13]
  wire [63:0] itlb_io_out_resp_bits_rdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 426:13]
  wire [86:0] itlb_io_out_resp_bits_user; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 426:13]
  wire  itlb_io_mem_req_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 426:13]
  wire  itlb_io_mem_req_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 426:13]
  wire [31:0] itlb_io_mem_req_bits_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 426:13]
  wire [3:0] itlb_io_mem_req_bits_cmd; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 426:13]
  wire [63:0] itlb_io_mem_req_bits_wdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 426:13]
  wire  itlb_io_mem_resp_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 426:13]
  wire [3:0] itlb_io_mem_resp_bits_cmd; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 426:13]
  wire [63:0] itlb_io_mem_resp_bits_rdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 426:13]
  wire  itlb_io_flush; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 426:13]
  wire [1:0] itlb_io_csrMMU_priviledgeMode; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 426:13]
  wire  itlb_io_csrMMU_loadPF; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 426:13]
  wire  itlb_io_csrMMU_storePF; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 426:13]
  wire  itlb_io_cacheEmpty; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 426:13]
  wire  itlb_io_ipf; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 426:13]
  wire [63:0] itlb_CSRSATP; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 426:13]
  wire  itlb_DISPLAY_ENABLE; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 426:13]
  wire  itlb_MOUFlushTLB; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 426:13]
  wire  io_imem_cache_clock; // @[src/main/scala/nutcore/mem/Cache.scala 668:35]
  wire  io_imem_cache_reset; // @[src/main/scala/nutcore/mem/Cache.scala 668:35]
  wire  io_imem_cache_io_in_req_ready; // @[src/main/scala/nutcore/mem/Cache.scala 668:35]
  wire  io_imem_cache_io_in_req_valid; // @[src/main/scala/nutcore/mem/Cache.scala 668:35]
  wire [31:0] io_imem_cache_io_in_req_bits_addr; // @[src/main/scala/nutcore/mem/Cache.scala 668:35]
  wire [86:0] io_imem_cache_io_in_req_bits_user; // @[src/main/scala/nutcore/mem/Cache.scala 668:35]
  wire  io_imem_cache_io_in_resp_ready; // @[src/main/scala/nutcore/mem/Cache.scala 668:35]
  wire  io_imem_cache_io_in_resp_valid; // @[src/main/scala/nutcore/mem/Cache.scala 668:35]
  wire [63:0] io_imem_cache_io_in_resp_bits_rdata; // @[src/main/scala/nutcore/mem/Cache.scala 668:35]
  wire [86:0] io_imem_cache_io_in_resp_bits_user; // @[src/main/scala/nutcore/mem/Cache.scala 668:35]
  wire [1:0] io_imem_cache_io_flush; // @[src/main/scala/nutcore/mem/Cache.scala 668:35]
  wire  io_imem_cache_io_out_mem_req_ready; // @[src/main/scala/nutcore/mem/Cache.scala 668:35]
  wire  io_imem_cache_io_out_mem_req_valid; // @[src/main/scala/nutcore/mem/Cache.scala 668:35]
  wire [31:0] io_imem_cache_io_out_mem_req_bits_addr; // @[src/main/scala/nutcore/mem/Cache.scala 668:35]
  wire [3:0] io_imem_cache_io_out_mem_req_bits_cmd; // @[src/main/scala/nutcore/mem/Cache.scala 668:35]
  wire [63:0] io_imem_cache_io_out_mem_req_bits_wdata; // @[src/main/scala/nutcore/mem/Cache.scala 668:35]
  wire  io_imem_cache_io_out_mem_resp_valid; // @[src/main/scala/nutcore/mem/Cache.scala 668:35]
  wire [3:0] io_imem_cache_io_out_mem_resp_bits_cmd; // @[src/main/scala/nutcore/mem/Cache.scala 668:35]
  wire [63:0] io_imem_cache_io_out_mem_resp_bits_rdata; // @[src/main/scala/nutcore/mem/Cache.scala 668:35]
  wire  io_imem_cache_io_mmio_req_ready; // @[src/main/scala/nutcore/mem/Cache.scala 668:35]
  wire  io_imem_cache_io_mmio_req_valid; // @[src/main/scala/nutcore/mem/Cache.scala 668:35]
  wire [31:0] io_imem_cache_io_mmio_req_bits_addr; // @[src/main/scala/nutcore/mem/Cache.scala 668:35]
  wire  io_imem_cache_io_mmio_resp_valid; // @[src/main/scala/nutcore/mem/Cache.scala 668:35]
  wire [63:0] io_imem_cache_io_mmio_resp_bits_rdata; // @[src/main/scala/nutcore/mem/Cache.scala 668:35]
  wire  io_imem_cache_io_empty; // @[src/main/scala/nutcore/mem/Cache.scala 668:35]
  wire  io_imem_cache_DISPLAY_ENABLE; // @[src/main/scala/nutcore/mem/Cache.scala 668:35]
  wire  io_imem_cache_MOUFlushICache; // @[src/main/scala/nutcore/mem/Cache.scala 668:35]
  wire  dtlb_clock; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 426:13]
  wire  dtlb_reset; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 426:13]
  wire  dtlb_io_in_req_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 426:13]
  wire  dtlb_io_in_req_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 426:13]
  wire [38:0] dtlb_io_in_req_bits_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 426:13]
  wire [2:0] dtlb_io_in_req_bits_size; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 426:13]
  wire [3:0] dtlb_io_in_req_bits_cmd; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 426:13]
  wire [7:0] dtlb_io_in_req_bits_wmask; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 426:13]
  wire [63:0] dtlb_io_in_req_bits_wdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 426:13]
  wire  dtlb_io_in_resp_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 426:13]
  wire [3:0] dtlb_io_in_resp_bits_cmd; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 426:13]
  wire [63:0] dtlb_io_in_resp_bits_rdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 426:13]
  wire  dtlb_io_out_req_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 426:13]
  wire  dtlb_io_out_req_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 426:13]
  wire [31:0] dtlb_io_out_req_bits_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 426:13]
  wire [2:0] dtlb_io_out_req_bits_size; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 426:13]
  wire [3:0] dtlb_io_out_req_bits_cmd; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 426:13]
  wire [7:0] dtlb_io_out_req_bits_wmask; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 426:13]
  wire [63:0] dtlb_io_out_req_bits_wdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 426:13]
  wire  dtlb_io_out_resp_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 426:13]
  wire  dtlb_io_out_resp_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 426:13]
  wire [3:0] dtlb_io_out_resp_bits_cmd; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 426:13]
  wire [63:0] dtlb_io_out_resp_bits_rdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 426:13]
  wire  dtlb_io_mem_req_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 426:13]
  wire  dtlb_io_mem_req_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 426:13]
  wire [31:0] dtlb_io_mem_req_bits_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 426:13]
  wire [3:0] dtlb_io_mem_req_bits_cmd; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 426:13]
  wire [63:0] dtlb_io_mem_req_bits_wdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 426:13]
  wire  dtlb_io_mem_resp_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 426:13]
  wire [3:0] dtlb_io_mem_resp_bits_cmd; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 426:13]
  wire [63:0] dtlb_io_mem_resp_bits_rdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 426:13]
  wire [1:0] dtlb_io_csrMMU_priviledgeMode; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 426:13]
  wire  dtlb_io_csrMMU_status_sum; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 426:13]
  wire  dtlb_io_csrMMU_status_mxr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 426:13]
  wire  dtlb_io_csrMMU_loadPF; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 426:13]
  wire  dtlb_io_csrMMU_storePF; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 426:13]
  wire [38:0] dtlb_io_csrMMU_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 426:13]
  wire  dtlb_io_cacheEmpty; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 426:13]
  wire  dtlb_io_ipf; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 426:13]
  wire  dtlb__WIRE_4; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 426:13]
  wire [63:0] dtlb_CSRSATP; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 426:13]
  wire  dtlb_DISPLAY_ENABLE; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 426:13]
  wire  dtlb__WIRE_1_1; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 426:13]
  wire  dtlb_MOUFlushTLB; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 426:13]
  wire  dtlb__WIRE_2_3; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 426:13]
  wire  dtlb__WIRE_16; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 426:13]
  wire  io_dmem_cache_clock; // @[src/main/scala/nutcore/mem/Cache.scala 668:35]
  wire  io_dmem_cache_reset; // @[src/main/scala/nutcore/mem/Cache.scala 668:35]
  wire  io_dmem_cache_io_in_req_ready; // @[src/main/scala/nutcore/mem/Cache.scala 668:35]
  wire  io_dmem_cache_io_in_req_valid; // @[src/main/scala/nutcore/mem/Cache.scala 668:35]
  wire [31:0] io_dmem_cache_io_in_req_bits_addr; // @[src/main/scala/nutcore/mem/Cache.scala 668:35]
  wire [2:0] io_dmem_cache_io_in_req_bits_size; // @[src/main/scala/nutcore/mem/Cache.scala 668:35]
  wire [3:0] io_dmem_cache_io_in_req_bits_cmd; // @[src/main/scala/nutcore/mem/Cache.scala 668:35]
  wire [7:0] io_dmem_cache_io_in_req_bits_wmask; // @[src/main/scala/nutcore/mem/Cache.scala 668:35]
  wire [63:0] io_dmem_cache_io_in_req_bits_wdata; // @[src/main/scala/nutcore/mem/Cache.scala 668:35]
  wire  io_dmem_cache_io_in_resp_ready; // @[src/main/scala/nutcore/mem/Cache.scala 668:35]
  wire  io_dmem_cache_io_in_resp_valid; // @[src/main/scala/nutcore/mem/Cache.scala 668:35]
  wire [3:0] io_dmem_cache_io_in_resp_bits_cmd; // @[src/main/scala/nutcore/mem/Cache.scala 668:35]
  wire [63:0] io_dmem_cache_io_in_resp_bits_rdata; // @[src/main/scala/nutcore/mem/Cache.scala 668:35]
  wire  io_dmem_cache_io_out_mem_req_ready; // @[src/main/scala/nutcore/mem/Cache.scala 668:35]
  wire  io_dmem_cache_io_out_mem_req_valid; // @[src/main/scala/nutcore/mem/Cache.scala 668:35]
  wire [31:0] io_dmem_cache_io_out_mem_req_bits_addr; // @[src/main/scala/nutcore/mem/Cache.scala 668:35]
  wire [3:0] io_dmem_cache_io_out_mem_req_bits_cmd; // @[src/main/scala/nutcore/mem/Cache.scala 668:35]
  wire [63:0] io_dmem_cache_io_out_mem_req_bits_wdata; // @[src/main/scala/nutcore/mem/Cache.scala 668:35]
  wire  io_dmem_cache_io_out_mem_resp_valid; // @[src/main/scala/nutcore/mem/Cache.scala 668:35]
  wire [3:0] io_dmem_cache_io_out_mem_resp_bits_cmd; // @[src/main/scala/nutcore/mem/Cache.scala 668:35]
  wire [63:0] io_dmem_cache_io_out_mem_resp_bits_rdata; // @[src/main/scala/nutcore/mem/Cache.scala 668:35]
  wire  io_dmem_cache_io_out_coh_req_ready; // @[src/main/scala/nutcore/mem/Cache.scala 668:35]
  wire  io_dmem_cache_io_out_coh_req_valid; // @[src/main/scala/nutcore/mem/Cache.scala 668:35]
  wire [31:0] io_dmem_cache_io_out_coh_req_bits_addr; // @[src/main/scala/nutcore/mem/Cache.scala 668:35]
  wire [63:0] io_dmem_cache_io_out_coh_req_bits_wdata; // @[src/main/scala/nutcore/mem/Cache.scala 668:35]
  wire  io_dmem_cache_io_out_coh_resp_valid; // @[src/main/scala/nutcore/mem/Cache.scala 668:35]
  wire [3:0] io_dmem_cache_io_out_coh_resp_bits_cmd; // @[src/main/scala/nutcore/mem/Cache.scala 668:35]
  wire [63:0] io_dmem_cache_io_out_coh_resp_bits_rdata; // @[src/main/scala/nutcore/mem/Cache.scala 668:35]
  wire  io_dmem_cache_io_mmio_req_ready; // @[src/main/scala/nutcore/mem/Cache.scala 668:35]
  wire  io_dmem_cache_io_mmio_req_valid; // @[src/main/scala/nutcore/mem/Cache.scala 668:35]
  wire [31:0] io_dmem_cache_io_mmio_req_bits_addr; // @[src/main/scala/nutcore/mem/Cache.scala 668:35]
  wire [2:0] io_dmem_cache_io_mmio_req_bits_size; // @[src/main/scala/nutcore/mem/Cache.scala 668:35]
  wire [3:0] io_dmem_cache_io_mmio_req_bits_cmd; // @[src/main/scala/nutcore/mem/Cache.scala 668:35]
  wire [7:0] io_dmem_cache_io_mmio_req_bits_wmask; // @[src/main/scala/nutcore/mem/Cache.scala 668:35]
  wire [63:0] io_dmem_cache_io_mmio_req_bits_wdata; // @[src/main/scala/nutcore/mem/Cache.scala 668:35]
  wire  io_dmem_cache_io_mmio_resp_valid; // @[src/main/scala/nutcore/mem/Cache.scala 668:35]
  wire [63:0] io_dmem_cache_io_mmio_resp_bits_rdata; // @[src/main/scala/nutcore/mem/Cache.scala 668:35]
  wire  io_dmem_cache_io_empty; // @[src/main/scala/nutcore/mem/Cache.scala 668:35]
  wire  io_dmem_cache_DISPLAY_ENABLE; // @[src/main/scala/nutcore/mem/Cache.scala 668:35]
  wire  io_dmem_cache__WIRE_17; // @[src/main/scala/nutcore/mem/Cache.scala 668:35]
  reg [63:0] dataBuffer_0_cf_instr; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [38:0] dataBuffer_0_cf_pc; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [38:0] dataBuffer_0_cf_pnpc; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_0_cf_exceptionVec_1; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_0_cf_exceptionVec_2; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_0_cf_exceptionVec_12; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_0_cf_intrVec_0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_0_cf_intrVec_1; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_0_cf_intrVec_2; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_0_cf_intrVec_3; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_0_cf_intrVec_4; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_0_cf_intrVec_5; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_0_cf_intrVec_6; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_0_cf_intrVec_7; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_0_cf_intrVec_8; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_0_cf_intrVec_9; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_0_cf_intrVec_10; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_0_cf_intrVec_11; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [3:0] dataBuffer_0_cf_brIdx; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_0_cf_crossPageIPFFix; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_0_ctrl_src1Type; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_0_ctrl_src2Type; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [2:0] dataBuffer_0_ctrl_fuType; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [6:0] dataBuffer_0_ctrl_fuOpType; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [4:0] dataBuffer_0_ctrl_rfSrc1; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [4:0] dataBuffer_0_ctrl_rfSrc2; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_0_ctrl_rfWen; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [4:0] dataBuffer_0_ctrl_rfDest; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_0_ctrl_isNutCoreTrap; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [63:0] dataBuffer_0_data_imm; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [63:0] dataBuffer_1_cf_instr; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [38:0] dataBuffer_1_cf_pc; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [38:0] dataBuffer_1_cf_pnpc; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_1_cf_exceptionVec_1; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_1_cf_exceptionVec_2; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_1_cf_exceptionVec_12; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_1_cf_intrVec_0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_1_cf_intrVec_1; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_1_cf_intrVec_2; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_1_cf_intrVec_3; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_1_cf_intrVec_4; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_1_cf_intrVec_5; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_1_cf_intrVec_6; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_1_cf_intrVec_7; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_1_cf_intrVec_8; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_1_cf_intrVec_9; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_1_cf_intrVec_10; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_1_cf_intrVec_11; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [3:0] dataBuffer_1_cf_brIdx; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_1_cf_crossPageIPFFix; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_1_ctrl_src1Type; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_1_ctrl_src2Type; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [2:0] dataBuffer_1_ctrl_fuType; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [6:0] dataBuffer_1_ctrl_fuOpType; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [4:0] dataBuffer_1_ctrl_rfSrc1; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [4:0] dataBuffer_1_ctrl_rfSrc2; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_1_ctrl_rfWen; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [4:0] dataBuffer_1_ctrl_rfDest; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_1_ctrl_isNutCoreTrap; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [63:0] dataBuffer_1_data_imm; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [63:0] dataBuffer_2_cf_instr; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [38:0] dataBuffer_2_cf_pc; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [38:0] dataBuffer_2_cf_pnpc; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_2_cf_exceptionVec_1; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_2_cf_exceptionVec_2; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_2_cf_exceptionVec_12; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_2_cf_intrVec_0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_2_cf_intrVec_1; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_2_cf_intrVec_2; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_2_cf_intrVec_3; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_2_cf_intrVec_4; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_2_cf_intrVec_5; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_2_cf_intrVec_6; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_2_cf_intrVec_7; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_2_cf_intrVec_8; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_2_cf_intrVec_9; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_2_cf_intrVec_10; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_2_cf_intrVec_11; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [3:0] dataBuffer_2_cf_brIdx; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_2_cf_crossPageIPFFix; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_2_ctrl_src1Type; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_2_ctrl_src2Type; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [2:0] dataBuffer_2_ctrl_fuType; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [6:0] dataBuffer_2_ctrl_fuOpType; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [4:0] dataBuffer_2_ctrl_rfSrc1; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [4:0] dataBuffer_2_ctrl_rfSrc2; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_2_ctrl_rfWen; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [4:0] dataBuffer_2_ctrl_rfDest; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_2_ctrl_isNutCoreTrap; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [63:0] dataBuffer_2_data_imm; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [63:0] dataBuffer_3_cf_instr; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [38:0] dataBuffer_3_cf_pc; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [38:0] dataBuffer_3_cf_pnpc; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_3_cf_exceptionVec_1; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_3_cf_exceptionVec_2; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_3_cf_exceptionVec_12; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_3_cf_intrVec_0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_3_cf_intrVec_1; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_3_cf_intrVec_2; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_3_cf_intrVec_3; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_3_cf_intrVec_4; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_3_cf_intrVec_5; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_3_cf_intrVec_6; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_3_cf_intrVec_7; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_3_cf_intrVec_8; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_3_cf_intrVec_9; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_3_cf_intrVec_10; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_3_cf_intrVec_11; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [3:0] dataBuffer_3_cf_brIdx; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_3_cf_crossPageIPFFix; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_3_ctrl_src1Type; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_3_ctrl_src2Type; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [2:0] dataBuffer_3_ctrl_fuType; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [6:0] dataBuffer_3_ctrl_fuOpType; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [4:0] dataBuffer_3_ctrl_rfSrc1; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [4:0] dataBuffer_3_ctrl_rfSrc2; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_3_ctrl_rfWen; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [4:0] dataBuffer_3_ctrl_rfDest; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_3_ctrl_isNutCoreTrap; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [63:0] dataBuffer_3_data_imm; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [1:0] ringBufferHead; // @[src/main/scala/utils/PipelineVector.scala 30:33]
  reg [1:0] ringBufferTail; // @[src/main/scala/utils/PipelineVector.scala 31:33]
  wire [1:0] _ringBufferAllowin_T_1 = ringBufferHead + 2'h1; // @[src/main/scala/utils/PipelineVector.scala 33:63]
  wire [1:0] _ringBufferAllowin_T_4 = ringBufferHead + 2'h2; // @[src/main/scala/utils/PipelineVector.scala 33:63]
  wire  ringBufferAllowin = _ringBufferAllowin_T_1 != ringBufferTail & _ringBufferAllowin_T_4 != ringBufferTail; // @[src/main/scala/utils/PipelineVector.scala 33:124]
  wire  needEnqueue_0 = frontend_io_out_0_valid; // @[src/main/scala/utils/PipelineVector.scala 36:27 37:20]
  wire [1:0] enqueueSize = {{1'd0}, needEnqueue_0}; // @[src/main/scala/utils/PipelineVector.scala 40:44]
  wire  enqueueFire_0 = enqueueSize >= 2'h1; // @[src/main/scala/utils/PipelineVector.scala 41:53]
  wire  enqueueFire_1 = enqueueSize >= 2'h2; // @[src/main/scala/utils/PipelineVector.scala 41:53]
  wire  wen = frontend_io_out_0_ready & frontend_io_out_0_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  wire [2:0] _T_1 = {{1'd0}, ringBufferHead}; // @[src/main/scala/utils/PipelineVector.scala 45:45]
  wire [63:0] _dataBuffer_T_cf_instr = needEnqueue_0 ? frontend_io_out_0_bits_cf_instr : 64'h0; // @[src/main/scala/utils/PipelineVector.scala 45:69]
  wire [38:0] _dataBuffer_T_cf_pc = needEnqueue_0 ? frontend_io_out_0_bits_cf_pc : 39'h0; // @[src/main/scala/utils/PipelineVector.scala 45:69]
  wire [38:0] _dataBuffer_T_cf_pnpc = needEnqueue_0 ? frontend_io_out_0_bits_cf_pnpc : 39'h0; // @[src/main/scala/utils/PipelineVector.scala 45:69]
  wire  _dataBuffer_T_cf_intrVec_0 = needEnqueue_0 ? frontend_io_out_0_bits_cf_intrVec_0 :
    frontend_io_out_1_bits_cf_intrVec_0; // @[src/main/scala/utils/PipelineVector.scala 45:69]
  wire  _dataBuffer_T_cf_intrVec_1 = needEnqueue_0 ? frontend_io_out_0_bits_cf_intrVec_1 :
    frontend_io_out_1_bits_cf_intrVec_1; // @[src/main/scala/utils/PipelineVector.scala 45:69]
  wire  _dataBuffer_T_cf_intrVec_2 = needEnqueue_0 ? frontend_io_out_0_bits_cf_intrVec_2 :
    frontend_io_out_1_bits_cf_intrVec_2; // @[src/main/scala/utils/PipelineVector.scala 45:69]
  wire  _dataBuffer_T_cf_intrVec_3 = needEnqueue_0 ? frontend_io_out_0_bits_cf_intrVec_3 :
    frontend_io_out_1_bits_cf_intrVec_3; // @[src/main/scala/utils/PipelineVector.scala 45:69]
  wire  _dataBuffer_T_cf_intrVec_4 = needEnqueue_0 ? frontend_io_out_0_bits_cf_intrVec_4 :
    frontend_io_out_1_bits_cf_intrVec_4; // @[src/main/scala/utils/PipelineVector.scala 45:69]
  wire  _dataBuffer_T_cf_intrVec_5 = needEnqueue_0 ? frontend_io_out_0_bits_cf_intrVec_5 :
    frontend_io_out_1_bits_cf_intrVec_5; // @[src/main/scala/utils/PipelineVector.scala 45:69]
  wire  _dataBuffer_T_cf_intrVec_6 = needEnqueue_0 ? frontend_io_out_0_bits_cf_intrVec_6 :
    frontend_io_out_1_bits_cf_intrVec_6; // @[src/main/scala/utils/PipelineVector.scala 45:69]
  wire  _dataBuffer_T_cf_intrVec_7 = needEnqueue_0 ? frontend_io_out_0_bits_cf_intrVec_7 :
    frontend_io_out_1_bits_cf_intrVec_7; // @[src/main/scala/utils/PipelineVector.scala 45:69]
  wire  _dataBuffer_T_cf_intrVec_8 = needEnqueue_0 ? frontend_io_out_0_bits_cf_intrVec_8 :
    frontend_io_out_1_bits_cf_intrVec_8; // @[src/main/scala/utils/PipelineVector.scala 45:69]
  wire  _dataBuffer_T_cf_intrVec_9 = needEnqueue_0 ? frontend_io_out_0_bits_cf_intrVec_9 :
    frontend_io_out_1_bits_cf_intrVec_9; // @[src/main/scala/utils/PipelineVector.scala 45:69]
  wire  _dataBuffer_T_cf_intrVec_10 = needEnqueue_0 ? frontend_io_out_0_bits_cf_intrVec_10 :
    frontend_io_out_1_bits_cf_intrVec_10; // @[src/main/scala/utils/PipelineVector.scala 45:69]
  wire  _dataBuffer_T_cf_intrVec_11 = needEnqueue_0 ? frontend_io_out_0_bits_cf_intrVec_11 :
    frontend_io_out_1_bits_cf_intrVec_11; // @[src/main/scala/utils/PipelineVector.scala 45:69]
  wire [3:0] _dataBuffer_T_cf_brIdx = needEnqueue_0 ? frontend_io_out_0_bits_cf_brIdx : 4'h0; // @[src/main/scala/utils/PipelineVector.scala 45:69]
  wire  _dataBuffer_T_ctrl_src1Type = needEnqueue_0 ? frontend_io_out_0_bits_ctrl_src1Type : 1'h1; // @[src/main/scala/utils/PipelineVector.scala 45:69]
  wire  _dataBuffer_T_ctrl_src2Type = needEnqueue_0 ? frontend_io_out_0_bits_ctrl_src2Type : 1'h1; // @[src/main/scala/utils/PipelineVector.scala 45:69]
  wire [2:0] _dataBuffer_T_ctrl_fuType = needEnqueue_0 ? frontend_io_out_0_bits_ctrl_fuType : 3'h3; // @[src/main/scala/utils/PipelineVector.scala 45:69]
  wire [6:0] _dataBuffer_T_ctrl_fuOpType = needEnqueue_0 ? frontend_io_out_0_bits_ctrl_fuOpType : 7'h0; // @[src/main/scala/utils/PipelineVector.scala 45:69]
  wire [4:0] _dataBuffer_T_ctrl_rfSrc1 = needEnqueue_0 ? frontend_io_out_0_bits_ctrl_rfSrc1 : 5'h0; // @[src/main/scala/utils/PipelineVector.scala 45:69]
  wire [4:0] _dataBuffer_T_ctrl_rfSrc2 = needEnqueue_0 ? frontend_io_out_0_bits_ctrl_rfSrc2 : 5'h0; // @[src/main/scala/utils/PipelineVector.scala 45:69]
  wire [4:0] _dataBuffer_T_ctrl_rfDest = needEnqueue_0 ? frontend_io_out_0_bits_ctrl_rfDest : 5'h0; // @[src/main/scala/utils/PipelineVector.scala 45:69]
  wire [63:0] _dataBuffer_T_data_imm = needEnqueue_0 ? frontend_io_out_0_bits_data_imm : 64'h0; // @[src/main/scala/utils/PipelineVector.scala 45:69]
  wire [63:0] _GEN_0 = 2'h0 == _T_1[1:0] ? _dataBuffer_T_cf_instr : dataBuffer_0_cf_instr; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire [63:0] _GEN_1 = 2'h1 == _T_1[1:0] ? _dataBuffer_T_cf_instr : dataBuffer_1_cf_instr; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire [63:0] _GEN_2 = 2'h2 == _T_1[1:0] ? _dataBuffer_T_cf_instr : dataBuffer_2_cf_instr; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire [63:0] _GEN_3 = 2'h3 == _T_1[1:0] ? _dataBuffer_T_cf_instr : dataBuffer_3_cf_instr; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire [38:0] _GEN_4 = 2'h0 == _T_1[1:0] ? _dataBuffer_T_cf_pc : dataBuffer_0_cf_pc; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire [38:0] _GEN_5 = 2'h1 == _T_1[1:0] ? _dataBuffer_T_cf_pc : dataBuffer_1_cf_pc; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire [38:0] _GEN_6 = 2'h2 == _T_1[1:0] ? _dataBuffer_T_cf_pc : dataBuffer_2_cf_pc; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire [38:0] _GEN_7 = 2'h3 == _T_1[1:0] ? _dataBuffer_T_cf_pc : dataBuffer_3_cf_pc; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire [38:0] _GEN_8 = 2'h0 == _T_1[1:0] ? _dataBuffer_T_cf_pnpc : dataBuffer_0_cf_pnpc; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire [38:0] _GEN_9 = 2'h1 == _T_1[1:0] ? _dataBuffer_T_cf_pnpc : dataBuffer_1_cf_pnpc; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire [38:0] _GEN_10 = 2'h2 == _T_1[1:0] ? _dataBuffer_T_cf_pnpc : dataBuffer_2_cf_pnpc; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire [38:0] _GEN_11 = 2'h3 == _T_1[1:0] ? _dataBuffer_T_cf_pnpc : dataBuffer_3_cf_pnpc; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_28 = 2'h0 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_cf_exceptionVec_1 :
    dataBuffer_0_cf_exceptionVec_1; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_29 = 2'h1 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_cf_exceptionVec_1 :
    dataBuffer_1_cf_exceptionVec_1; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_30 = 2'h2 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_cf_exceptionVec_1 :
    dataBuffer_2_cf_exceptionVec_1; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_31 = 2'h3 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_cf_exceptionVec_1 :
    dataBuffer_3_cf_exceptionVec_1; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_32 = 2'h0 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_cf_exceptionVec_2 :
    dataBuffer_0_cf_exceptionVec_2; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_33 = 2'h1 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_cf_exceptionVec_2 :
    dataBuffer_1_cf_exceptionVec_2; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_34 = 2'h2 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_cf_exceptionVec_2 :
    dataBuffer_2_cf_exceptionVec_2; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_35 = 2'h3 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_cf_exceptionVec_2 :
    dataBuffer_3_cf_exceptionVec_2; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_72 = 2'h0 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_cf_exceptionVec_12 :
    dataBuffer_0_cf_exceptionVec_12; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_73 = 2'h1 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_cf_exceptionVec_12 :
    dataBuffer_1_cf_exceptionVec_12; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_74 = 2'h2 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_cf_exceptionVec_12 :
    dataBuffer_2_cf_exceptionVec_12; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_75 = 2'h3 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_cf_exceptionVec_12 :
    dataBuffer_3_cf_exceptionVec_12; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_88 = 2'h0 == _T_1[1:0] ? _dataBuffer_T_cf_intrVec_0 : dataBuffer_0_cf_intrVec_0; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_89 = 2'h1 == _T_1[1:0] ? _dataBuffer_T_cf_intrVec_0 : dataBuffer_1_cf_intrVec_0; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_90 = 2'h2 == _T_1[1:0] ? _dataBuffer_T_cf_intrVec_0 : dataBuffer_2_cf_intrVec_0; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_91 = 2'h3 == _T_1[1:0] ? _dataBuffer_T_cf_intrVec_0 : dataBuffer_3_cf_intrVec_0; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_92 = 2'h0 == _T_1[1:0] ? _dataBuffer_T_cf_intrVec_1 : dataBuffer_0_cf_intrVec_1; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_93 = 2'h1 == _T_1[1:0] ? _dataBuffer_T_cf_intrVec_1 : dataBuffer_1_cf_intrVec_1; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_94 = 2'h2 == _T_1[1:0] ? _dataBuffer_T_cf_intrVec_1 : dataBuffer_2_cf_intrVec_1; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_95 = 2'h3 == _T_1[1:0] ? _dataBuffer_T_cf_intrVec_1 : dataBuffer_3_cf_intrVec_1; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_96 = 2'h0 == _T_1[1:0] ? _dataBuffer_T_cf_intrVec_2 : dataBuffer_0_cf_intrVec_2; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_97 = 2'h1 == _T_1[1:0] ? _dataBuffer_T_cf_intrVec_2 : dataBuffer_1_cf_intrVec_2; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_98 = 2'h2 == _T_1[1:0] ? _dataBuffer_T_cf_intrVec_2 : dataBuffer_2_cf_intrVec_2; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_99 = 2'h3 == _T_1[1:0] ? _dataBuffer_T_cf_intrVec_2 : dataBuffer_3_cf_intrVec_2; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_100 = 2'h0 == _T_1[1:0] ? _dataBuffer_T_cf_intrVec_3 : dataBuffer_0_cf_intrVec_3; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_101 = 2'h1 == _T_1[1:0] ? _dataBuffer_T_cf_intrVec_3 : dataBuffer_1_cf_intrVec_3; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_102 = 2'h2 == _T_1[1:0] ? _dataBuffer_T_cf_intrVec_3 : dataBuffer_2_cf_intrVec_3; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_103 = 2'h3 == _T_1[1:0] ? _dataBuffer_T_cf_intrVec_3 : dataBuffer_3_cf_intrVec_3; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_104 = 2'h0 == _T_1[1:0] ? _dataBuffer_T_cf_intrVec_4 : dataBuffer_0_cf_intrVec_4; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_105 = 2'h1 == _T_1[1:0] ? _dataBuffer_T_cf_intrVec_4 : dataBuffer_1_cf_intrVec_4; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_106 = 2'h2 == _T_1[1:0] ? _dataBuffer_T_cf_intrVec_4 : dataBuffer_2_cf_intrVec_4; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_107 = 2'h3 == _T_1[1:0] ? _dataBuffer_T_cf_intrVec_4 : dataBuffer_3_cf_intrVec_4; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_108 = 2'h0 == _T_1[1:0] ? _dataBuffer_T_cf_intrVec_5 : dataBuffer_0_cf_intrVec_5; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_109 = 2'h1 == _T_1[1:0] ? _dataBuffer_T_cf_intrVec_5 : dataBuffer_1_cf_intrVec_5; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_110 = 2'h2 == _T_1[1:0] ? _dataBuffer_T_cf_intrVec_5 : dataBuffer_2_cf_intrVec_5; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_111 = 2'h3 == _T_1[1:0] ? _dataBuffer_T_cf_intrVec_5 : dataBuffer_3_cf_intrVec_5; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_112 = 2'h0 == _T_1[1:0] ? _dataBuffer_T_cf_intrVec_6 : dataBuffer_0_cf_intrVec_6; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_113 = 2'h1 == _T_1[1:0] ? _dataBuffer_T_cf_intrVec_6 : dataBuffer_1_cf_intrVec_6; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_114 = 2'h2 == _T_1[1:0] ? _dataBuffer_T_cf_intrVec_6 : dataBuffer_2_cf_intrVec_6; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_115 = 2'h3 == _T_1[1:0] ? _dataBuffer_T_cf_intrVec_6 : dataBuffer_3_cf_intrVec_6; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_116 = 2'h0 == _T_1[1:0] ? _dataBuffer_T_cf_intrVec_7 : dataBuffer_0_cf_intrVec_7; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_117 = 2'h1 == _T_1[1:0] ? _dataBuffer_T_cf_intrVec_7 : dataBuffer_1_cf_intrVec_7; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_118 = 2'h2 == _T_1[1:0] ? _dataBuffer_T_cf_intrVec_7 : dataBuffer_2_cf_intrVec_7; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_119 = 2'h3 == _T_1[1:0] ? _dataBuffer_T_cf_intrVec_7 : dataBuffer_3_cf_intrVec_7; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_120 = 2'h0 == _T_1[1:0] ? _dataBuffer_T_cf_intrVec_8 : dataBuffer_0_cf_intrVec_8; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_121 = 2'h1 == _T_1[1:0] ? _dataBuffer_T_cf_intrVec_8 : dataBuffer_1_cf_intrVec_8; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_122 = 2'h2 == _T_1[1:0] ? _dataBuffer_T_cf_intrVec_8 : dataBuffer_2_cf_intrVec_8; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_123 = 2'h3 == _T_1[1:0] ? _dataBuffer_T_cf_intrVec_8 : dataBuffer_3_cf_intrVec_8; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_124 = 2'h0 == _T_1[1:0] ? _dataBuffer_T_cf_intrVec_9 : dataBuffer_0_cf_intrVec_9; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_125 = 2'h1 == _T_1[1:0] ? _dataBuffer_T_cf_intrVec_9 : dataBuffer_1_cf_intrVec_9; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_126 = 2'h2 == _T_1[1:0] ? _dataBuffer_T_cf_intrVec_9 : dataBuffer_2_cf_intrVec_9; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_127 = 2'h3 == _T_1[1:0] ? _dataBuffer_T_cf_intrVec_9 : dataBuffer_3_cf_intrVec_9; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_128 = 2'h0 == _T_1[1:0] ? _dataBuffer_T_cf_intrVec_10 : dataBuffer_0_cf_intrVec_10; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_129 = 2'h1 == _T_1[1:0] ? _dataBuffer_T_cf_intrVec_10 : dataBuffer_1_cf_intrVec_10; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_130 = 2'h2 == _T_1[1:0] ? _dataBuffer_T_cf_intrVec_10 : dataBuffer_2_cf_intrVec_10; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_131 = 2'h3 == _T_1[1:0] ? _dataBuffer_T_cf_intrVec_10 : dataBuffer_3_cf_intrVec_10; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_132 = 2'h0 == _T_1[1:0] ? _dataBuffer_T_cf_intrVec_11 : dataBuffer_0_cf_intrVec_11; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_133 = 2'h1 == _T_1[1:0] ? _dataBuffer_T_cf_intrVec_11 : dataBuffer_1_cf_intrVec_11; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_134 = 2'h2 == _T_1[1:0] ? _dataBuffer_T_cf_intrVec_11 : dataBuffer_2_cf_intrVec_11; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_135 = 2'h3 == _T_1[1:0] ? _dataBuffer_T_cf_intrVec_11 : dataBuffer_3_cf_intrVec_11; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire [3:0] _GEN_136 = 2'h0 == _T_1[1:0] ? _dataBuffer_T_cf_brIdx : dataBuffer_0_cf_brIdx; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire [3:0] _GEN_137 = 2'h1 == _T_1[1:0] ? _dataBuffer_T_cf_brIdx : dataBuffer_1_cf_brIdx; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire [3:0] _GEN_138 = 2'h2 == _T_1[1:0] ? _dataBuffer_T_cf_brIdx : dataBuffer_2_cf_brIdx; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire [3:0] _GEN_139 = 2'h3 == _T_1[1:0] ? _dataBuffer_T_cf_brIdx : dataBuffer_3_cf_brIdx; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_144 = 2'h0 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_cf_crossPageIPFFix :
    dataBuffer_0_cf_crossPageIPFFix; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_145 = 2'h1 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_cf_crossPageIPFFix :
    dataBuffer_1_cf_crossPageIPFFix; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_146 = 2'h2 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_cf_crossPageIPFFix :
    dataBuffer_2_cf_crossPageIPFFix; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_147 = 2'h3 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_cf_crossPageIPFFix :
    dataBuffer_3_cf_crossPageIPFFix; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_156 = 2'h0 == _T_1[1:0] ? _dataBuffer_T_ctrl_src1Type : dataBuffer_0_ctrl_src1Type; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_157 = 2'h1 == _T_1[1:0] ? _dataBuffer_T_ctrl_src1Type : dataBuffer_1_ctrl_src1Type; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_158 = 2'h2 == _T_1[1:0] ? _dataBuffer_T_ctrl_src1Type : dataBuffer_2_ctrl_src1Type; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_159 = 2'h3 == _T_1[1:0] ? _dataBuffer_T_ctrl_src1Type : dataBuffer_3_ctrl_src1Type; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_160 = 2'h0 == _T_1[1:0] ? _dataBuffer_T_ctrl_src2Type : dataBuffer_0_ctrl_src2Type; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_161 = 2'h1 == _T_1[1:0] ? _dataBuffer_T_ctrl_src2Type : dataBuffer_1_ctrl_src2Type; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_162 = 2'h2 == _T_1[1:0] ? _dataBuffer_T_ctrl_src2Type : dataBuffer_2_ctrl_src2Type; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_163 = 2'h3 == _T_1[1:0] ? _dataBuffer_T_ctrl_src2Type : dataBuffer_3_ctrl_src2Type; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire [2:0] _GEN_164 = 2'h0 == _T_1[1:0] ? _dataBuffer_T_ctrl_fuType : dataBuffer_0_ctrl_fuType; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire [2:0] _GEN_165 = 2'h1 == _T_1[1:0] ? _dataBuffer_T_ctrl_fuType : dataBuffer_1_ctrl_fuType; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire [2:0] _GEN_166 = 2'h2 == _T_1[1:0] ? _dataBuffer_T_ctrl_fuType : dataBuffer_2_ctrl_fuType; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire [2:0] _GEN_167 = 2'h3 == _T_1[1:0] ? _dataBuffer_T_ctrl_fuType : dataBuffer_3_ctrl_fuType; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire [6:0] _GEN_168 = 2'h0 == _T_1[1:0] ? _dataBuffer_T_ctrl_fuOpType : dataBuffer_0_ctrl_fuOpType; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire [6:0] _GEN_169 = 2'h1 == _T_1[1:0] ? _dataBuffer_T_ctrl_fuOpType : dataBuffer_1_ctrl_fuOpType; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire [6:0] _GEN_170 = 2'h2 == _T_1[1:0] ? _dataBuffer_T_ctrl_fuOpType : dataBuffer_2_ctrl_fuOpType; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire [6:0] _GEN_171 = 2'h3 == _T_1[1:0] ? _dataBuffer_T_ctrl_fuOpType : dataBuffer_3_ctrl_fuOpType; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire [4:0] _GEN_172 = 2'h0 == _T_1[1:0] ? _dataBuffer_T_ctrl_rfSrc1 : dataBuffer_0_ctrl_rfSrc1; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire [4:0] _GEN_173 = 2'h1 == _T_1[1:0] ? _dataBuffer_T_ctrl_rfSrc1 : dataBuffer_1_ctrl_rfSrc1; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire [4:0] _GEN_174 = 2'h2 == _T_1[1:0] ? _dataBuffer_T_ctrl_rfSrc1 : dataBuffer_2_ctrl_rfSrc1; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire [4:0] _GEN_175 = 2'h3 == _T_1[1:0] ? _dataBuffer_T_ctrl_rfSrc1 : dataBuffer_3_ctrl_rfSrc1; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire [4:0] _GEN_176 = 2'h0 == _T_1[1:0] ? _dataBuffer_T_ctrl_rfSrc2 : dataBuffer_0_ctrl_rfSrc2; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire [4:0] _GEN_177 = 2'h1 == _T_1[1:0] ? _dataBuffer_T_ctrl_rfSrc2 : dataBuffer_1_ctrl_rfSrc2; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire [4:0] _GEN_178 = 2'h2 == _T_1[1:0] ? _dataBuffer_T_ctrl_rfSrc2 : dataBuffer_2_ctrl_rfSrc2; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire [4:0] _GEN_179 = 2'h3 == _T_1[1:0] ? _dataBuffer_T_ctrl_rfSrc2 : dataBuffer_3_ctrl_rfSrc2; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_180 = 2'h0 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_ctrl_rfWen : dataBuffer_0_ctrl_rfWen; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_181 = 2'h1 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_ctrl_rfWen : dataBuffer_1_ctrl_rfWen; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_182 = 2'h2 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_ctrl_rfWen : dataBuffer_2_ctrl_rfWen; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_183 = 2'h3 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_ctrl_rfWen : dataBuffer_3_ctrl_rfWen; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire [4:0] _GEN_184 = 2'h0 == _T_1[1:0] ? _dataBuffer_T_ctrl_rfDest : dataBuffer_0_ctrl_rfDest; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire [4:0] _GEN_185 = 2'h1 == _T_1[1:0] ? _dataBuffer_T_ctrl_rfDest : dataBuffer_1_ctrl_rfDest; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire [4:0] _GEN_186 = 2'h2 == _T_1[1:0] ? _dataBuffer_T_ctrl_rfDest : dataBuffer_2_ctrl_rfDest; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire [4:0] _GEN_187 = 2'h3 == _T_1[1:0] ? _dataBuffer_T_ctrl_rfDest : dataBuffer_3_ctrl_rfDest; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_188 = 2'h0 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_ctrl_isNutCoreTrap :
    dataBuffer_0_ctrl_isNutCoreTrap; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_189 = 2'h1 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_ctrl_isNutCoreTrap :
    dataBuffer_1_ctrl_isNutCoreTrap; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_190 = 2'h2 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_ctrl_isNutCoreTrap :
    dataBuffer_2_ctrl_isNutCoreTrap; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_191 = 2'h3 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_ctrl_isNutCoreTrap :
    dataBuffer_3_ctrl_isNutCoreTrap; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire [63:0] _GEN_216 = 2'h0 == _T_1[1:0] ? _dataBuffer_T_data_imm : dataBuffer_0_data_imm; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire [63:0] _GEN_217 = 2'h1 == _T_1[1:0] ? _dataBuffer_T_data_imm : dataBuffer_1_data_imm; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire [63:0] _GEN_218 = 2'h2 == _T_1[1:0] ? _dataBuffer_T_data_imm : dataBuffer_2_data_imm; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire [63:0] _GEN_219 = 2'h3 == _T_1[1:0] ? _dataBuffer_T_data_imm : dataBuffer_3_data_imm; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire [63:0] _GEN_220 = enqueueFire_0 ? _GEN_0 : dataBuffer_0_cf_instr; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [63:0] _GEN_221 = enqueueFire_0 ? _GEN_1 : dataBuffer_1_cf_instr; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [63:0] _GEN_222 = enqueueFire_0 ? _GEN_2 : dataBuffer_2_cf_instr; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [63:0] _GEN_223 = enqueueFire_0 ? _GEN_3 : dataBuffer_3_cf_instr; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [38:0] _GEN_224 = enqueueFire_0 ? _GEN_4 : dataBuffer_0_cf_pc; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [38:0] _GEN_225 = enqueueFire_0 ? _GEN_5 : dataBuffer_1_cf_pc; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [38:0] _GEN_226 = enqueueFire_0 ? _GEN_6 : dataBuffer_2_cf_pc; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [38:0] _GEN_227 = enqueueFire_0 ? _GEN_7 : dataBuffer_3_cf_pc; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [38:0] _GEN_228 = enqueueFire_0 ? _GEN_8 : dataBuffer_0_cf_pnpc; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [38:0] _GEN_229 = enqueueFire_0 ? _GEN_9 : dataBuffer_1_cf_pnpc; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [38:0] _GEN_230 = enqueueFire_0 ? _GEN_10 : dataBuffer_2_cf_pnpc; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [38:0] _GEN_231 = enqueueFire_0 ? _GEN_11 : dataBuffer_3_cf_pnpc; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_248 = enqueueFire_0 ? _GEN_28 : dataBuffer_0_cf_exceptionVec_1; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_249 = enqueueFire_0 ? _GEN_29 : dataBuffer_1_cf_exceptionVec_1; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_250 = enqueueFire_0 ? _GEN_30 : dataBuffer_2_cf_exceptionVec_1; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_251 = enqueueFire_0 ? _GEN_31 : dataBuffer_3_cf_exceptionVec_1; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_252 = enqueueFire_0 ? _GEN_32 : dataBuffer_0_cf_exceptionVec_2; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_253 = enqueueFire_0 ? _GEN_33 : dataBuffer_1_cf_exceptionVec_2; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_254 = enqueueFire_0 ? _GEN_34 : dataBuffer_2_cf_exceptionVec_2; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_255 = enqueueFire_0 ? _GEN_35 : dataBuffer_3_cf_exceptionVec_2; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_292 = enqueueFire_0 ? _GEN_72 : dataBuffer_0_cf_exceptionVec_12; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_293 = enqueueFire_0 ? _GEN_73 : dataBuffer_1_cf_exceptionVec_12; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_294 = enqueueFire_0 ? _GEN_74 : dataBuffer_2_cf_exceptionVec_12; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_295 = enqueueFire_0 ? _GEN_75 : dataBuffer_3_cf_exceptionVec_12; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_308 = enqueueFire_0 ? _GEN_88 : dataBuffer_0_cf_intrVec_0; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_309 = enqueueFire_0 ? _GEN_89 : dataBuffer_1_cf_intrVec_0; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_310 = enqueueFire_0 ? _GEN_90 : dataBuffer_2_cf_intrVec_0; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_311 = enqueueFire_0 ? _GEN_91 : dataBuffer_3_cf_intrVec_0; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_312 = enqueueFire_0 ? _GEN_92 : dataBuffer_0_cf_intrVec_1; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_313 = enqueueFire_0 ? _GEN_93 : dataBuffer_1_cf_intrVec_1; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_314 = enqueueFire_0 ? _GEN_94 : dataBuffer_2_cf_intrVec_1; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_315 = enqueueFire_0 ? _GEN_95 : dataBuffer_3_cf_intrVec_1; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_316 = enqueueFire_0 ? _GEN_96 : dataBuffer_0_cf_intrVec_2; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_317 = enqueueFire_0 ? _GEN_97 : dataBuffer_1_cf_intrVec_2; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_318 = enqueueFire_0 ? _GEN_98 : dataBuffer_2_cf_intrVec_2; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_319 = enqueueFire_0 ? _GEN_99 : dataBuffer_3_cf_intrVec_2; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_320 = enqueueFire_0 ? _GEN_100 : dataBuffer_0_cf_intrVec_3; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_321 = enqueueFire_0 ? _GEN_101 : dataBuffer_1_cf_intrVec_3; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_322 = enqueueFire_0 ? _GEN_102 : dataBuffer_2_cf_intrVec_3; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_323 = enqueueFire_0 ? _GEN_103 : dataBuffer_3_cf_intrVec_3; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_324 = enqueueFire_0 ? _GEN_104 : dataBuffer_0_cf_intrVec_4; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_325 = enqueueFire_0 ? _GEN_105 : dataBuffer_1_cf_intrVec_4; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_326 = enqueueFire_0 ? _GEN_106 : dataBuffer_2_cf_intrVec_4; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_327 = enqueueFire_0 ? _GEN_107 : dataBuffer_3_cf_intrVec_4; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_328 = enqueueFire_0 ? _GEN_108 : dataBuffer_0_cf_intrVec_5; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_329 = enqueueFire_0 ? _GEN_109 : dataBuffer_1_cf_intrVec_5; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_330 = enqueueFire_0 ? _GEN_110 : dataBuffer_2_cf_intrVec_5; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_331 = enqueueFire_0 ? _GEN_111 : dataBuffer_3_cf_intrVec_5; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_332 = enqueueFire_0 ? _GEN_112 : dataBuffer_0_cf_intrVec_6; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_333 = enqueueFire_0 ? _GEN_113 : dataBuffer_1_cf_intrVec_6; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_334 = enqueueFire_0 ? _GEN_114 : dataBuffer_2_cf_intrVec_6; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_335 = enqueueFire_0 ? _GEN_115 : dataBuffer_3_cf_intrVec_6; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_336 = enqueueFire_0 ? _GEN_116 : dataBuffer_0_cf_intrVec_7; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_337 = enqueueFire_0 ? _GEN_117 : dataBuffer_1_cf_intrVec_7; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_338 = enqueueFire_0 ? _GEN_118 : dataBuffer_2_cf_intrVec_7; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_339 = enqueueFire_0 ? _GEN_119 : dataBuffer_3_cf_intrVec_7; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_340 = enqueueFire_0 ? _GEN_120 : dataBuffer_0_cf_intrVec_8; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_341 = enqueueFire_0 ? _GEN_121 : dataBuffer_1_cf_intrVec_8; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_342 = enqueueFire_0 ? _GEN_122 : dataBuffer_2_cf_intrVec_8; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_343 = enqueueFire_0 ? _GEN_123 : dataBuffer_3_cf_intrVec_8; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_344 = enqueueFire_0 ? _GEN_124 : dataBuffer_0_cf_intrVec_9; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_345 = enqueueFire_0 ? _GEN_125 : dataBuffer_1_cf_intrVec_9; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_346 = enqueueFire_0 ? _GEN_126 : dataBuffer_2_cf_intrVec_9; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_347 = enqueueFire_0 ? _GEN_127 : dataBuffer_3_cf_intrVec_9; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_348 = enqueueFire_0 ? _GEN_128 : dataBuffer_0_cf_intrVec_10; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_349 = enqueueFire_0 ? _GEN_129 : dataBuffer_1_cf_intrVec_10; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_350 = enqueueFire_0 ? _GEN_130 : dataBuffer_2_cf_intrVec_10; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_351 = enqueueFire_0 ? _GEN_131 : dataBuffer_3_cf_intrVec_10; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_352 = enqueueFire_0 ? _GEN_132 : dataBuffer_0_cf_intrVec_11; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_353 = enqueueFire_0 ? _GEN_133 : dataBuffer_1_cf_intrVec_11; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_354 = enqueueFire_0 ? _GEN_134 : dataBuffer_2_cf_intrVec_11; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_355 = enqueueFire_0 ? _GEN_135 : dataBuffer_3_cf_intrVec_11; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [3:0] _GEN_356 = enqueueFire_0 ? _GEN_136 : dataBuffer_0_cf_brIdx; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [3:0] _GEN_357 = enqueueFire_0 ? _GEN_137 : dataBuffer_1_cf_brIdx; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [3:0] _GEN_358 = enqueueFire_0 ? _GEN_138 : dataBuffer_2_cf_brIdx; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [3:0] _GEN_359 = enqueueFire_0 ? _GEN_139 : dataBuffer_3_cf_brIdx; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_364 = enqueueFire_0 ? _GEN_144 : dataBuffer_0_cf_crossPageIPFFix; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_365 = enqueueFire_0 ? _GEN_145 : dataBuffer_1_cf_crossPageIPFFix; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_366 = enqueueFire_0 ? _GEN_146 : dataBuffer_2_cf_crossPageIPFFix; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_367 = enqueueFire_0 ? _GEN_147 : dataBuffer_3_cf_crossPageIPFFix; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_376 = enqueueFire_0 ? _GEN_156 : dataBuffer_0_ctrl_src1Type; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_377 = enqueueFire_0 ? _GEN_157 : dataBuffer_1_ctrl_src1Type; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_378 = enqueueFire_0 ? _GEN_158 : dataBuffer_2_ctrl_src1Type; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_379 = enqueueFire_0 ? _GEN_159 : dataBuffer_3_ctrl_src1Type; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_380 = enqueueFire_0 ? _GEN_160 : dataBuffer_0_ctrl_src2Type; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_381 = enqueueFire_0 ? _GEN_161 : dataBuffer_1_ctrl_src2Type; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_382 = enqueueFire_0 ? _GEN_162 : dataBuffer_2_ctrl_src2Type; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_383 = enqueueFire_0 ? _GEN_163 : dataBuffer_3_ctrl_src2Type; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [2:0] _GEN_384 = enqueueFire_0 ? _GEN_164 : dataBuffer_0_ctrl_fuType; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [2:0] _GEN_385 = enqueueFire_0 ? _GEN_165 : dataBuffer_1_ctrl_fuType; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [2:0] _GEN_386 = enqueueFire_0 ? _GEN_166 : dataBuffer_2_ctrl_fuType; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [2:0] _GEN_387 = enqueueFire_0 ? _GEN_167 : dataBuffer_3_ctrl_fuType; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [6:0] _GEN_388 = enqueueFire_0 ? _GEN_168 : dataBuffer_0_ctrl_fuOpType; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [6:0] _GEN_389 = enqueueFire_0 ? _GEN_169 : dataBuffer_1_ctrl_fuOpType; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [6:0] _GEN_390 = enqueueFire_0 ? _GEN_170 : dataBuffer_2_ctrl_fuOpType; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [6:0] _GEN_391 = enqueueFire_0 ? _GEN_171 : dataBuffer_3_ctrl_fuOpType; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [4:0] _GEN_392 = enqueueFire_0 ? _GEN_172 : dataBuffer_0_ctrl_rfSrc1; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [4:0] _GEN_393 = enqueueFire_0 ? _GEN_173 : dataBuffer_1_ctrl_rfSrc1; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [4:0] _GEN_394 = enqueueFire_0 ? _GEN_174 : dataBuffer_2_ctrl_rfSrc1; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [4:0] _GEN_395 = enqueueFire_0 ? _GEN_175 : dataBuffer_3_ctrl_rfSrc1; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [4:0] _GEN_396 = enqueueFire_0 ? _GEN_176 : dataBuffer_0_ctrl_rfSrc2; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [4:0] _GEN_397 = enqueueFire_0 ? _GEN_177 : dataBuffer_1_ctrl_rfSrc2; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [4:0] _GEN_398 = enqueueFire_0 ? _GEN_178 : dataBuffer_2_ctrl_rfSrc2; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [4:0] _GEN_399 = enqueueFire_0 ? _GEN_179 : dataBuffer_3_ctrl_rfSrc2; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_400 = enqueueFire_0 ? _GEN_180 : dataBuffer_0_ctrl_rfWen; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_401 = enqueueFire_0 ? _GEN_181 : dataBuffer_1_ctrl_rfWen; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_402 = enqueueFire_0 ? _GEN_182 : dataBuffer_2_ctrl_rfWen; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_403 = enqueueFire_0 ? _GEN_183 : dataBuffer_3_ctrl_rfWen; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [4:0] _GEN_404 = enqueueFire_0 ? _GEN_184 : dataBuffer_0_ctrl_rfDest; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [4:0] _GEN_405 = enqueueFire_0 ? _GEN_185 : dataBuffer_1_ctrl_rfDest; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [4:0] _GEN_406 = enqueueFire_0 ? _GEN_186 : dataBuffer_2_ctrl_rfDest; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [4:0] _GEN_407 = enqueueFire_0 ? _GEN_187 : dataBuffer_3_ctrl_rfDest; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_408 = enqueueFire_0 ? _GEN_188 : dataBuffer_0_ctrl_isNutCoreTrap; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_409 = enqueueFire_0 ? _GEN_189 : dataBuffer_1_ctrl_isNutCoreTrap; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_410 = enqueueFire_0 ? _GEN_190 : dataBuffer_2_ctrl_isNutCoreTrap; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_411 = enqueueFire_0 ? _GEN_191 : dataBuffer_3_ctrl_isNutCoreTrap; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [63:0] _GEN_436 = enqueueFire_0 ? _GEN_216 : dataBuffer_0_data_imm; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [63:0] _GEN_437 = enqueueFire_0 ? _GEN_217 : dataBuffer_1_data_imm; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [63:0] _GEN_438 = enqueueFire_0 ? _GEN_218 : dataBuffer_2_data_imm; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [63:0] _GEN_439 = enqueueFire_0 ? _GEN_219 : dataBuffer_3_data_imm; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [1:0] _T_4 = 2'h1 + ringBufferHead; // @[src/main/scala/utils/PipelineVector.scala 46:45]
  wire [1:0] _ringBufferHead_T_1 = ringBufferHead + enqueueSize; // @[src/main/scala/utils/PipelineVector.scala 47:42]
  wire [63:0] _GEN_1102 = 2'h1 == ringBufferTail ? dataBuffer_1_data_imm : dataBuffer_0_data_imm; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire [63:0] _GEN_1103 = 2'h2 == ringBufferTail ? dataBuffer_2_data_imm : _GEN_1102; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire  _GEN_1130 = 2'h1 == ringBufferTail ? dataBuffer_1_ctrl_isNutCoreTrap : dataBuffer_0_ctrl_isNutCoreTrap; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire  _GEN_1131 = 2'h2 == ringBufferTail ? dataBuffer_2_ctrl_isNutCoreTrap : _GEN_1130; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire [4:0] _GEN_1134 = 2'h1 == ringBufferTail ? dataBuffer_1_ctrl_rfDest : dataBuffer_0_ctrl_rfDest; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire [4:0] _GEN_1135 = 2'h2 == ringBufferTail ? dataBuffer_2_ctrl_rfDest : _GEN_1134; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire  _GEN_1138 = 2'h1 == ringBufferTail ? dataBuffer_1_ctrl_rfWen : dataBuffer_0_ctrl_rfWen; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire  _GEN_1139 = 2'h2 == ringBufferTail ? dataBuffer_2_ctrl_rfWen : _GEN_1138; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire [4:0] _GEN_1142 = 2'h1 == ringBufferTail ? dataBuffer_1_ctrl_rfSrc2 : dataBuffer_0_ctrl_rfSrc2; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire [4:0] _GEN_1143 = 2'h2 == ringBufferTail ? dataBuffer_2_ctrl_rfSrc2 : _GEN_1142; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire [4:0] _GEN_1146 = 2'h1 == ringBufferTail ? dataBuffer_1_ctrl_rfSrc1 : dataBuffer_0_ctrl_rfSrc1; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire [4:0] _GEN_1147 = 2'h2 == ringBufferTail ? dataBuffer_2_ctrl_rfSrc1 : _GEN_1146; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire [6:0] _GEN_1150 = 2'h1 == ringBufferTail ? dataBuffer_1_ctrl_fuOpType : dataBuffer_0_ctrl_fuOpType; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire [6:0] _GEN_1151 = 2'h2 == ringBufferTail ? dataBuffer_2_ctrl_fuOpType : _GEN_1150; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire [2:0] _GEN_1154 = 2'h1 == ringBufferTail ? dataBuffer_1_ctrl_fuType : dataBuffer_0_ctrl_fuType; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire [2:0] _GEN_1155 = 2'h2 == ringBufferTail ? dataBuffer_2_ctrl_fuType : _GEN_1154; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire  _GEN_1158 = 2'h1 == ringBufferTail ? dataBuffer_1_ctrl_src2Type : dataBuffer_0_ctrl_src2Type; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire  _GEN_1159 = 2'h2 == ringBufferTail ? dataBuffer_2_ctrl_src2Type : _GEN_1158; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire  _GEN_1162 = 2'h1 == ringBufferTail ? dataBuffer_1_ctrl_src1Type : dataBuffer_0_ctrl_src1Type; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire  _GEN_1163 = 2'h2 == ringBufferTail ? dataBuffer_2_ctrl_src1Type : _GEN_1162; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire  _GEN_1174 = 2'h1 == ringBufferTail ? dataBuffer_1_cf_crossPageIPFFix : dataBuffer_0_cf_crossPageIPFFix; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire  _GEN_1175 = 2'h2 == ringBufferTail ? dataBuffer_2_cf_crossPageIPFFix : _GEN_1174; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire [3:0] _GEN_1182 = 2'h1 == ringBufferTail ? dataBuffer_1_cf_brIdx : dataBuffer_0_cf_brIdx; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire [3:0] _GEN_1183 = 2'h2 == ringBufferTail ? dataBuffer_2_cf_brIdx : _GEN_1182; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire  _GEN_1186 = 2'h1 == ringBufferTail ? dataBuffer_1_cf_intrVec_0 : dataBuffer_0_cf_intrVec_0; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire  _GEN_1187 = 2'h2 == ringBufferTail ? dataBuffer_2_cf_intrVec_0 : _GEN_1186; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire  _GEN_1190 = 2'h1 == ringBufferTail ? dataBuffer_1_cf_intrVec_1 : dataBuffer_0_cf_intrVec_1; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire  _GEN_1191 = 2'h2 == ringBufferTail ? dataBuffer_2_cf_intrVec_1 : _GEN_1190; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire  _GEN_1194 = 2'h1 == ringBufferTail ? dataBuffer_1_cf_intrVec_2 : dataBuffer_0_cf_intrVec_2; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire  _GEN_1195 = 2'h2 == ringBufferTail ? dataBuffer_2_cf_intrVec_2 : _GEN_1194; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire  _GEN_1198 = 2'h1 == ringBufferTail ? dataBuffer_1_cf_intrVec_3 : dataBuffer_0_cf_intrVec_3; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire  _GEN_1199 = 2'h2 == ringBufferTail ? dataBuffer_2_cf_intrVec_3 : _GEN_1198; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire  _GEN_1202 = 2'h1 == ringBufferTail ? dataBuffer_1_cf_intrVec_4 : dataBuffer_0_cf_intrVec_4; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire  _GEN_1203 = 2'h2 == ringBufferTail ? dataBuffer_2_cf_intrVec_4 : _GEN_1202; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire  _GEN_1206 = 2'h1 == ringBufferTail ? dataBuffer_1_cf_intrVec_5 : dataBuffer_0_cf_intrVec_5; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire  _GEN_1207 = 2'h2 == ringBufferTail ? dataBuffer_2_cf_intrVec_5 : _GEN_1206; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire  _GEN_1210 = 2'h1 == ringBufferTail ? dataBuffer_1_cf_intrVec_6 : dataBuffer_0_cf_intrVec_6; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire  _GEN_1211 = 2'h2 == ringBufferTail ? dataBuffer_2_cf_intrVec_6 : _GEN_1210; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire  _GEN_1214 = 2'h1 == ringBufferTail ? dataBuffer_1_cf_intrVec_7 : dataBuffer_0_cf_intrVec_7; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire  _GEN_1215 = 2'h2 == ringBufferTail ? dataBuffer_2_cf_intrVec_7 : _GEN_1214; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire  _GEN_1218 = 2'h1 == ringBufferTail ? dataBuffer_1_cf_intrVec_8 : dataBuffer_0_cf_intrVec_8; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire  _GEN_1219 = 2'h2 == ringBufferTail ? dataBuffer_2_cf_intrVec_8 : _GEN_1218; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire  _GEN_1222 = 2'h1 == ringBufferTail ? dataBuffer_1_cf_intrVec_9 : dataBuffer_0_cf_intrVec_9; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire  _GEN_1223 = 2'h2 == ringBufferTail ? dataBuffer_2_cf_intrVec_9 : _GEN_1222; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire  _GEN_1226 = 2'h1 == ringBufferTail ? dataBuffer_1_cf_intrVec_10 : dataBuffer_0_cf_intrVec_10; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire  _GEN_1227 = 2'h2 == ringBufferTail ? dataBuffer_2_cf_intrVec_10 : _GEN_1226; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire  _GEN_1230 = 2'h1 == ringBufferTail ? dataBuffer_1_cf_intrVec_11 : dataBuffer_0_cf_intrVec_11; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire  _GEN_1231 = 2'h2 == ringBufferTail ? dataBuffer_2_cf_intrVec_11 : _GEN_1230; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire  _GEN_1238 = 2'h1 == ringBufferTail ? dataBuffer_1_cf_exceptionVec_1 : dataBuffer_0_cf_exceptionVec_1; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire  _GEN_1239 = 2'h2 == ringBufferTail ? dataBuffer_2_cf_exceptionVec_1 : _GEN_1238; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire  _GEN_1242 = 2'h1 == ringBufferTail ? dataBuffer_1_cf_exceptionVec_2 : dataBuffer_0_cf_exceptionVec_2; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire  _GEN_1243 = 2'h2 == ringBufferTail ? dataBuffer_2_cf_exceptionVec_2 : _GEN_1242; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire  _GEN_1282 = 2'h1 == ringBufferTail ? dataBuffer_1_cf_exceptionVec_12 : dataBuffer_0_cf_exceptionVec_12; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire  _GEN_1283 = 2'h2 == ringBufferTail ? dataBuffer_2_cf_exceptionVec_12 : _GEN_1282; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire [38:0] _GEN_1310 = 2'h1 == ringBufferTail ? dataBuffer_1_cf_pnpc : dataBuffer_0_cf_pnpc; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire [38:0] _GEN_1311 = 2'h2 == ringBufferTail ? dataBuffer_2_cf_pnpc : _GEN_1310; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire [38:0] _GEN_1314 = 2'h1 == ringBufferTail ? dataBuffer_1_cf_pc : dataBuffer_0_cf_pc; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire [38:0] _GEN_1315 = 2'h2 == ringBufferTail ? dataBuffer_2_cf_pc : _GEN_1314; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire [63:0] _GEN_1318 = 2'h1 == ringBufferTail ? dataBuffer_1_cf_instr : dataBuffer_0_cf_instr; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire [63:0] _GEN_1319 = 2'h2 == ringBufferTail ? dataBuffer_2_cf_instr : _GEN_1318; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire  _dequeueSize_T = backend_io_in_0_ready & backend_io_in_0_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  wire [1:0] dequeueSize = {{1'd0}, _dequeueSize_T}; // @[src/main/scala/utils/PipelineVector.scala 64:40]
  wire  dequeueFire = dequeueSize > 2'h0; // @[src/main/scala/utils/PipelineVector.scala 65:35]
  wire [1:0] _ringBufferTail_T_1 = ringBufferTail + dequeueSize; // @[src/main/scala/utils/PipelineVector.scala 67:42]
  wire [3:0] _T_6 = 3'h4 + _T_1; // @[src/main/scala/utils/PipelineVector.scala 77:84]
  wire [3:0] _GEN_1553 = {{2'd0}, ringBufferTail}; // @[src/main/scala/utils/PipelineVector.scala 77:109]
  wire [3:0] _T_8 = _T_6 - _GEN_1553; // @[src/main/scala/utils/PipelineVector.scala 77:109]
  wire [3:0] _GEN_12 = _T_8 % 4'h4; // @[src/main/scala/utils/PipelineVector.scala 77:134]
  wire  _T_11 = ~reset; // @[src/main/scala/utils/PipelineVector.scala 77:15]
  reg [63:0] c; // @[src/main/scala/utils/GTimer.scala 24:20]
  wire [63:0] _c_T_1 = c + 64'h1; // @[src/main/scala/utils/GTimer.scala 25:12]
  Frontend_inorder frontend ( // @[src/main/scala/nutcore/NutCore.scala 104:34]
    .clock(frontend_clock),
    .reset(frontend_reset),
    .io_imem_req_ready(frontend_io_imem_req_ready),
    .io_imem_req_valid(frontend_io_imem_req_valid),
    .io_imem_req_bits_addr(frontend_io_imem_req_bits_addr),
    .io_imem_req_bits_user(frontend_io_imem_req_bits_user),
    .io_imem_resp_ready(frontend_io_imem_resp_ready),
    .io_imem_resp_valid(frontend_io_imem_resp_valid),
    .io_imem_resp_bits_rdata(frontend_io_imem_resp_bits_rdata),
    .io_imem_resp_bits_user(frontend_io_imem_resp_bits_user),
    .io_out_0_ready(frontend_io_out_0_ready),
    .io_out_0_valid(frontend_io_out_0_valid),
    .io_out_0_bits_cf_instr(frontend_io_out_0_bits_cf_instr),
    .io_out_0_bits_cf_pc(frontend_io_out_0_bits_cf_pc),
    .io_out_0_bits_cf_pnpc(frontend_io_out_0_bits_cf_pnpc),
    .io_out_0_bits_cf_exceptionVec_1(frontend_io_out_0_bits_cf_exceptionVec_1),
    .io_out_0_bits_cf_exceptionVec_2(frontend_io_out_0_bits_cf_exceptionVec_2),
    .io_out_0_bits_cf_exceptionVec_12(frontend_io_out_0_bits_cf_exceptionVec_12),
    .io_out_0_bits_cf_intrVec_0(frontend_io_out_0_bits_cf_intrVec_0),
    .io_out_0_bits_cf_intrVec_1(frontend_io_out_0_bits_cf_intrVec_1),
    .io_out_0_bits_cf_intrVec_2(frontend_io_out_0_bits_cf_intrVec_2),
    .io_out_0_bits_cf_intrVec_3(frontend_io_out_0_bits_cf_intrVec_3),
    .io_out_0_bits_cf_intrVec_4(frontend_io_out_0_bits_cf_intrVec_4),
    .io_out_0_bits_cf_intrVec_5(frontend_io_out_0_bits_cf_intrVec_5),
    .io_out_0_bits_cf_intrVec_6(frontend_io_out_0_bits_cf_intrVec_6),
    .io_out_0_bits_cf_intrVec_7(frontend_io_out_0_bits_cf_intrVec_7),
    .io_out_0_bits_cf_intrVec_8(frontend_io_out_0_bits_cf_intrVec_8),
    .io_out_0_bits_cf_intrVec_9(frontend_io_out_0_bits_cf_intrVec_9),
    .io_out_0_bits_cf_intrVec_10(frontend_io_out_0_bits_cf_intrVec_10),
    .io_out_0_bits_cf_intrVec_11(frontend_io_out_0_bits_cf_intrVec_11),
    .io_out_0_bits_cf_brIdx(frontend_io_out_0_bits_cf_brIdx),
    .io_out_0_bits_cf_crossPageIPFFix(frontend_io_out_0_bits_cf_crossPageIPFFix),
    .io_out_0_bits_ctrl_src1Type(frontend_io_out_0_bits_ctrl_src1Type),
    .io_out_0_bits_ctrl_src2Type(frontend_io_out_0_bits_ctrl_src2Type),
    .io_out_0_bits_ctrl_fuType(frontend_io_out_0_bits_ctrl_fuType),
    .io_out_0_bits_ctrl_fuOpType(frontend_io_out_0_bits_ctrl_fuOpType),
    .io_out_0_bits_ctrl_rfSrc1(frontend_io_out_0_bits_ctrl_rfSrc1),
    .io_out_0_bits_ctrl_rfSrc2(frontend_io_out_0_bits_ctrl_rfSrc2),
    .io_out_0_bits_ctrl_rfWen(frontend_io_out_0_bits_ctrl_rfWen),
    .io_out_0_bits_ctrl_rfDest(frontend_io_out_0_bits_ctrl_rfDest),
    .io_out_0_bits_ctrl_isNutCoreTrap(frontend_io_out_0_bits_ctrl_isNutCoreTrap),
    .io_out_0_bits_data_imm(frontend_io_out_0_bits_data_imm),
    .io_out_1_bits_cf_intrVec_0(frontend_io_out_1_bits_cf_intrVec_0),
    .io_out_1_bits_cf_intrVec_1(frontend_io_out_1_bits_cf_intrVec_1),
    .io_out_1_bits_cf_intrVec_2(frontend_io_out_1_bits_cf_intrVec_2),
    .io_out_1_bits_cf_intrVec_3(frontend_io_out_1_bits_cf_intrVec_3),
    .io_out_1_bits_cf_intrVec_4(frontend_io_out_1_bits_cf_intrVec_4),
    .io_out_1_bits_cf_intrVec_5(frontend_io_out_1_bits_cf_intrVec_5),
    .io_out_1_bits_cf_intrVec_6(frontend_io_out_1_bits_cf_intrVec_6),
    .io_out_1_bits_cf_intrVec_7(frontend_io_out_1_bits_cf_intrVec_7),
    .io_out_1_bits_cf_intrVec_8(frontend_io_out_1_bits_cf_intrVec_8),
    .io_out_1_bits_cf_intrVec_9(frontend_io_out_1_bits_cf_intrVec_9),
    .io_out_1_bits_cf_intrVec_10(frontend_io_out_1_bits_cf_intrVec_10),
    .io_out_1_bits_cf_intrVec_11(frontend_io_out_1_bits_cf_intrVec_11),
    .io_flushVec(frontend_io_flushVec),
    .io_redirect_target(frontend_io_redirect_target),
    .io_redirect_valid(frontend_io_redirect_valid),
    .io_ipf(frontend_io_ipf),
    .REG_valid(frontend_REG_valid),
    .REG_pc(frontend_REG_pc),
    .REG_isMissPredict(frontend_REG_isMissPredict),
    .REG_actualTarget(frontend_REG_actualTarget),
    .REG_actualTaken(frontend_REG_actualTaken),
    .REG_fuOpType(frontend_REG_fuOpType),
    .REG_btbType(frontend_REG_btbType),
    .REG_isRVC(frontend_REG_isRVC),
    ._WIRE_0(frontend__WIRE_0),
    .DISPLAY_ENABLE(frontend_DISPLAY_ENABLE),
    ._WIRE_7(frontend__WIRE_7),
    ._WIRE_11(frontend__WIRE_11),
    ._WIRE_1_4(frontend__WIRE_1_4),
    ._WIRE_14(frontend__WIRE_14),
    ._WIRE_2_2(frontend__WIRE_2_2),
    .r_0(frontend_r_0)
  );
  Backend_inorder backend ( // @[src/main/scala/nutcore/NutCore.scala 147:25]
    .clock(backend_clock),
    .reset(backend_reset),
    .io_in_0_ready(backend_io_in_0_ready),
    .io_in_0_valid(backend_io_in_0_valid),
    .io_in_0_bits_cf_instr(backend_io_in_0_bits_cf_instr),
    .io_in_0_bits_cf_pc(backend_io_in_0_bits_cf_pc),
    .io_in_0_bits_cf_pnpc(backend_io_in_0_bits_cf_pnpc),
    .io_in_0_bits_cf_exceptionVec_1(backend_io_in_0_bits_cf_exceptionVec_1),
    .io_in_0_bits_cf_exceptionVec_2(backend_io_in_0_bits_cf_exceptionVec_2),
    .io_in_0_bits_cf_exceptionVec_12(backend_io_in_0_bits_cf_exceptionVec_12),
    .io_in_0_bits_cf_intrVec_0(backend_io_in_0_bits_cf_intrVec_0),
    .io_in_0_bits_cf_intrVec_1(backend_io_in_0_bits_cf_intrVec_1),
    .io_in_0_bits_cf_intrVec_2(backend_io_in_0_bits_cf_intrVec_2),
    .io_in_0_bits_cf_intrVec_3(backend_io_in_0_bits_cf_intrVec_3),
    .io_in_0_bits_cf_intrVec_4(backend_io_in_0_bits_cf_intrVec_4),
    .io_in_0_bits_cf_intrVec_5(backend_io_in_0_bits_cf_intrVec_5),
    .io_in_0_bits_cf_intrVec_6(backend_io_in_0_bits_cf_intrVec_6),
    .io_in_0_bits_cf_intrVec_7(backend_io_in_0_bits_cf_intrVec_7),
    .io_in_0_bits_cf_intrVec_8(backend_io_in_0_bits_cf_intrVec_8),
    .io_in_0_bits_cf_intrVec_9(backend_io_in_0_bits_cf_intrVec_9),
    .io_in_0_bits_cf_intrVec_10(backend_io_in_0_bits_cf_intrVec_10),
    .io_in_0_bits_cf_intrVec_11(backend_io_in_0_bits_cf_intrVec_11),
    .io_in_0_bits_cf_brIdx(backend_io_in_0_bits_cf_brIdx),
    .io_in_0_bits_cf_crossPageIPFFix(backend_io_in_0_bits_cf_crossPageIPFFix),
    .io_in_0_bits_ctrl_src1Type(backend_io_in_0_bits_ctrl_src1Type),
    .io_in_0_bits_ctrl_src2Type(backend_io_in_0_bits_ctrl_src2Type),
    .io_in_0_bits_ctrl_fuType(backend_io_in_0_bits_ctrl_fuType),
    .io_in_0_bits_ctrl_fuOpType(backend_io_in_0_bits_ctrl_fuOpType),
    .io_in_0_bits_ctrl_rfSrc1(backend_io_in_0_bits_ctrl_rfSrc1),
    .io_in_0_bits_ctrl_rfSrc2(backend_io_in_0_bits_ctrl_rfSrc2),
    .io_in_0_bits_ctrl_rfWen(backend_io_in_0_bits_ctrl_rfWen),
    .io_in_0_bits_ctrl_rfDest(backend_io_in_0_bits_ctrl_rfDest),
    .io_in_0_bits_ctrl_isNutCoreTrap(backend_io_in_0_bits_ctrl_isNutCoreTrap),
    .io_in_0_bits_data_imm(backend_io_in_0_bits_data_imm),
    .io_flush(backend_io_flush),
    .io_dmem_req_ready(backend_io_dmem_req_ready),
    .io_dmem_req_valid(backend_io_dmem_req_valid),
    .io_dmem_req_bits_addr(backend_io_dmem_req_bits_addr),
    .io_dmem_req_bits_size(backend_io_dmem_req_bits_size),
    .io_dmem_req_bits_cmd(backend_io_dmem_req_bits_cmd),
    .io_dmem_req_bits_wmask(backend_io_dmem_req_bits_wmask),
    .io_dmem_req_bits_wdata(backend_io_dmem_req_bits_wdata),
    .io_dmem_resp_valid(backend_io_dmem_resp_valid),
    .io_dmem_resp_bits_rdata(backend_io_dmem_resp_bits_rdata),
    .io_memMMU_imem_priviledgeMode(backend_io_memMMU_imem_priviledgeMode),
    .io_memMMU_dmem_priviledgeMode(backend_io_memMMU_dmem_priviledgeMode),
    .io_memMMU_dmem_status_sum(backend_io_memMMU_dmem_status_sum),
    .io_memMMU_dmem_status_mxr(backend_io_memMMU_dmem_status_mxr),
    .io_memMMU_dmem_loadPF(backend_io_memMMU_dmem_loadPF),
    .io_memMMU_dmem_storePF(backend_io_memMMU_dmem_storePF),
    .io_memMMU_dmem_addr(backend_io_memMMU_dmem_addr),
    .io_redirect_target(backend_io_redirect_target),
    .io_redirect_valid(backend_io_redirect_valid),
    .io_extra_meip_0(backend_io_extra_meip_0),
    .REG_valid(backend_REG_valid),
    .REG_pc(backend_REG_pc),
    .REG_isMissPredict(backend_REG_isMissPredict),
    .REG_actualTarget(backend_REG_actualTarget),
    .REG_actualTaken(backend_REG_actualTaken),
    .REG_fuOpType(backend_REG_fuOpType),
    .REG_btbType(backend_REG_btbType),
    .REG_isRVC(backend_REG_isRVC),
    ._WIRE_1(backend__WIRE_1),
    .satp(backend_satp),
    ._WIRE_4(backend__WIRE_4),
    ._WIRE_1_1(backend__WIRE_1_1),
    ._WIRE_7(backend__WIRE_7),
    .io_extra_mtip(backend_io_extra_mtip),
    ._WIRE_11(backend__WIRE_11),
    ._WIRE_1_4(backend__WIRE_1_4),
    ._WIRE_14(backend__WIRE_14),
    ._WIRE_2_2(backend__WIRE_2_2),
    ._WIRE_16(backend__WIRE_16),
    ._WIRE_17(backend__WIRE_17),
    .r_0(backend_r_0),
    .io_extra_msip(backend_io_extra_msip)
  );
  SimpleBusCrossbarNto1 mmioXbar ( // @[src/main/scala/nutcore/NutCore.scala 151:26]
    .clock(mmioXbar_clock),
    .reset(mmioXbar_reset),
    .io_in_0_req_ready(mmioXbar_io_in_0_req_ready),
    .io_in_0_req_valid(mmioXbar_io_in_0_req_valid),
    .io_in_0_req_bits_addr(mmioXbar_io_in_0_req_bits_addr),
    .io_in_0_req_bits_cmd(mmioXbar_io_in_0_req_bits_cmd),
    .io_in_0_req_bits_wmask(mmioXbar_io_in_0_req_bits_wmask),
    .io_in_0_req_bits_wdata(mmioXbar_io_in_0_req_bits_wdata),
    .io_in_0_resp_valid(mmioXbar_io_in_0_resp_valid),
    .io_in_0_resp_bits_cmd(mmioXbar_io_in_0_resp_bits_cmd),
    .io_in_0_resp_bits_rdata(mmioXbar_io_in_0_resp_bits_rdata),
    .io_in_1_req_ready(mmioXbar_io_in_1_req_ready),
    .io_in_1_req_valid(mmioXbar_io_in_1_req_valid),
    .io_in_1_req_bits_addr(mmioXbar_io_in_1_req_bits_addr),
    .io_in_1_req_bits_size(mmioXbar_io_in_1_req_bits_size),
    .io_in_1_req_bits_cmd(mmioXbar_io_in_1_req_bits_cmd),
    .io_in_1_req_bits_wmask(mmioXbar_io_in_1_req_bits_wmask),
    .io_in_1_req_bits_wdata(mmioXbar_io_in_1_req_bits_wdata),
    .io_in_1_resp_valid(mmioXbar_io_in_1_resp_valid),
    .io_in_1_resp_bits_cmd(mmioXbar_io_in_1_resp_bits_cmd),
    .io_in_1_resp_bits_rdata(mmioXbar_io_in_1_resp_bits_rdata),
    .io_out_req_ready(mmioXbar_io_out_req_ready),
    .io_out_req_valid(mmioXbar_io_out_req_valid),
    .io_out_req_bits_addr(mmioXbar_io_out_req_bits_addr),
    .io_out_req_bits_size(mmioXbar_io_out_req_bits_size),
    .io_out_req_bits_cmd(mmioXbar_io_out_req_bits_cmd),
    .io_out_req_bits_wmask(mmioXbar_io_out_req_bits_wmask),
    .io_out_req_bits_wdata(mmioXbar_io_out_req_bits_wdata),
    .io_out_resp_ready(mmioXbar_io_out_resp_ready),
    .io_out_resp_valid(mmioXbar_io_out_resp_valid),
    .io_out_resp_bits_cmd(mmioXbar_io_out_resp_bits_cmd),
    .io_out_resp_bits_rdata(mmioXbar_io_out_resp_bits_rdata)
  );
  SimpleBusCrossbarNto1_1 dmemXbar ( // @[src/main/scala/nutcore/NutCore.scala 152:26]
    .clock(dmemXbar_clock),
    .reset(dmemXbar_reset),
    .io_in_0_req_ready(dmemXbar_io_in_0_req_ready),
    .io_in_0_req_valid(dmemXbar_io_in_0_req_valid),
    .io_in_0_req_bits_addr(dmemXbar_io_in_0_req_bits_addr),
    .io_in_0_req_bits_size(dmemXbar_io_in_0_req_bits_size),
    .io_in_0_req_bits_cmd(dmemXbar_io_in_0_req_bits_cmd),
    .io_in_0_req_bits_wmask(dmemXbar_io_in_0_req_bits_wmask),
    .io_in_0_req_bits_wdata(dmemXbar_io_in_0_req_bits_wdata),
    .io_in_0_resp_valid(dmemXbar_io_in_0_resp_valid),
    .io_in_0_resp_bits_cmd(dmemXbar_io_in_0_resp_bits_cmd),
    .io_in_0_resp_bits_rdata(dmemXbar_io_in_0_resp_bits_rdata),
    .io_in_1_req_ready(dmemXbar_io_in_1_req_ready),
    .io_in_1_req_valid(dmemXbar_io_in_1_req_valid),
    .io_in_1_req_bits_addr(dmemXbar_io_in_1_req_bits_addr),
    .io_in_1_req_bits_cmd(dmemXbar_io_in_1_req_bits_cmd),
    .io_in_1_req_bits_wdata(dmemXbar_io_in_1_req_bits_wdata),
    .io_in_1_resp_valid(dmemXbar_io_in_1_resp_valid),
    .io_in_1_resp_bits_cmd(dmemXbar_io_in_1_resp_bits_cmd),
    .io_in_1_resp_bits_rdata(dmemXbar_io_in_1_resp_bits_rdata),
    .io_in_2_req_ready(dmemXbar_io_in_2_req_ready),
    .io_in_2_req_valid(dmemXbar_io_in_2_req_valid),
    .io_in_2_req_bits_addr(dmemXbar_io_in_2_req_bits_addr),
    .io_in_2_req_bits_cmd(dmemXbar_io_in_2_req_bits_cmd),
    .io_in_2_req_bits_wdata(dmemXbar_io_in_2_req_bits_wdata),
    .io_in_2_resp_valid(dmemXbar_io_in_2_resp_valid),
    .io_in_2_resp_bits_cmd(dmemXbar_io_in_2_resp_bits_cmd),
    .io_in_2_resp_bits_rdata(dmemXbar_io_in_2_resp_bits_rdata),
    .io_in_3_req_ready(dmemXbar_io_in_3_req_ready),
    .io_in_3_req_valid(dmemXbar_io_in_3_req_valid),
    .io_in_3_req_bits_addr(dmemXbar_io_in_3_req_bits_addr),
    .io_in_3_req_bits_size(dmemXbar_io_in_3_req_bits_size),
    .io_in_3_req_bits_cmd(dmemXbar_io_in_3_req_bits_cmd),
    .io_in_3_req_bits_wmask(dmemXbar_io_in_3_req_bits_wmask),
    .io_in_3_req_bits_wdata(dmemXbar_io_in_3_req_bits_wdata),
    .io_in_3_resp_ready(dmemXbar_io_in_3_resp_ready),
    .io_in_3_resp_valid(dmemXbar_io_in_3_resp_valid),
    .io_in_3_resp_bits_cmd(dmemXbar_io_in_3_resp_bits_cmd),
    .io_in_3_resp_bits_rdata(dmemXbar_io_in_3_resp_bits_rdata),
    .io_out_req_ready(dmemXbar_io_out_req_ready),
    .io_out_req_valid(dmemXbar_io_out_req_valid),
    .io_out_req_bits_addr(dmemXbar_io_out_req_bits_addr),
    .io_out_req_bits_size(dmemXbar_io_out_req_bits_size),
    .io_out_req_bits_cmd(dmemXbar_io_out_req_bits_cmd),
    .io_out_req_bits_wmask(dmemXbar_io_out_req_bits_wmask),
    .io_out_req_bits_wdata(dmemXbar_io_out_req_bits_wdata),
    .io_out_resp_ready(dmemXbar_io_out_resp_ready),
    .io_out_resp_valid(dmemXbar_io_out_resp_valid),
    .io_out_resp_bits_cmd(dmemXbar_io_out_resp_bits_cmd),
    .io_out_resp_bits_rdata(dmemXbar_io_out_resp_bits_rdata)
  );
  EmbeddedTLB itlb ( // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 426:13]
    .clock(itlb_clock),
    .reset(itlb_reset),
    .io_in_req_ready(itlb_io_in_req_ready),
    .io_in_req_valid(itlb_io_in_req_valid),
    .io_in_req_bits_addr(itlb_io_in_req_bits_addr),
    .io_in_req_bits_user(itlb_io_in_req_bits_user),
    .io_in_resp_ready(itlb_io_in_resp_ready),
    .io_in_resp_valid(itlb_io_in_resp_valid),
    .io_in_resp_bits_cmd(itlb_io_in_resp_bits_cmd),
    .io_in_resp_bits_rdata(itlb_io_in_resp_bits_rdata),
    .io_in_resp_bits_user(itlb_io_in_resp_bits_user),
    .io_out_req_ready(itlb_io_out_req_ready),
    .io_out_req_valid(itlb_io_out_req_valid),
    .io_out_req_bits_addr(itlb_io_out_req_bits_addr),
    .io_out_req_bits_cmd(itlb_io_out_req_bits_cmd),
    .io_out_req_bits_wdata(itlb_io_out_req_bits_wdata),
    .io_out_req_bits_user(itlb_io_out_req_bits_user),
    .io_out_resp_ready(itlb_io_out_resp_ready),
    .io_out_resp_valid(itlb_io_out_resp_valid),
    .io_out_resp_bits_rdata(itlb_io_out_resp_bits_rdata),
    .io_out_resp_bits_user(itlb_io_out_resp_bits_user),
    .io_mem_req_ready(itlb_io_mem_req_ready),
    .io_mem_req_valid(itlb_io_mem_req_valid),
    .io_mem_req_bits_addr(itlb_io_mem_req_bits_addr),
    .io_mem_req_bits_cmd(itlb_io_mem_req_bits_cmd),
    .io_mem_req_bits_wdata(itlb_io_mem_req_bits_wdata),
    .io_mem_resp_valid(itlb_io_mem_resp_valid),
    .io_mem_resp_bits_cmd(itlb_io_mem_resp_bits_cmd),
    .io_mem_resp_bits_rdata(itlb_io_mem_resp_bits_rdata),
    .io_flush(itlb_io_flush),
    .io_csrMMU_priviledgeMode(itlb_io_csrMMU_priviledgeMode),
    .io_csrMMU_loadPF(itlb_io_csrMMU_loadPF),
    .io_csrMMU_storePF(itlb_io_csrMMU_storePF),
    .io_cacheEmpty(itlb_io_cacheEmpty),
    .io_ipf(itlb_io_ipf),
    .CSRSATP(itlb_CSRSATP),
    .DISPLAY_ENABLE(itlb_DISPLAY_ENABLE),
    .MOUFlushTLB(itlb_MOUFlushTLB)
  );
  Cache io_imem_cache ( // @[src/main/scala/nutcore/mem/Cache.scala 668:35]
    .clock(io_imem_cache_clock),
    .reset(io_imem_cache_reset),
    .io_in_req_ready(io_imem_cache_io_in_req_ready),
    .io_in_req_valid(io_imem_cache_io_in_req_valid),
    .io_in_req_bits_addr(io_imem_cache_io_in_req_bits_addr),
    .io_in_req_bits_user(io_imem_cache_io_in_req_bits_user),
    .io_in_resp_ready(io_imem_cache_io_in_resp_ready),
    .io_in_resp_valid(io_imem_cache_io_in_resp_valid),
    .io_in_resp_bits_rdata(io_imem_cache_io_in_resp_bits_rdata),
    .io_in_resp_bits_user(io_imem_cache_io_in_resp_bits_user),
    .io_flush(io_imem_cache_io_flush),
    .io_out_mem_req_ready(io_imem_cache_io_out_mem_req_ready),
    .io_out_mem_req_valid(io_imem_cache_io_out_mem_req_valid),
    .io_out_mem_req_bits_addr(io_imem_cache_io_out_mem_req_bits_addr),
    .io_out_mem_req_bits_cmd(io_imem_cache_io_out_mem_req_bits_cmd),
    .io_out_mem_req_bits_wdata(io_imem_cache_io_out_mem_req_bits_wdata),
    .io_out_mem_resp_valid(io_imem_cache_io_out_mem_resp_valid),
    .io_out_mem_resp_bits_cmd(io_imem_cache_io_out_mem_resp_bits_cmd),
    .io_out_mem_resp_bits_rdata(io_imem_cache_io_out_mem_resp_bits_rdata),
    .io_mmio_req_ready(io_imem_cache_io_mmio_req_ready),
    .io_mmio_req_valid(io_imem_cache_io_mmio_req_valid),
    .io_mmio_req_bits_addr(io_imem_cache_io_mmio_req_bits_addr),
    .io_mmio_resp_valid(io_imem_cache_io_mmio_resp_valid),
    .io_mmio_resp_bits_rdata(io_imem_cache_io_mmio_resp_bits_rdata),
    .io_empty(io_imem_cache_io_empty),
    .DISPLAY_ENABLE(io_imem_cache_DISPLAY_ENABLE),
    .MOUFlushICache(io_imem_cache_MOUFlushICache)
  );
  EmbeddedTLB_1 dtlb ( // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 426:13]
    .clock(dtlb_clock),
    .reset(dtlb_reset),
    .io_in_req_ready(dtlb_io_in_req_ready),
    .io_in_req_valid(dtlb_io_in_req_valid),
    .io_in_req_bits_addr(dtlb_io_in_req_bits_addr),
    .io_in_req_bits_size(dtlb_io_in_req_bits_size),
    .io_in_req_bits_cmd(dtlb_io_in_req_bits_cmd),
    .io_in_req_bits_wmask(dtlb_io_in_req_bits_wmask),
    .io_in_req_bits_wdata(dtlb_io_in_req_bits_wdata),
    .io_in_resp_valid(dtlb_io_in_resp_valid),
    .io_in_resp_bits_cmd(dtlb_io_in_resp_bits_cmd),
    .io_in_resp_bits_rdata(dtlb_io_in_resp_bits_rdata),
    .io_out_req_ready(dtlb_io_out_req_ready),
    .io_out_req_valid(dtlb_io_out_req_valid),
    .io_out_req_bits_addr(dtlb_io_out_req_bits_addr),
    .io_out_req_bits_size(dtlb_io_out_req_bits_size),
    .io_out_req_bits_cmd(dtlb_io_out_req_bits_cmd),
    .io_out_req_bits_wmask(dtlb_io_out_req_bits_wmask),
    .io_out_req_bits_wdata(dtlb_io_out_req_bits_wdata),
    .io_out_resp_ready(dtlb_io_out_resp_ready),
    .io_out_resp_valid(dtlb_io_out_resp_valid),
    .io_out_resp_bits_cmd(dtlb_io_out_resp_bits_cmd),
    .io_out_resp_bits_rdata(dtlb_io_out_resp_bits_rdata),
    .io_mem_req_ready(dtlb_io_mem_req_ready),
    .io_mem_req_valid(dtlb_io_mem_req_valid),
    .io_mem_req_bits_addr(dtlb_io_mem_req_bits_addr),
    .io_mem_req_bits_cmd(dtlb_io_mem_req_bits_cmd),
    .io_mem_req_bits_wdata(dtlb_io_mem_req_bits_wdata),
    .io_mem_resp_valid(dtlb_io_mem_resp_valid),
    .io_mem_resp_bits_cmd(dtlb_io_mem_resp_bits_cmd),
    .io_mem_resp_bits_rdata(dtlb_io_mem_resp_bits_rdata),
    .io_csrMMU_priviledgeMode(dtlb_io_csrMMU_priviledgeMode),
    .io_csrMMU_status_sum(dtlb_io_csrMMU_status_sum),
    .io_csrMMU_status_mxr(dtlb_io_csrMMU_status_mxr),
    .io_csrMMU_loadPF(dtlb_io_csrMMU_loadPF),
    .io_csrMMU_storePF(dtlb_io_csrMMU_storePF),
    .io_csrMMU_addr(dtlb_io_csrMMU_addr),
    .io_cacheEmpty(dtlb_io_cacheEmpty),
    .io_ipf(dtlb_io_ipf),
    ._WIRE_4(dtlb__WIRE_4),
    .CSRSATP(dtlb_CSRSATP),
    .DISPLAY_ENABLE(dtlb_DISPLAY_ENABLE),
    ._WIRE_1_1(dtlb__WIRE_1_1),
    .MOUFlushTLB(dtlb_MOUFlushTLB),
    ._WIRE_2_3(dtlb__WIRE_2_3),
    ._WIRE_16(dtlb__WIRE_16)
  );
  Cache_1 io_dmem_cache ( // @[src/main/scala/nutcore/mem/Cache.scala 668:35]
    .clock(io_dmem_cache_clock),
    .reset(io_dmem_cache_reset),
    .io_in_req_ready(io_dmem_cache_io_in_req_ready),
    .io_in_req_valid(io_dmem_cache_io_in_req_valid),
    .io_in_req_bits_addr(io_dmem_cache_io_in_req_bits_addr),
    .io_in_req_bits_size(io_dmem_cache_io_in_req_bits_size),
    .io_in_req_bits_cmd(io_dmem_cache_io_in_req_bits_cmd),
    .io_in_req_bits_wmask(io_dmem_cache_io_in_req_bits_wmask),
    .io_in_req_bits_wdata(io_dmem_cache_io_in_req_bits_wdata),
    .io_in_resp_ready(io_dmem_cache_io_in_resp_ready),
    .io_in_resp_valid(io_dmem_cache_io_in_resp_valid),
    .io_in_resp_bits_cmd(io_dmem_cache_io_in_resp_bits_cmd),
    .io_in_resp_bits_rdata(io_dmem_cache_io_in_resp_bits_rdata),
    .io_out_mem_req_ready(io_dmem_cache_io_out_mem_req_ready),
    .io_out_mem_req_valid(io_dmem_cache_io_out_mem_req_valid),
    .io_out_mem_req_bits_addr(io_dmem_cache_io_out_mem_req_bits_addr),
    .io_out_mem_req_bits_cmd(io_dmem_cache_io_out_mem_req_bits_cmd),
    .io_out_mem_req_bits_wdata(io_dmem_cache_io_out_mem_req_bits_wdata),
    .io_out_mem_resp_valid(io_dmem_cache_io_out_mem_resp_valid),
    .io_out_mem_resp_bits_cmd(io_dmem_cache_io_out_mem_resp_bits_cmd),
    .io_out_mem_resp_bits_rdata(io_dmem_cache_io_out_mem_resp_bits_rdata),
    .io_out_coh_req_ready(io_dmem_cache_io_out_coh_req_ready),
    .io_out_coh_req_valid(io_dmem_cache_io_out_coh_req_valid),
    .io_out_coh_req_bits_addr(io_dmem_cache_io_out_coh_req_bits_addr),
    .io_out_coh_req_bits_wdata(io_dmem_cache_io_out_coh_req_bits_wdata),
    .io_out_coh_resp_valid(io_dmem_cache_io_out_coh_resp_valid),
    .io_out_coh_resp_bits_cmd(io_dmem_cache_io_out_coh_resp_bits_cmd),
    .io_out_coh_resp_bits_rdata(io_dmem_cache_io_out_coh_resp_bits_rdata),
    .io_mmio_req_ready(io_dmem_cache_io_mmio_req_ready),
    .io_mmio_req_valid(io_dmem_cache_io_mmio_req_valid),
    .io_mmio_req_bits_addr(io_dmem_cache_io_mmio_req_bits_addr),
    .io_mmio_req_bits_size(io_dmem_cache_io_mmio_req_bits_size),
    .io_mmio_req_bits_cmd(io_dmem_cache_io_mmio_req_bits_cmd),
    .io_mmio_req_bits_wmask(io_dmem_cache_io_mmio_req_bits_wmask),
    .io_mmio_req_bits_wdata(io_dmem_cache_io_mmio_req_bits_wdata),
    .io_mmio_resp_valid(io_dmem_cache_io_mmio_resp_valid),
    .io_mmio_resp_bits_rdata(io_dmem_cache_io_mmio_resp_bits_rdata),
    .io_empty(io_dmem_cache_io_empty),
    .DISPLAY_ENABLE(io_dmem_cache_DISPLAY_ENABLE),
    ._WIRE_17(io_dmem_cache__WIRE_17)
  );
  assign io_imem_mem_req_valid = io_imem_cache_io_out_mem_req_valid; // @[src/main/scala/nutcore/NutCore.scala 156:13]
  assign io_imem_mem_req_bits_addr = io_imem_cache_io_out_mem_req_bits_addr; // @[src/main/scala/nutcore/NutCore.scala 156:13]
  assign io_imem_mem_req_bits_cmd = io_imem_cache_io_out_mem_req_bits_cmd; // @[src/main/scala/nutcore/NutCore.scala 156:13]
  assign io_imem_mem_req_bits_wdata = io_imem_cache_io_out_mem_req_bits_wdata; // @[src/main/scala/nutcore/NutCore.scala 156:13]
  assign io_dmem_mem_req_valid = io_dmem_cache_io_out_mem_req_valid; // @[src/main/scala/nutcore/NutCore.scala 161:13]
  assign io_dmem_mem_req_bits_addr = io_dmem_cache_io_out_mem_req_bits_addr; // @[src/main/scala/nutcore/NutCore.scala 161:13]
  assign io_dmem_mem_req_bits_cmd = io_dmem_cache_io_out_mem_req_bits_cmd; // @[src/main/scala/nutcore/NutCore.scala 161:13]
  assign io_dmem_mem_req_bits_wdata = io_dmem_cache_io_out_mem_req_bits_wdata; // @[src/main/scala/nutcore/NutCore.scala 161:13]
  assign io_dmem_coh_req_ready = io_dmem_cache_io_out_coh_req_ready; // @[src/main/scala/nutcore/NutCore.scala 161:13]
  assign io_dmem_coh_resp_valid = io_dmem_cache_io_out_coh_resp_valid; // @[src/main/scala/nutcore/NutCore.scala 161:13]
  assign io_dmem_coh_resp_bits_cmd = io_dmem_cache_io_out_coh_resp_bits_cmd; // @[src/main/scala/nutcore/NutCore.scala 161:13]
  assign io_dmem_coh_resp_bits_rdata = io_dmem_cache_io_out_coh_resp_bits_rdata; // @[src/main/scala/nutcore/NutCore.scala 161:13]
  assign io_mmio_req_valid = mmioXbar_io_out_req_valid; // @[src/main/scala/nutcore/NutCore.scala 170:13]
  assign io_mmio_req_bits_addr = mmioXbar_io_out_req_bits_addr; // @[src/main/scala/nutcore/NutCore.scala 170:13]
  assign io_mmio_req_bits_size = mmioXbar_io_out_req_bits_size; // @[src/main/scala/nutcore/NutCore.scala 170:13]
  assign io_mmio_req_bits_cmd = mmioXbar_io_out_req_bits_cmd; // @[src/main/scala/nutcore/NutCore.scala 170:13]
  assign io_mmio_req_bits_wmask = mmioXbar_io_out_req_bits_wmask; // @[src/main/scala/nutcore/NutCore.scala 170:13]
  assign io_mmio_req_bits_wdata = mmioXbar_io_out_req_bits_wdata; // @[src/main/scala/nutcore/NutCore.scala 170:13]
  assign io_frontend_req_ready = dmemXbar_io_in_3_req_ready; // @[src/main/scala/nutcore/NutCore.scala 168:23]
  assign io_frontend_resp_valid = dmemXbar_io_in_3_resp_valid; // @[src/main/scala/nutcore/NutCore.scala 168:23]
  assign io_frontend_resp_bits_cmd = dmemXbar_io_in_3_resp_bits_cmd; // @[src/main/scala/nutcore/NutCore.scala 168:23]
  assign io_frontend_resp_bits_rdata = dmemXbar_io_in_3_resp_bits_rdata; // @[src/main/scala/nutcore/NutCore.scala 168:23]
  assign _WIRE_0 = frontend__WIRE_0;
  assign frontend_clock = clock;
  assign frontend_reset = reset;
  assign frontend_io_imem_req_ready = itlb_io_in_req_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 430:15]
  assign frontend_io_imem_resp_valid = itlb_io_in_resp_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 430:15]
  assign frontend_io_imem_resp_bits_rdata = itlb_io_in_resp_bits_rdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 430:15]
  assign frontend_io_imem_resp_bits_user = itlb_io_in_resp_bits_user; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 430:15]
  assign frontend_io_out_0_ready = ringBufferAllowin | ~frontend_io_out_0_valid; // @[src/main/scala/utils/PipelineVector.scala 50:36]
  assign frontend_io_redirect_target = backend_io_redirect_target; // @[src/main/scala/nutcore/NutCore.scala 164:26]
  assign frontend_io_redirect_valid = backend_io_redirect_valid; // @[src/main/scala/nutcore/NutCore.scala 164:26]
  assign frontend_io_ipf = itlb_io_ipf; // @[src/main/scala/nutcore/NutCore.scala 155:21]
  assign frontend_REG_valid = backend_REG_valid;
  assign frontend_REG_pc = backend_REG_pc;
  assign frontend_REG_isMissPredict = backend_REG_isMissPredict;
  assign frontend_REG_actualTarget = backend_REG_actualTarget;
  assign frontend_REG_actualTaken = backend_REG_actualTaken;
  assign frontend_REG_fuOpType = backend_REG_fuOpType;
  assign frontend_REG_btbType = backend_REG_btbType;
  assign frontend_REG_isRVC = backend_REG_isRVC;
  assign frontend_DISPLAY_ENABLE = DISPLAY_ENABLE;
  assign frontend__WIRE_11 = backend__WIRE_11;
  assign frontend__WIRE_1_4 = backend__WIRE_1_4;
  assign frontend__WIRE_14 = backend__WIRE_14;
  assign frontend__WIRE_2_2 = dtlb__WIRE_2_3;
  assign backend_clock = clock;
  assign backend_reset = reset;
  assign backend_io_in_0_valid = ringBufferHead != ringBufferTail; // @[src/main/scala/utils/PipelineVector.scala 56:34]
  assign backend_io_in_0_bits_cf_instr = 2'h3 == ringBufferTail ? dataBuffer_3_cf_instr : _GEN_1319; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  assign backend_io_in_0_bits_cf_pc = 2'h3 == ringBufferTail ? dataBuffer_3_cf_pc : _GEN_1315; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  assign backend_io_in_0_bits_cf_pnpc = 2'h3 == ringBufferTail ? dataBuffer_3_cf_pnpc : _GEN_1311; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  assign backend_io_in_0_bits_cf_exceptionVec_1 = 2'h3 == ringBufferTail ? dataBuffer_3_cf_exceptionVec_1 : _GEN_1239; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  assign backend_io_in_0_bits_cf_exceptionVec_2 = 2'h3 == ringBufferTail ? dataBuffer_3_cf_exceptionVec_2 : _GEN_1243; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  assign backend_io_in_0_bits_cf_exceptionVec_12 = 2'h3 == ringBufferTail ? dataBuffer_3_cf_exceptionVec_12 : _GEN_1283; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  assign backend_io_in_0_bits_cf_intrVec_0 = 2'h3 == ringBufferTail ? dataBuffer_3_cf_intrVec_0 : _GEN_1187; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  assign backend_io_in_0_bits_cf_intrVec_1 = 2'h3 == ringBufferTail ? dataBuffer_3_cf_intrVec_1 : _GEN_1191; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  assign backend_io_in_0_bits_cf_intrVec_2 = 2'h3 == ringBufferTail ? dataBuffer_3_cf_intrVec_2 : _GEN_1195; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  assign backend_io_in_0_bits_cf_intrVec_3 = 2'h3 == ringBufferTail ? dataBuffer_3_cf_intrVec_3 : _GEN_1199; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  assign backend_io_in_0_bits_cf_intrVec_4 = 2'h3 == ringBufferTail ? dataBuffer_3_cf_intrVec_4 : _GEN_1203; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  assign backend_io_in_0_bits_cf_intrVec_5 = 2'h3 == ringBufferTail ? dataBuffer_3_cf_intrVec_5 : _GEN_1207; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  assign backend_io_in_0_bits_cf_intrVec_6 = 2'h3 == ringBufferTail ? dataBuffer_3_cf_intrVec_6 : _GEN_1211; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  assign backend_io_in_0_bits_cf_intrVec_7 = 2'h3 == ringBufferTail ? dataBuffer_3_cf_intrVec_7 : _GEN_1215; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  assign backend_io_in_0_bits_cf_intrVec_8 = 2'h3 == ringBufferTail ? dataBuffer_3_cf_intrVec_8 : _GEN_1219; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  assign backend_io_in_0_bits_cf_intrVec_9 = 2'h3 == ringBufferTail ? dataBuffer_3_cf_intrVec_9 : _GEN_1223; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  assign backend_io_in_0_bits_cf_intrVec_10 = 2'h3 == ringBufferTail ? dataBuffer_3_cf_intrVec_10 : _GEN_1227; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  assign backend_io_in_0_bits_cf_intrVec_11 = 2'h3 == ringBufferTail ? dataBuffer_3_cf_intrVec_11 : _GEN_1231; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  assign backend_io_in_0_bits_cf_brIdx = 2'h3 == ringBufferTail ? dataBuffer_3_cf_brIdx : _GEN_1183; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  assign backend_io_in_0_bits_cf_crossPageIPFFix = 2'h3 == ringBufferTail ? dataBuffer_3_cf_crossPageIPFFix : _GEN_1175; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  assign backend_io_in_0_bits_ctrl_src1Type = 2'h3 == ringBufferTail ? dataBuffer_3_ctrl_src1Type : _GEN_1163; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  assign backend_io_in_0_bits_ctrl_src2Type = 2'h3 == ringBufferTail ? dataBuffer_3_ctrl_src2Type : _GEN_1159; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  assign backend_io_in_0_bits_ctrl_fuType = 2'h3 == ringBufferTail ? dataBuffer_3_ctrl_fuType : _GEN_1155; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  assign backend_io_in_0_bits_ctrl_fuOpType = 2'h3 == ringBufferTail ? dataBuffer_3_ctrl_fuOpType : _GEN_1151; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  assign backend_io_in_0_bits_ctrl_rfSrc1 = 2'h3 == ringBufferTail ? dataBuffer_3_ctrl_rfSrc1 : _GEN_1147; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  assign backend_io_in_0_bits_ctrl_rfSrc2 = 2'h3 == ringBufferTail ? dataBuffer_3_ctrl_rfSrc2 : _GEN_1143; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  assign backend_io_in_0_bits_ctrl_rfWen = 2'h3 == ringBufferTail ? dataBuffer_3_ctrl_rfWen : _GEN_1139; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  assign backend_io_in_0_bits_ctrl_rfDest = 2'h3 == ringBufferTail ? dataBuffer_3_ctrl_rfDest : _GEN_1135; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  assign backend_io_in_0_bits_ctrl_isNutCoreTrap = 2'h3 == ringBufferTail ? dataBuffer_3_ctrl_isNutCoreTrap : _GEN_1131; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  assign backend_io_in_0_bits_data_imm = 2'h3 == ringBufferTail ? dataBuffer_3_data_imm : _GEN_1103; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  assign backend_io_flush = frontend_io_flushVec[3:2]; // @[src/main/scala/nutcore/NutCore.scala 165:45]
  assign backend_io_dmem_req_ready = dtlb_io_in_req_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 430:15]
  assign backend_io_dmem_resp_valid = dtlb_io_in_resp_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 430:15]
  assign backend_io_dmem_resp_bits_rdata = dtlb_io_in_resp_bits_rdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 430:15]
  assign backend_io_memMMU_dmem_loadPF = dtlb_io_csrMMU_loadPF; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 433:19]
  assign backend_io_memMMU_dmem_storePF = dtlb_io_csrMMU_storePF; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 433:19]
  assign backend_io_memMMU_dmem_addr = dtlb_io_csrMMU_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 433:19]
  assign backend_io_extra_meip_0 = io_extra_meip_0;
  assign backend__WIRE_4 = DISPLAY_ENABLE;
  assign backend__WIRE_1_1 = dtlb__WIRE_1_1;
  assign backend__WIRE_7 = frontend__WIRE_7;
  assign backend_io_extra_mtip = io_extra_mtip;
  assign backend__WIRE_2_2 = dtlb__WIRE_2_3;
  assign backend__WIRE_16 = dtlb__WIRE_16;
  assign backend__WIRE_17 = io_dmem_cache__WIRE_17;
  assign backend_r_0 = frontend_r_0;
  assign backend_io_extra_msip = io_extra_msip;
  assign mmioXbar_clock = clock;
  assign mmioXbar_reset = reset;
  assign mmioXbar_io_in_0_req_valid = io_imem_cache_io_mmio_req_valid; // @[src/main/scala/nutcore/mem/Cache.scala 675:13]
  assign mmioXbar_io_in_0_req_bits_addr = io_imem_cache_io_mmio_req_bits_addr; // @[src/main/scala/nutcore/mem/Cache.scala 675:13]
  assign mmioXbar_io_in_0_req_bits_cmd = 4'h0; // @[src/main/scala/nutcore/mem/Cache.scala 675:13]
  assign mmioXbar_io_in_0_req_bits_wmask = 8'h0; // @[src/main/scala/nutcore/mem/Cache.scala 675:13]
  assign mmioXbar_io_in_0_req_bits_wdata = 64'h0; // @[src/main/scala/nutcore/mem/Cache.scala 675:13]
  assign mmioXbar_io_in_1_req_valid = io_dmem_cache_io_mmio_req_valid; // @[src/main/scala/nutcore/mem/Cache.scala 675:13]
  assign mmioXbar_io_in_1_req_bits_addr = io_dmem_cache_io_mmio_req_bits_addr; // @[src/main/scala/nutcore/mem/Cache.scala 675:13]
  assign mmioXbar_io_in_1_req_bits_size = io_dmem_cache_io_mmio_req_bits_size; // @[src/main/scala/nutcore/mem/Cache.scala 675:13]
  assign mmioXbar_io_in_1_req_bits_cmd = io_dmem_cache_io_mmio_req_bits_cmd; // @[src/main/scala/nutcore/mem/Cache.scala 675:13]
  assign mmioXbar_io_in_1_req_bits_wmask = io_dmem_cache_io_mmio_req_bits_wmask; // @[src/main/scala/nutcore/mem/Cache.scala 675:13]
  assign mmioXbar_io_in_1_req_bits_wdata = io_dmem_cache_io_mmio_req_bits_wdata; // @[src/main/scala/nutcore/mem/Cache.scala 675:13]
  assign mmioXbar_io_out_req_ready = io_mmio_req_ready; // @[src/main/scala/nutcore/NutCore.scala 170:13]
  assign mmioXbar_io_out_resp_valid = io_mmio_resp_valid; // @[src/main/scala/nutcore/NutCore.scala 170:13]
  assign mmioXbar_io_out_resp_bits_cmd = io_mmio_resp_bits_cmd; // @[src/main/scala/nutcore/NutCore.scala 170:13]
  assign mmioXbar_io_out_resp_bits_rdata = io_mmio_resp_bits_rdata; // @[src/main/scala/nutcore/NutCore.scala 170:13]
  assign dmemXbar_clock = clock;
  assign dmemXbar_reset = reset;
  assign dmemXbar_io_in_0_req_valid = dtlb_io_out_req_valid; // @[src/main/scala/nutcore/NutCore.scala 160:23]
  assign dmemXbar_io_in_0_req_bits_addr = dtlb_io_out_req_bits_addr; // @[src/main/scala/nutcore/NutCore.scala 160:23]
  assign dmemXbar_io_in_0_req_bits_size = dtlb_io_out_req_bits_size; // @[src/main/scala/nutcore/NutCore.scala 160:23]
  assign dmemXbar_io_in_0_req_bits_cmd = dtlb_io_out_req_bits_cmd; // @[src/main/scala/nutcore/NutCore.scala 160:23]
  assign dmemXbar_io_in_0_req_bits_wmask = dtlb_io_out_req_bits_wmask; // @[src/main/scala/nutcore/NutCore.scala 160:23]
  assign dmemXbar_io_in_0_req_bits_wdata = dtlb_io_out_req_bits_wdata; // @[src/main/scala/nutcore/NutCore.scala 160:23]
  assign dmemXbar_io_in_1_req_valid = itlb_io_mem_req_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 431:16]
  assign dmemXbar_io_in_1_req_bits_addr = itlb_io_mem_req_bits_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 431:16]
  assign dmemXbar_io_in_1_req_bits_cmd = itlb_io_mem_req_bits_cmd; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 431:16]
  assign dmemXbar_io_in_1_req_bits_wdata = itlb_io_mem_req_bits_wdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 431:16]
  assign dmemXbar_io_in_2_req_valid = dtlb_io_mem_req_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 431:16]
  assign dmemXbar_io_in_2_req_bits_addr = dtlb_io_mem_req_bits_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 431:16]
  assign dmemXbar_io_in_2_req_bits_cmd = dtlb_io_mem_req_bits_cmd; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 431:16]
  assign dmemXbar_io_in_2_req_bits_wdata = dtlb_io_mem_req_bits_wdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 431:16]
  assign dmemXbar_io_in_3_req_valid = io_frontend_req_valid; // @[src/main/scala/nutcore/NutCore.scala 168:23]
  assign dmemXbar_io_in_3_req_bits_addr = io_frontend_req_bits_addr; // @[src/main/scala/nutcore/NutCore.scala 168:23]
  assign dmemXbar_io_in_3_req_bits_size = io_frontend_req_bits_size; // @[src/main/scala/nutcore/NutCore.scala 168:23]
  assign dmemXbar_io_in_3_req_bits_cmd = io_frontend_req_bits_cmd; // @[src/main/scala/nutcore/NutCore.scala 168:23]
  assign dmemXbar_io_in_3_req_bits_wmask = io_frontend_req_bits_wmask; // @[src/main/scala/nutcore/NutCore.scala 168:23]
  assign dmemXbar_io_in_3_req_bits_wdata = io_frontend_req_bits_wdata; // @[src/main/scala/nutcore/NutCore.scala 168:23]
  assign dmemXbar_io_in_3_resp_ready = io_frontend_resp_ready; // @[src/main/scala/nutcore/NutCore.scala 168:23]
  assign dmemXbar_io_out_req_ready = io_dmem_cache_io_in_req_ready; // @[src/main/scala/nutcore/mem/Cache.scala 674:17]
  assign dmemXbar_io_out_resp_valid = io_dmem_cache_io_in_resp_valid; // @[src/main/scala/nutcore/mem/Cache.scala 674:17]
  assign dmemXbar_io_out_resp_bits_cmd = io_dmem_cache_io_in_resp_bits_cmd; // @[src/main/scala/nutcore/mem/Cache.scala 674:17]
  assign dmemXbar_io_out_resp_bits_rdata = io_dmem_cache_io_in_resp_bits_rdata; // @[src/main/scala/nutcore/mem/Cache.scala 674:17]
  assign itlb_clock = clock;
  assign itlb_reset = reset;
  assign itlb_io_in_req_valid = frontend_io_imem_req_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 430:15]
  assign itlb_io_in_req_bits_addr = frontend_io_imem_req_bits_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 430:15]
  assign itlb_io_in_req_bits_user = frontend_io_imem_req_bits_user; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 430:15]
  assign itlb_io_in_resp_ready = frontend_io_imem_resp_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 430:15]
  assign itlb_io_out_req_ready = io_imem_cache_io_in_req_ready; // @[src/main/scala/nutcore/mem/Cache.scala 674:17]
  assign itlb_io_out_resp_valid = io_imem_cache_io_in_resp_valid; // @[src/main/scala/nutcore/mem/Cache.scala 674:17]
  assign itlb_io_out_resp_bits_rdata = io_imem_cache_io_in_resp_bits_rdata; // @[src/main/scala/nutcore/mem/Cache.scala 674:17]
  assign itlb_io_out_resp_bits_user = io_imem_cache_io_in_resp_bits_user; // @[src/main/scala/nutcore/mem/Cache.scala 674:17]
  assign itlb_io_mem_req_ready = dmemXbar_io_in_1_req_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 431:16]
  assign itlb_io_mem_resp_valid = dmemXbar_io_in_1_resp_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 431:16]
  assign itlb_io_mem_resp_bits_cmd = dmemXbar_io_in_1_resp_bits_cmd; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 431:16]
  assign itlb_io_mem_resp_bits_rdata = dmemXbar_io_in_1_resp_bits_rdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 431:16]
  assign itlb_io_flush = frontend_io_flushVec[0]; // @[src/main/scala/nutcore/NutCore.scala 154:104]
  assign itlb_io_csrMMU_priviledgeMode = backend_io_memMMU_imem_priviledgeMode; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 433:19]
  assign itlb_io_cacheEmpty = io_imem_cache_io_empty; // @[src/main/scala/nutcore/mem/Cache.scala 676:11]
  assign itlb_CSRSATP = backend_satp;
  assign itlb_DISPLAY_ENABLE = DISPLAY_ENABLE;
  assign itlb_MOUFlushTLB = backend__WIRE_1_4;
  assign io_imem_cache_clock = clock;
  assign io_imem_cache_reset = reset;
  assign io_imem_cache_io_in_req_valid = itlb_io_out_req_valid; // @[src/main/scala/nutcore/mem/Cache.scala 674:17]
  assign io_imem_cache_io_in_req_bits_addr = itlb_io_out_req_bits_addr; // @[src/main/scala/nutcore/mem/Cache.scala 674:17]
  assign io_imem_cache_io_in_req_bits_user = itlb_io_out_req_bits_user; // @[src/main/scala/nutcore/mem/Cache.scala 674:17]
  assign io_imem_cache_io_in_resp_ready = itlb_io_out_resp_ready; // @[src/main/scala/nutcore/mem/Cache.scala 674:17]
  assign io_imem_cache_io_flush = frontend_io_flushVec[0] ? 2'h3 : 2'h0; // @[src/main/scala/nutcore/NutCore.scala 156:83]
  assign io_imem_cache_io_out_mem_req_ready = io_imem_mem_req_ready; // @[src/main/scala/nutcore/NutCore.scala 156:13]
  assign io_imem_cache_io_out_mem_resp_valid = io_imem_mem_resp_valid; // @[src/main/scala/nutcore/NutCore.scala 156:13]
  assign io_imem_cache_io_out_mem_resp_bits_cmd = io_imem_mem_resp_bits_cmd; // @[src/main/scala/nutcore/NutCore.scala 156:13]
  assign io_imem_cache_io_out_mem_resp_bits_rdata = io_imem_mem_resp_bits_rdata; // @[src/main/scala/nutcore/NutCore.scala 156:13]
  assign io_imem_cache_io_mmio_req_ready = mmioXbar_io_in_0_req_ready; // @[src/main/scala/nutcore/mem/Cache.scala 675:13]
  assign io_imem_cache_io_mmio_resp_valid = mmioXbar_io_in_0_resp_valid; // @[src/main/scala/nutcore/mem/Cache.scala 675:13]
  assign io_imem_cache_io_mmio_resp_bits_rdata = mmioXbar_io_in_0_resp_bits_rdata; // @[src/main/scala/nutcore/mem/Cache.scala 675:13]
  assign io_imem_cache_DISPLAY_ENABLE = DISPLAY_ENABLE;
  assign io_imem_cache_MOUFlushICache = backend__WIRE_11;
  assign dtlb_clock = clock;
  assign dtlb_reset = reset;
  assign dtlb_io_in_req_valid = backend_io_dmem_req_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 430:15]
  assign dtlb_io_in_req_bits_addr = backend_io_dmem_req_bits_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 430:15]
  assign dtlb_io_in_req_bits_size = backend_io_dmem_req_bits_size; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 430:15]
  assign dtlb_io_in_req_bits_cmd = backend_io_dmem_req_bits_cmd; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 430:15]
  assign dtlb_io_in_req_bits_wmask = backend_io_dmem_req_bits_wmask; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 430:15]
  assign dtlb_io_in_req_bits_wdata = backend_io_dmem_req_bits_wdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 430:15]
  assign dtlb_io_out_req_ready = dmemXbar_io_in_0_req_ready; // @[src/main/scala/nutcore/NutCore.scala 160:23]
  assign dtlb_io_out_resp_valid = dmemXbar_io_in_0_resp_valid; // @[src/main/scala/nutcore/NutCore.scala 160:23]
  assign dtlb_io_out_resp_bits_cmd = dmemXbar_io_in_0_resp_bits_cmd; // @[src/main/scala/nutcore/NutCore.scala 160:23]
  assign dtlb_io_out_resp_bits_rdata = dmemXbar_io_in_0_resp_bits_rdata; // @[src/main/scala/nutcore/NutCore.scala 160:23]
  assign dtlb_io_mem_req_ready = dmemXbar_io_in_2_req_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 431:16]
  assign dtlb_io_mem_resp_valid = dmemXbar_io_in_2_resp_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 431:16]
  assign dtlb_io_mem_resp_bits_cmd = dmemXbar_io_in_2_resp_bits_cmd; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 431:16]
  assign dtlb_io_mem_resp_bits_rdata = dmemXbar_io_in_2_resp_bits_rdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 431:16]
  assign dtlb_io_csrMMU_priviledgeMode = backend_io_memMMU_dmem_priviledgeMode; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 433:19]
  assign dtlb_io_csrMMU_status_sum = backend_io_memMMU_dmem_status_sum; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 433:19]
  assign dtlb_io_csrMMU_status_mxr = backend_io_memMMU_dmem_status_mxr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 433:19]
  assign dtlb_io_cacheEmpty = io_dmem_cache_io_empty; // @[src/main/scala/nutcore/mem/Cache.scala 676:11]
  assign dtlb__WIRE_4 = backend__WIRE_1;
  assign dtlb_CSRSATP = backend_satp;
  assign dtlb_DISPLAY_ENABLE = DISPLAY_ENABLE;
  assign dtlb_MOUFlushTLB = backend__WIRE_1_4;
  assign io_dmem_cache_clock = clock;
  assign io_dmem_cache_reset = reset;
  assign io_dmem_cache_io_in_req_valid = dmemXbar_io_out_req_valid; // @[src/main/scala/nutcore/mem/Cache.scala 674:17]
  assign io_dmem_cache_io_in_req_bits_addr = dmemXbar_io_out_req_bits_addr; // @[src/main/scala/nutcore/mem/Cache.scala 674:17]
  assign io_dmem_cache_io_in_req_bits_size = dmemXbar_io_out_req_bits_size; // @[src/main/scala/nutcore/mem/Cache.scala 674:17]
  assign io_dmem_cache_io_in_req_bits_cmd = dmemXbar_io_out_req_bits_cmd; // @[src/main/scala/nutcore/mem/Cache.scala 674:17]
  assign io_dmem_cache_io_in_req_bits_wmask = dmemXbar_io_out_req_bits_wmask; // @[src/main/scala/nutcore/mem/Cache.scala 674:17]
  assign io_dmem_cache_io_in_req_bits_wdata = dmemXbar_io_out_req_bits_wdata; // @[src/main/scala/nutcore/mem/Cache.scala 674:17]
  assign io_dmem_cache_io_in_resp_ready = dmemXbar_io_out_resp_ready; // @[src/main/scala/nutcore/mem/Cache.scala 674:17]
  assign io_dmem_cache_io_out_mem_req_ready = io_dmem_mem_req_ready; // @[src/main/scala/nutcore/NutCore.scala 161:13]
  assign io_dmem_cache_io_out_mem_resp_valid = io_dmem_mem_resp_valid; // @[src/main/scala/nutcore/NutCore.scala 161:13]
  assign io_dmem_cache_io_out_mem_resp_bits_cmd = io_dmem_mem_resp_bits_cmd; // @[src/main/scala/nutcore/NutCore.scala 161:13]
  assign io_dmem_cache_io_out_mem_resp_bits_rdata = io_dmem_mem_resp_bits_rdata; // @[src/main/scala/nutcore/NutCore.scala 161:13]
  assign io_dmem_cache_io_out_coh_req_valid = io_dmem_coh_req_valid; // @[src/main/scala/nutcore/NutCore.scala 161:13]
  assign io_dmem_cache_io_out_coh_req_bits_addr = io_dmem_coh_req_bits_addr; // @[src/main/scala/nutcore/NutCore.scala 161:13]
  assign io_dmem_cache_io_out_coh_req_bits_wdata = io_dmem_coh_req_bits_wdata; // @[src/main/scala/nutcore/NutCore.scala 161:13]
  assign io_dmem_cache_io_mmio_req_ready = mmioXbar_io_in_1_req_ready; // @[src/main/scala/nutcore/mem/Cache.scala 675:13]
  assign io_dmem_cache_io_mmio_resp_valid = mmioXbar_io_in_1_resp_valid; // @[src/main/scala/nutcore/mem/Cache.scala 675:13]
  assign io_dmem_cache_io_mmio_resp_bits_rdata = mmioXbar_io_in_1_resp_bits_rdata; // @[src/main/scala/nutcore/mem/Cache.scala 675:13]
  assign io_dmem_cache_DISPLAY_ENABLE = DISPLAY_ENABLE;
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_0_cf_instr <= 64'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h0 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_0_cf_instr <= 64'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_0_cf_instr <= _GEN_220;
        end
      end else begin
        dataBuffer_0_cf_instr <= _GEN_220;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_0_cf_pc <= 39'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h0 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_0_cf_pc <= 39'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_0_cf_pc <= _GEN_224;
        end
      end else begin
        dataBuffer_0_cf_pc <= _GEN_224;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_0_cf_pnpc <= 39'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h0 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_0_cf_pnpc <= 39'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_0_cf_pnpc <= _GEN_228;
        end
      end else begin
        dataBuffer_0_cf_pnpc <= _GEN_228;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_0_cf_exceptionVec_1 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h0 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_0_cf_exceptionVec_1 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_0_cf_exceptionVec_1 <= _GEN_248;
        end
      end else begin
        dataBuffer_0_cf_exceptionVec_1 <= _GEN_248;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_0_cf_exceptionVec_2 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h0 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_0_cf_exceptionVec_2 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_0_cf_exceptionVec_2 <= _GEN_252;
        end
      end else begin
        dataBuffer_0_cf_exceptionVec_2 <= _GEN_252;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_0_cf_exceptionVec_12 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h0 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_0_cf_exceptionVec_12 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_0_cf_exceptionVec_12 <= _GEN_292;
        end
      end else begin
        dataBuffer_0_cf_exceptionVec_12 <= _GEN_292;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_0_cf_intrVec_0 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h0 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_0_cf_intrVec_0 <= frontend_io_out_1_bits_cf_intrVec_0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_0_cf_intrVec_0 <= _GEN_308;
        end
      end else begin
        dataBuffer_0_cf_intrVec_0 <= _GEN_308;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_0_cf_intrVec_1 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h0 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_0_cf_intrVec_1 <= frontend_io_out_1_bits_cf_intrVec_1; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_0_cf_intrVec_1 <= _GEN_312;
        end
      end else begin
        dataBuffer_0_cf_intrVec_1 <= _GEN_312;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_0_cf_intrVec_2 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h0 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_0_cf_intrVec_2 <= frontend_io_out_1_bits_cf_intrVec_2; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_0_cf_intrVec_2 <= _GEN_316;
        end
      end else begin
        dataBuffer_0_cf_intrVec_2 <= _GEN_316;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_0_cf_intrVec_3 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h0 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_0_cf_intrVec_3 <= frontend_io_out_1_bits_cf_intrVec_3; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_0_cf_intrVec_3 <= _GEN_320;
        end
      end else begin
        dataBuffer_0_cf_intrVec_3 <= _GEN_320;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_0_cf_intrVec_4 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h0 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_0_cf_intrVec_4 <= frontend_io_out_1_bits_cf_intrVec_4; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_0_cf_intrVec_4 <= _GEN_324;
        end
      end else begin
        dataBuffer_0_cf_intrVec_4 <= _GEN_324;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_0_cf_intrVec_5 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h0 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_0_cf_intrVec_5 <= frontend_io_out_1_bits_cf_intrVec_5; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_0_cf_intrVec_5 <= _GEN_328;
        end
      end else begin
        dataBuffer_0_cf_intrVec_5 <= _GEN_328;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_0_cf_intrVec_6 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h0 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_0_cf_intrVec_6 <= frontend_io_out_1_bits_cf_intrVec_6; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_0_cf_intrVec_6 <= _GEN_332;
        end
      end else begin
        dataBuffer_0_cf_intrVec_6 <= _GEN_332;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_0_cf_intrVec_7 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h0 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_0_cf_intrVec_7 <= frontend_io_out_1_bits_cf_intrVec_7; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_0_cf_intrVec_7 <= _GEN_336;
        end
      end else begin
        dataBuffer_0_cf_intrVec_7 <= _GEN_336;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_0_cf_intrVec_8 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h0 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_0_cf_intrVec_8 <= frontend_io_out_1_bits_cf_intrVec_8; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_0_cf_intrVec_8 <= _GEN_340;
        end
      end else begin
        dataBuffer_0_cf_intrVec_8 <= _GEN_340;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_0_cf_intrVec_9 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h0 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_0_cf_intrVec_9 <= frontend_io_out_1_bits_cf_intrVec_9; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_0_cf_intrVec_9 <= _GEN_344;
        end
      end else begin
        dataBuffer_0_cf_intrVec_9 <= _GEN_344;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_0_cf_intrVec_10 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h0 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_0_cf_intrVec_10 <= frontend_io_out_1_bits_cf_intrVec_10; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_0_cf_intrVec_10 <= _GEN_348;
        end
      end else begin
        dataBuffer_0_cf_intrVec_10 <= _GEN_348;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_0_cf_intrVec_11 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h0 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_0_cf_intrVec_11 <= frontend_io_out_1_bits_cf_intrVec_11; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_0_cf_intrVec_11 <= _GEN_352;
        end
      end else begin
        dataBuffer_0_cf_intrVec_11 <= _GEN_352;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_0_cf_brIdx <= 4'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h0 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_0_cf_brIdx <= 4'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_0_cf_brIdx <= _GEN_356;
        end
      end else begin
        dataBuffer_0_cf_brIdx <= _GEN_356;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_0_cf_crossPageIPFFix <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h0 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_0_cf_crossPageIPFFix <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_0_cf_crossPageIPFFix <= _GEN_364;
        end
      end else begin
        dataBuffer_0_cf_crossPageIPFFix <= _GEN_364;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_0_ctrl_src1Type <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        dataBuffer_0_ctrl_src1Type <= 2'h0 == _T_4 | _GEN_376;
      end else if (enqueueFire_0) begin // @[src/main/scala/utils/PipelineVector.scala 45:29]
        dataBuffer_0_ctrl_src1Type <= _GEN_156;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_0_ctrl_src2Type <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        dataBuffer_0_ctrl_src2Type <= 2'h0 == _T_4 | _GEN_380;
      end else if (enqueueFire_0) begin // @[src/main/scala/utils/PipelineVector.scala 45:29]
        dataBuffer_0_ctrl_src2Type <= _GEN_160;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_0_ctrl_fuType <= 3'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h0 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_0_ctrl_fuType <= 3'h3; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_0_ctrl_fuType <= _GEN_384;
        end
      end else begin
        dataBuffer_0_ctrl_fuType <= _GEN_384;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_0_ctrl_fuOpType <= 7'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h0 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_0_ctrl_fuOpType <= 7'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_0_ctrl_fuOpType <= _GEN_388;
        end
      end else begin
        dataBuffer_0_ctrl_fuOpType <= _GEN_388;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_0_ctrl_rfSrc1 <= 5'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h0 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_0_ctrl_rfSrc1 <= 5'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_0_ctrl_rfSrc1 <= _GEN_392;
        end
      end else begin
        dataBuffer_0_ctrl_rfSrc1 <= _GEN_392;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_0_ctrl_rfSrc2 <= 5'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h0 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_0_ctrl_rfSrc2 <= 5'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_0_ctrl_rfSrc2 <= _GEN_396;
        end
      end else begin
        dataBuffer_0_ctrl_rfSrc2 <= _GEN_396;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_0_ctrl_rfWen <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h0 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_0_ctrl_rfWen <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_0_ctrl_rfWen <= _GEN_400;
        end
      end else begin
        dataBuffer_0_ctrl_rfWen <= _GEN_400;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_0_ctrl_rfDest <= 5'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h0 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_0_ctrl_rfDest <= 5'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_0_ctrl_rfDest <= _GEN_404;
        end
      end else begin
        dataBuffer_0_ctrl_rfDest <= _GEN_404;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_0_ctrl_isNutCoreTrap <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h0 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_0_ctrl_isNutCoreTrap <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_0_ctrl_isNutCoreTrap <= _GEN_408;
        end
      end else begin
        dataBuffer_0_ctrl_isNutCoreTrap <= _GEN_408;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_0_data_imm <= 64'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h0 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_0_data_imm <= 64'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_0_data_imm <= _GEN_436;
        end
      end else begin
        dataBuffer_0_data_imm <= _GEN_436;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_1_cf_instr <= 64'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h1 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_1_cf_instr <= 64'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_1_cf_instr <= _GEN_221;
        end
      end else begin
        dataBuffer_1_cf_instr <= _GEN_221;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_1_cf_pc <= 39'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h1 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_1_cf_pc <= 39'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_1_cf_pc <= _GEN_225;
        end
      end else begin
        dataBuffer_1_cf_pc <= _GEN_225;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_1_cf_pnpc <= 39'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h1 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_1_cf_pnpc <= 39'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_1_cf_pnpc <= _GEN_229;
        end
      end else begin
        dataBuffer_1_cf_pnpc <= _GEN_229;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_1_cf_exceptionVec_1 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h1 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_1_cf_exceptionVec_1 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_1_cf_exceptionVec_1 <= _GEN_249;
        end
      end else begin
        dataBuffer_1_cf_exceptionVec_1 <= _GEN_249;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_1_cf_exceptionVec_2 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h1 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_1_cf_exceptionVec_2 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_1_cf_exceptionVec_2 <= _GEN_253;
        end
      end else begin
        dataBuffer_1_cf_exceptionVec_2 <= _GEN_253;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_1_cf_exceptionVec_12 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h1 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_1_cf_exceptionVec_12 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_1_cf_exceptionVec_12 <= _GEN_293;
        end
      end else begin
        dataBuffer_1_cf_exceptionVec_12 <= _GEN_293;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_1_cf_intrVec_0 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h1 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_1_cf_intrVec_0 <= frontend_io_out_1_bits_cf_intrVec_0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_1_cf_intrVec_0 <= _GEN_309;
        end
      end else begin
        dataBuffer_1_cf_intrVec_0 <= _GEN_309;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_1_cf_intrVec_1 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h1 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_1_cf_intrVec_1 <= frontend_io_out_1_bits_cf_intrVec_1; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_1_cf_intrVec_1 <= _GEN_313;
        end
      end else begin
        dataBuffer_1_cf_intrVec_1 <= _GEN_313;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_1_cf_intrVec_2 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h1 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_1_cf_intrVec_2 <= frontend_io_out_1_bits_cf_intrVec_2; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_1_cf_intrVec_2 <= _GEN_317;
        end
      end else begin
        dataBuffer_1_cf_intrVec_2 <= _GEN_317;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_1_cf_intrVec_3 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h1 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_1_cf_intrVec_3 <= frontend_io_out_1_bits_cf_intrVec_3; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_1_cf_intrVec_3 <= _GEN_321;
        end
      end else begin
        dataBuffer_1_cf_intrVec_3 <= _GEN_321;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_1_cf_intrVec_4 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h1 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_1_cf_intrVec_4 <= frontend_io_out_1_bits_cf_intrVec_4; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_1_cf_intrVec_4 <= _GEN_325;
        end
      end else begin
        dataBuffer_1_cf_intrVec_4 <= _GEN_325;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_1_cf_intrVec_5 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h1 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_1_cf_intrVec_5 <= frontend_io_out_1_bits_cf_intrVec_5; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_1_cf_intrVec_5 <= _GEN_329;
        end
      end else begin
        dataBuffer_1_cf_intrVec_5 <= _GEN_329;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_1_cf_intrVec_6 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h1 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_1_cf_intrVec_6 <= frontend_io_out_1_bits_cf_intrVec_6; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_1_cf_intrVec_6 <= _GEN_333;
        end
      end else begin
        dataBuffer_1_cf_intrVec_6 <= _GEN_333;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_1_cf_intrVec_7 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h1 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_1_cf_intrVec_7 <= frontend_io_out_1_bits_cf_intrVec_7; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_1_cf_intrVec_7 <= _GEN_337;
        end
      end else begin
        dataBuffer_1_cf_intrVec_7 <= _GEN_337;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_1_cf_intrVec_8 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h1 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_1_cf_intrVec_8 <= frontend_io_out_1_bits_cf_intrVec_8; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_1_cf_intrVec_8 <= _GEN_341;
        end
      end else begin
        dataBuffer_1_cf_intrVec_8 <= _GEN_341;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_1_cf_intrVec_9 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h1 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_1_cf_intrVec_9 <= frontend_io_out_1_bits_cf_intrVec_9; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_1_cf_intrVec_9 <= _GEN_345;
        end
      end else begin
        dataBuffer_1_cf_intrVec_9 <= _GEN_345;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_1_cf_intrVec_10 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h1 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_1_cf_intrVec_10 <= frontend_io_out_1_bits_cf_intrVec_10; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_1_cf_intrVec_10 <= _GEN_349;
        end
      end else begin
        dataBuffer_1_cf_intrVec_10 <= _GEN_349;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_1_cf_intrVec_11 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h1 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_1_cf_intrVec_11 <= frontend_io_out_1_bits_cf_intrVec_11; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_1_cf_intrVec_11 <= _GEN_353;
        end
      end else begin
        dataBuffer_1_cf_intrVec_11 <= _GEN_353;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_1_cf_brIdx <= 4'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h1 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_1_cf_brIdx <= 4'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_1_cf_brIdx <= _GEN_357;
        end
      end else begin
        dataBuffer_1_cf_brIdx <= _GEN_357;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_1_cf_crossPageIPFFix <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h1 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_1_cf_crossPageIPFFix <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_1_cf_crossPageIPFFix <= _GEN_365;
        end
      end else begin
        dataBuffer_1_cf_crossPageIPFFix <= _GEN_365;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_1_ctrl_src1Type <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        dataBuffer_1_ctrl_src1Type <= 2'h1 == _T_4 | _GEN_377;
      end else if (enqueueFire_0) begin // @[src/main/scala/utils/PipelineVector.scala 45:29]
        dataBuffer_1_ctrl_src1Type <= _GEN_157;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_1_ctrl_src2Type <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        dataBuffer_1_ctrl_src2Type <= 2'h1 == _T_4 | _GEN_381;
      end else if (enqueueFire_0) begin // @[src/main/scala/utils/PipelineVector.scala 45:29]
        dataBuffer_1_ctrl_src2Type <= _GEN_161;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_1_ctrl_fuType <= 3'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h1 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_1_ctrl_fuType <= 3'h3; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_1_ctrl_fuType <= _GEN_385;
        end
      end else begin
        dataBuffer_1_ctrl_fuType <= _GEN_385;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_1_ctrl_fuOpType <= 7'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h1 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_1_ctrl_fuOpType <= 7'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_1_ctrl_fuOpType <= _GEN_389;
        end
      end else begin
        dataBuffer_1_ctrl_fuOpType <= _GEN_389;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_1_ctrl_rfSrc1 <= 5'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h1 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_1_ctrl_rfSrc1 <= 5'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_1_ctrl_rfSrc1 <= _GEN_393;
        end
      end else begin
        dataBuffer_1_ctrl_rfSrc1 <= _GEN_393;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_1_ctrl_rfSrc2 <= 5'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h1 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_1_ctrl_rfSrc2 <= 5'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_1_ctrl_rfSrc2 <= _GEN_397;
        end
      end else begin
        dataBuffer_1_ctrl_rfSrc2 <= _GEN_397;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_1_ctrl_rfWen <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h1 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_1_ctrl_rfWen <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_1_ctrl_rfWen <= _GEN_401;
        end
      end else begin
        dataBuffer_1_ctrl_rfWen <= _GEN_401;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_1_ctrl_rfDest <= 5'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h1 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_1_ctrl_rfDest <= 5'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_1_ctrl_rfDest <= _GEN_405;
        end
      end else begin
        dataBuffer_1_ctrl_rfDest <= _GEN_405;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_1_ctrl_isNutCoreTrap <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h1 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_1_ctrl_isNutCoreTrap <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_1_ctrl_isNutCoreTrap <= _GEN_409;
        end
      end else begin
        dataBuffer_1_ctrl_isNutCoreTrap <= _GEN_409;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_1_data_imm <= 64'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h1 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_1_data_imm <= 64'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_1_data_imm <= _GEN_437;
        end
      end else begin
        dataBuffer_1_data_imm <= _GEN_437;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_2_cf_instr <= 64'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h2 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_2_cf_instr <= 64'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_2_cf_instr <= _GEN_222;
        end
      end else begin
        dataBuffer_2_cf_instr <= _GEN_222;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_2_cf_pc <= 39'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h2 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_2_cf_pc <= 39'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_2_cf_pc <= _GEN_226;
        end
      end else begin
        dataBuffer_2_cf_pc <= _GEN_226;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_2_cf_pnpc <= 39'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h2 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_2_cf_pnpc <= 39'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_2_cf_pnpc <= _GEN_230;
        end
      end else begin
        dataBuffer_2_cf_pnpc <= _GEN_230;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_2_cf_exceptionVec_1 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h2 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_2_cf_exceptionVec_1 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_2_cf_exceptionVec_1 <= _GEN_250;
        end
      end else begin
        dataBuffer_2_cf_exceptionVec_1 <= _GEN_250;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_2_cf_exceptionVec_2 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h2 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_2_cf_exceptionVec_2 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_2_cf_exceptionVec_2 <= _GEN_254;
        end
      end else begin
        dataBuffer_2_cf_exceptionVec_2 <= _GEN_254;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_2_cf_exceptionVec_12 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h2 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_2_cf_exceptionVec_12 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_2_cf_exceptionVec_12 <= _GEN_294;
        end
      end else begin
        dataBuffer_2_cf_exceptionVec_12 <= _GEN_294;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_2_cf_intrVec_0 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h2 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_2_cf_intrVec_0 <= frontend_io_out_1_bits_cf_intrVec_0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_2_cf_intrVec_0 <= _GEN_310;
        end
      end else begin
        dataBuffer_2_cf_intrVec_0 <= _GEN_310;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_2_cf_intrVec_1 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h2 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_2_cf_intrVec_1 <= frontend_io_out_1_bits_cf_intrVec_1; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_2_cf_intrVec_1 <= _GEN_314;
        end
      end else begin
        dataBuffer_2_cf_intrVec_1 <= _GEN_314;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_2_cf_intrVec_2 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h2 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_2_cf_intrVec_2 <= frontend_io_out_1_bits_cf_intrVec_2; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_2_cf_intrVec_2 <= _GEN_318;
        end
      end else begin
        dataBuffer_2_cf_intrVec_2 <= _GEN_318;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_2_cf_intrVec_3 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h2 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_2_cf_intrVec_3 <= frontend_io_out_1_bits_cf_intrVec_3; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_2_cf_intrVec_3 <= _GEN_322;
        end
      end else begin
        dataBuffer_2_cf_intrVec_3 <= _GEN_322;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_2_cf_intrVec_4 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h2 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_2_cf_intrVec_4 <= frontend_io_out_1_bits_cf_intrVec_4; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_2_cf_intrVec_4 <= _GEN_326;
        end
      end else begin
        dataBuffer_2_cf_intrVec_4 <= _GEN_326;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_2_cf_intrVec_5 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h2 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_2_cf_intrVec_5 <= frontend_io_out_1_bits_cf_intrVec_5; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_2_cf_intrVec_5 <= _GEN_330;
        end
      end else begin
        dataBuffer_2_cf_intrVec_5 <= _GEN_330;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_2_cf_intrVec_6 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h2 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_2_cf_intrVec_6 <= frontend_io_out_1_bits_cf_intrVec_6; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_2_cf_intrVec_6 <= _GEN_334;
        end
      end else begin
        dataBuffer_2_cf_intrVec_6 <= _GEN_334;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_2_cf_intrVec_7 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h2 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_2_cf_intrVec_7 <= frontend_io_out_1_bits_cf_intrVec_7; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_2_cf_intrVec_7 <= _GEN_338;
        end
      end else begin
        dataBuffer_2_cf_intrVec_7 <= _GEN_338;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_2_cf_intrVec_8 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h2 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_2_cf_intrVec_8 <= frontend_io_out_1_bits_cf_intrVec_8; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_2_cf_intrVec_8 <= _GEN_342;
        end
      end else begin
        dataBuffer_2_cf_intrVec_8 <= _GEN_342;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_2_cf_intrVec_9 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h2 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_2_cf_intrVec_9 <= frontend_io_out_1_bits_cf_intrVec_9; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_2_cf_intrVec_9 <= _GEN_346;
        end
      end else begin
        dataBuffer_2_cf_intrVec_9 <= _GEN_346;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_2_cf_intrVec_10 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h2 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_2_cf_intrVec_10 <= frontend_io_out_1_bits_cf_intrVec_10; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_2_cf_intrVec_10 <= _GEN_350;
        end
      end else begin
        dataBuffer_2_cf_intrVec_10 <= _GEN_350;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_2_cf_intrVec_11 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h2 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_2_cf_intrVec_11 <= frontend_io_out_1_bits_cf_intrVec_11; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_2_cf_intrVec_11 <= _GEN_354;
        end
      end else begin
        dataBuffer_2_cf_intrVec_11 <= _GEN_354;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_2_cf_brIdx <= 4'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h2 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_2_cf_brIdx <= 4'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_2_cf_brIdx <= _GEN_358;
        end
      end else begin
        dataBuffer_2_cf_brIdx <= _GEN_358;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_2_cf_crossPageIPFFix <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h2 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_2_cf_crossPageIPFFix <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_2_cf_crossPageIPFFix <= _GEN_366;
        end
      end else begin
        dataBuffer_2_cf_crossPageIPFFix <= _GEN_366;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_2_ctrl_src1Type <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        dataBuffer_2_ctrl_src1Type <= 2'h2 == _T_4 | _GEN_378;
      end else if (enqueueFire_0) begin // @[src/main/scala/utils/PipelineVector.scala 45:29]
        dataBuffer_2_ctrl_src1Type <= _GEN_158;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_2_ctrl_src2Type <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        dataBuffer_2_ctrl_src2Type <= 2'h2 == _T_4 | _GEN_382;
      end else if (enqueueFire_0) begin // @[src/main/scala/utils/PipelineVector.scala 45:29]
        dataBuffer_2_ctrl_src2Type <= _GEN_162;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_2_ctrl_fuType <= 3'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h2 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_2_ctrl_fuType <= 3'h3; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_2_ctrl_fuType <= _GEN_386;
        end
      end else begin
        dataBuffer_2_ctrl_fuType <= _GEN_386;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_2_ctrl_fuOpType <= 7'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h2 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_2_ctrl_fuOpType <= 7'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_2_ctrl_fuOpType <= _GEN_390;
        end
      end else begin
        dataBuffer_2_ctrl_fuOpType <= _GEN_390;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_2_ctrl_rfSrc1 <= 5'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h2 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_2_ctrl_rfSrc1 <= 5'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_2_ctrl_rfSrc1 <= _GEN_394;
        end
      end else begin
        dataBuffer_2_ctrl_rfSrc1 <= _GEN_394;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_2_ctrl_rfSrc2 <= 5'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h2 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_2_ctrl_rfSrc2 <= 5'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_2_ctrl_rfSrc2 <= _GEN_398;
        end
      end else begin
        dataBuffer_2_ctrl_rfSrc2 <= _GEN_398;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_2_ctrl_rfWen <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h2 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_2_ctrl_rfWen <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_2_ctrl_rfWen <= _GEN_402;
        end
      end else begin
        dataBuffer_2_ctrl_rfWen <= _GEN_402;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_2_ctrl_rfDest <= 5'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h2 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_2_ctrl_rfDest <= 5'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_2_ctrl_rfDest <= _GEN_406;
        end
      end else begin
        dataBuffer_2_ctrl_rfDest <= _GEN_406;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_2_ctrl_isNutCoreTrap <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h2 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_2_ctrl_isNutCoreTrap <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_2_ctrl_isNutCoreTrap <= _GEN_410;
        end
      end else begin
        dataBuffer_2_ctrl_isNutCoreTrap <= _GEN_410;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_2_data_imm <= 64'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h2 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_2_data_imm <= 64'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_2_data_imm <= _GEN_438;
        end
      end else begin
        dataBuffer_2_data_imm <= _GEN_438;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_3_cf_instr <= 64'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h3 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_3_cf_instr <= 64'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_3_cf_instr <= _GEN_223;
        end
      end else begin
        dataBuffer_3_cf_instr <= _GEN_223;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_3_cf_pc <= 39'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h3 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_3_cf_pc <= 39'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_3_cf_pc <= _GEN_227;
        end
      end else begin
        dataBuffer_3_cf_pc <= _GEN_227;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_3_cf_pnpc <= 39'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h3 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_3_cf_pnpc <= 39'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_3_cf_pnpc <= _GEN_231;
        end
      end else begin
        dataBuffer_3_cf_pnpc <= _GEN_231;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_3_cf_exceptionVec_1 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h3 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_3_cf_exceptionVec_1 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_3_cf_exceptionVec_1 <= _GEN_251;
        end
      end else begin
        dataBuffer_3_cf_exceptionVec_1 <= _GEN_251;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_3_cf_exceptionVec_2 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h3 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_3_cf_exceptionVec_2 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_3_cf_exceptionVec_2 <= _GEN_255;
        end
      end else begin
        dataBuffer_3_cf_exceptionVec_2 <= _GEN_255;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_3_cf_exceptionVec_12 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h3 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_3_cf_exceptionVec_12 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_3_cf_exceptionVec_12 <= _GEN_295;
        end
      end else begin
        dataBuffer_3_cf_exceptionVec_12 <= _GEN_295;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_3_cf_intrVec_0 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h3 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_3_cf_intrVec_0 <= frontend_io_out_1_bits_cf_intrVec_0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_3_cf_intrVec_0 <= _GEN_311;
        end
      end else begin
        dataBuffer_3_cf_intrVec_0 <= _GEN_311;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_3_cf_intrVec_1 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h3 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_3_cf_intrVec_1 <= frontend_io_out_1_bits_cf_intrVec_1; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_3_cf_intrVec_1 <= _GEN_315;
        end
      end else begin
        dataBuffer_3_cf_intrVec_1 <= _GEN_315;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_3_cf_intrVec_2 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h3 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_3_cf_intrVec_2 <= frontend_io_out_1_bits_cf_intrVec_2; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_3_cf_intrVec_2 <= _GEN_319;
        end
      end else begin
        dataBuffer_3_cf_intrVec_2 <= _GEN_319;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_3_cf_intrVec_3 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h3 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_3_cf_intrVec_3 <= frontend_io_out_1_bits_cf_intrVec_3; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_3_cf_intrVec_3 <= _GEN_323;
        end
      end else begin
        dataBuffer_3_cf_intrVec_3 <= _GEN_323;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_3_cf_intrVec_4 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h3 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_3_cf_intrVec_4 <= frontend_io_out_1_bits_cf_intrVec_4; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_3_cf_intrVec_4 <= _GEN_327;
        end
      end else begin
        dataBuffer_3_cf_intrVec_4 <= _GEN_327;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_3_cf_intrVec_5 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h3 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_3_cf_intrVec_5 <= frontend_io_out_1_bits_cf_intrVec_5; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_3_cf_intrVec_5 <= _GEN_331;
        end
      end else begin
        dataBuffer_3_cf_intrVec_5 <= _GEN_331;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_3_cf_intrVec_6 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h3 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_3_cf_intrVec_6 <= frontend_io_out_1_bits_cf_intrVec_6; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_3_cf_intrVec_6 <= _GEN_335;
        end
      end else begin
        dataBuffer_3_cf_intrVec_6 <= _GEN_335;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_3_cf_intrVec_7 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h3 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_3_cf_intrVec_7 <= frontend_io_out_1_bits_cf_intrVec_7; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_3_cf_intrVec_7 <= _GEN_339;
        end
      end else begin
        dataBuffer_3_cf_intrVec_7 <= _GEN_339;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_3_cf_intrVec_8 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h3 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_3_cf_intrVec_8 <= frontend_io_out_1_bits_cf_intrVec_8; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_3_cf_intrVec_8 <= _GEN_343;
        end
      end else begin
        dataBuffer_3_cf_intrVec_8 <= _GEN_343;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_3_cf_intrVec_9 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h3 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_3_cf_intrVec_9 <= frontend_io_out_1_bits_cf_intrVec_9; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_3_cf_intrVec_9 <= _GEN_347;
        end
      end else begin
        dataBuffer_3_cf_intrVec_9 <= _GEN_347;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_3_cf_intrVec_10 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h3 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_3_cf_intrVec_10 <= frontend_io_out_1_bits_cf_intrVec_10; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_3_cf_intrVec_10 <= _GEN_351;
        end
      end else begin
        dataBuffer_3_cf_intrVec_10 <= _GEN_351;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_3_cf_intrVec_11 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h3 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_3_cf_intrVec_11 <= frontend_io_out_1_bits_cf_intrVec_11; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_3_cf_intrVec_11 <= _GEN_355;
        end
      end else begin
        dataBuffer_3_cf_intrVec_11 <= _GEN_355;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_3_cf_brIdx <= 4'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h3 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_3_cf_brIdx <= 4'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_3_cf_brIdx <= _GEN_359;
        end
      end else begin
        dataBuffer_3_cf_brIdx <= _GEN_359;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_3_cf_crossPageIPFFix <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h3 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_3_cf_crossPageIPFFix <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_3_cf_crossPageIPFFix <= _GEN_367;
        end
      end else begin
        dataBuffer_3_cf_crossPageIPFFix <= _GEN_367;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_3_ctrl_src1Type <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        dataBuffer_3_ctrl_src1Type <= 2'h3 == _T_4 | _GEN_379;
      end else if (enqueueFire_0) begin // @[src/main/scala/utils/PipelineVector.scala 45:29]
        dataBuffer_3_ctrl_src1Type <= _GEN_159;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_3_ctrl_src2Type <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        dataBuffer_3_ctrl_src2Type <= 2'h3 == _T_4 | _GEN_383;
      end else if (enqueueFire_0) begin // @[src/main/scala/utils/PipelineVector.scala 45:29]
        dataBuffer_3_ctrl_src2Type <= _GEN_163;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_3_ctrl_fuType <= 3'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h3 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_3_ctrl_fuType <= 3'h3; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_3_ctrl_fuType <= _GEN_387;
        end
      end else begin
        dataBuffer_3_ctrl_fuType <= _GEN_387;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_3_ctrl_fuOpType <= 7'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h3 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_3_ctrl_fuOpType <= 7'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_3_ctrl_fuOpType <= _GEN_391;
        end
      end else begin
        dataBuffer_3_ctrl_fuOpType <= _GEN_391;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_3_ctrl_rfSrc1 <= 5'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h3 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_3_ctrl_rfSrc1 <= 5'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_3_ctrl_rfSrc1 <= _GEN_395;
        end
      end else begin
        dataBuffer_3_ctrl_rfSrc1 <= _GEN_395;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_3_ctrl_rfSrc2 <= 5'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h3 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_3_ctrl_rfSrc2 <= 5'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_3_ctrl_rfSrc2 <= _GEN_399;
        end
      end else begin
        dataBuffer_3_ctrl_rfSrc2 <= _GEN_399;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_3_ctrl_rfWen <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h3 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_3_ctrl_rfWen <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_3_ctrl_rfWen <= _GEN_403;
        end
      end else begin
        dataBuffer_3_ctrl_rfWen <= _GEN_403;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_3_ctrl_rfDest <= 5'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h3 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_3_ctrl_rfDest <= 5'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_3_ctrl_rfDest <= _GEN_407;
        end
      end else begin
        dataBuffer_3_ctrl_rfDest <= _GEN_407;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_3_ctrl_isNutCoreTrap <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h3 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_3_ctrl_isNutCoreTrap <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_3_ctrl_isNutCoreTrap <= _GEN_411;
        end
      end else begin
        dataBuffer_3_ctrl_isNutCoreTrap <= _GEN_411;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_3_data_imm <= 64'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h3 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_3_data_imm <= 64'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_3_data_imm <= _GEN_439;
        end
      end else begin
        dataBuffer_3_data_imm <= _GEN_439;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 30:33]
      ringBufferHead <= 2'h0; // @[src/main/scala/utils/PipelineVector.scala 30:33]
    end else if (frontend_io_flushVec[1]) begin // @[src/main/scala/utils/PipelineVector.scala 71:16]
      ringBufferHead <= 2'h0; // @[src/main/scala/utils/PipelineVector.scala 72:24]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      ringBufferHead <= _ringBufferHead_T_1; // @[src/main/scala/utils/PipelineVector.scala 47:24]
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 31:33]
      ringBufferTail <= 2'h0; // @[src/main/scala/utils/PipelineVector.scala 31:33]
    end else if (frontend_io_flushVec[1]) begin // @[src/main/scala/utils/PipelineVector.scala 71:16]
      ringBufferTail <= 2'h0; // @[src/main/scala/utils/PipelineVector.scala 73:24]
    end else if (dequeueFire) begin // @[src/main/scala/utils/PipelineVector.scala 66:22]
      ringBufferTail <= _ringBufferTail_T_1; // @[src/main/scala/utils/PipelineVector.scala 67:24]
    end
    if (reset) begin // @[src/main/scala/utils/GTimer.scala 24:20]
      c <= 64'h0; // @[src/main/scala/utils/GTimer.scala 24:20]
    end else begin
      c <= _c_T_1; // @[src/main/scala/utils/GTimer.scala 25:7]
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & ~reset) begin
          $fwrite(32'h80000002,"[DPQ] size %x head %x tail %x enq %x deq %x\n",_GEN_12[2:0],ringBufferHead,
            ringBufferTail,enqueueSize,dequeueSize); // @[src/main/scala/utils/PipelineVector.scala 77:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_11) begin
          $fwrite(32'h80000002,"[%d] NutCore: ",c); // @[src/main/scala/utils/Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_11) begin
          $fwrite(32'h80000002,"------------------------ BACKEND ------------------------\n"); // @[src/main/scala/utils/Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  dataBuffer_0_cf_instr = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  dataBuffer_0_cf_pc = _RAND_1[38:0];
  _RAND_2 = {2{`RANDOM}};
  dataBuffer_0_cf_pnpc = _RAND_2[38:0];
  _RAND_3 = {1{`RANDOM}};
  dataBuffer_0_cf_exceptionVec_1 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  dataBuffer_0_cf_exceptionVec_2 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  dataBuffer_0_cf_exceptionVec_12 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  dataBuffer_0_cf_intrVec_0 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  dataBuffer_0_cf_intrVec_1 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  dataBuffer_0_cf_intrVec_2 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  dataBuffer_0_cf_intrVec_3 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  dataBuffer_0_cf_intrVec_4 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  dataBuffer_0_cf_intrVec_5 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  dataBuffer_0_cf_intrVec_6 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  dataBuffer_0_cf_intrVec_7 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  dataBuffer_0_cf_intrVec_8 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  dataBuffer_0_cf_intrVec_9 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  dataBuffer_0_cf_intrVec_10 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  dataBuffer_0_cf_intrVec_11 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  dataBuffer_0_cf_brIdx = _RAND_18[3:0];
  _RAND_19 = {1{`RANDOM}};
  dataBuffer_0_cf_crossPageIPFFix = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  dataBuffer_0_ctrl_src1Type = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  dataBuffer_0_ctrl_src2Type = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  dataBuffer_0_ctrl_fuType = _RAND_22[2:0];
  _RAND_23 = {1{`RANDOM}};
  dataBuffer_0_ctrl_fuOpType = _RAND_23[6:0];
  _RAND_24 = {1{`RANDOM}};
  dataBuffer_0_ctrl_rfSrc1 = _RAND_24[4:0];
  _RAND_25 = {1{`RANDOM}};
  dataBuffer_0_ctrl_rfSrc2 = _RAND_25[4:0];
  _RAND_26 = {1{`RANDOM}};
  dataBuffer_0_ctrl_rfWen = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  dataBuffer_0_ctrl_rfDest = _RAND_27[4:0];
  _RAND_28 = {1{`RANDOM}};
  dataBuffer_0_ctrl_isNutCoreTrap = _RAND_28[0:0];
  _RAND_29 = {2{`RANDOM}};
  dataBuffer_0_data_imm = _RAND_29[63:0];
  _RAND_30 = {2{`RANDOM}};
  dataBuffer_1_cf_instr = _RAND_30[63:0];
  _RAND_31 = {2{`RANDOM}};
  dataBuffer_1_cf_pc = _RAND_31[38:0];
  _RAND_32 = {2{`RANDOM}};
  dataBuffer_1_cf_pnpc = _RAND_32[38:0];
  _RAND_33 = {1{`RANDOM}};
  dataBuffer_1_cf_exceptionVec_1 = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  dataBuffer_1_cf_exceptionVec_2 = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  dataBuffer_1_cf_exceptionVec_12 = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  dataBuffer_1_cf_intrVec_0 = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  dataBuffer_1_cf_intrVec_1 = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  dataBuffer_1_cf_intrVec_2 = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  dataBuffer_1_cf_intrVec_3 = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  dataBuffer_1_cf_intrVec_4 = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  dataBuffer_1_cf_intrVec_5 = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  dataBuffer_1_cf_intrVec_6 = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  dataBuffer_1_cf_intrVec_7 = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  dataBuffer_1_cf_intrVec_8 = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  dataBuffer_1_cf_intrVec_9 = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  dataBuffer_1_cf_intrVec_10 = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  dataBuffer_1_cf_intrVec_11 = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  dataBuffer_1_cf_brIdx = _RAND_48[3:0];
  _RAND_49 = {1{`RANDOM}};
  dataBuffer_1_cf_crossPageIPFFix = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  dataBuffer_1_ctrl_src1Type = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  dataBuffer_1_ctrl_src2Type = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  dataBuffer_1_ctrl_fuType = _RAND_52[2:0];
  _RAND_53 = {1{`RANDOM}};
  dataBuffer_1_ctrl_fuOpType = _RAND_53[6:0];
  _RAND_54 = {1{`RANDOM}};
  dataBuffer_1_ctrl_rfSrc1 = _RAND_54[4:0];
  _RAND_55 = {1{`RANDOM}};
  dataBuffer_1_ctrl_rfSrc2 = _RAND_55[4:0];
  _RAND_56 = {1{`RANDOM}};
  dataBuffer_1_ctrl_rfWen = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  dataBuffer_1_ctrl_rfDest = _RAND_57[4:0];
  _RAND_58 = {1{`RANDOM}};
  dataBuffer_1_ctrl_isNutCoreTrap = _RAND_58[0:0];
  _RAND_59 = {2{`RANDOM}};
  dataBuffer_1_data_imm = _RAND_59[63:0];
  _RAND_60 = {2{`RANDOM}};
  dataBuffer_2_cf_instr = _RAND_60[63:0];
  _RAND_61 = {2{`RANDOM}};
  dataBuffer_2_cf_pc = _RAND_61[38:0];
  _RAND_62 = {2{`RANDOM}};
  dataBuffer_2_cf_pnpc = _RAND_62[38:0];
  _RAND_63 = {1{`RANDOM}};
  dataBuffer_2_cf_exceptionVec_1 = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  dataBuffer_2_cf_exceptionVec_2 = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  dataBuffer_2_cf_exceptionVec_12 = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  dataBuffer_2_cf_intrVec_0 = _RAND_66[0:0];
  _RAND_67 = {1{`RANDOM}};
  dataBuffer_2_cf_intrVec_1 = _RAND_67[0:0];
  _RAND_68 = {1{`RANDOM}};
  dataBuffer_2_cf_intrVec_2 = _RAND_68[0:0];
  _RAND_69 = {1{`RANDOM}};
  dataBuffer_2_cf_intrVec_3 = _RAND_69[0:0];
  _RAND_70 = {1{`RANDOM}};
  dataBuffer_2_cf_intrVec_4 = _RAND_70[0:0];
  _RAND_71 = {1{`RANDOM}};
  dataBuffer_2_cf_intrVec_5 = _RAND_71[0:0];
  _RAND_72 = {1{`RANDOM}};
  dataBuffer_2_cf_intrVec_6 = _RAND_72[0:0];
  _RAND_73 = {1{`RANDOM}};
  dataBuffer_2_cf_intrVec_7 = _RAND_73[0:0];
  _RAND_74 = {1{`RANDOM}};
  dataBuffer_2_cf_intrVec_8 = _RAND_74[0:0];
  _RAND_75 = {1{`RANDOM}};
  dataBuffer_2_cf_intrVec_9 = _RAND_75[0:0];
  _RAND_76 = {1{`RANDOM}};
  dataBuffer_2_cf_intrVec_10 = _RAND_76[0:0];
  _RAND_77 = {1{`RANDOM}};
  dataBuffer_2_cf_intrVec_11 = _RAND_77[0:0];
  _RAND_78 = {1{`RANDOM}};
  dataBuffer_2_cf_brIdx = _RAND_78[3:0];
  _RAND_79 = {1{`RANDOM}};
  dataBuffer_2_cf_crossPageIPFFix = _RAND_79[0:0];
  _RAND_80 = {1{`RANDOM}};
  dataBuffer_2_ctrl_src1Type = _RAND_80[0:0];
  _RAND_81 = {1{`RANDOM}};
  dataBuffer_2_ctrl_src2Type = _RAND_81[0:0];
  _RAND_82 = {1{`RANDOM}};
  dataBuffer_2_ctrl_fuType = _RAND_82[2:0];
  _RAND_83 = {1{`RANDOM}};
  dataBuffer_2_ctrl_fuOpType = _RAND_83[6:0];
  _RAND_84 = {1{`RANDOM}};
  dataBuffer_2_ctrl_rfSrc1 = _RAND_84[4:0];
  _RAND_85 = {1{`RANDOM}};
  dataBuffer_2_ctrl_rfSrc2 = _RAND_85[4:0];
  _RAND_86 = {1{`RANDOM}};
  dataBuffer_2_ctrl_rfWen = _RAND_86[0:0];
  _RAND_87 = {1{`RANDOM}};
  dataBuffer_2_ctrl_rfDest = _RAND_87[4:0];
  _RAND_88 = {1{`RANDOM}};
  dataBuffer_2_ctrl_isNutCoreTrap = _RAND_88[0:0];
  _RAND_89 = {2{`RANDOM}};
  dataBuffer_2_data_imm = _RAND_89[63:0];
  _RAND_90 = {2{`RANDOM}};
  dataBuffer_3_cf_instr = _RAND_90[63:0];
  _RAND_91 = {2{`RANDOM}};
  dataBuffer_3_cf_pc = _RAND_91[38:0];
  _RAND_92 = {2{`RANDOM}};
  dataBuffer_3_cf_pnpc = _RAND_92[38:0];
  _RAND_93 = {1{`RANDOM}};
  dataBuffer_3_cf_exceptionVec_1 = _RAND_93[0:0];
  _RAND_94 = {1{`RANDOM}};
  dataBuffer_3_cf_exceptionVec_2 = _RAND_94[0:0];
  _RAND_95 = {1{`RANDOM}};
  dataBuffer_3_cf_exceptionVec_12 = _RAND_95[0:0];
  _RAND_96 = {1{`RANDOM}};
  dataBuffer_3_cf_intrVec_0 = _RAND_96[0:0];
  _RAND_97 = {1{`RANDOM}};
  dataBuffer_3_cf_intrVec_1 = _RAND_97[0:0];
  _RAND_98 = {1{`RANDOM}};
  dataBuffer_3_cf_intrVec_2 = _RAND_98[0:0];
  _RAND_99 = {1{`RANDOM}};
  dataBuffer_3_cf_intrVec_3 = _RAND_99[0:0];
  _RAND_100 = {1{`RANDOM}};
  dataBuffer_3_cf_intrVec_4 = _RAND_100[0:0];
  _RAND_101 = {1{`RANDOM}};
  dataBuffer_3_cf_intrVec_5 = _RAND_101[0:0];
  _RAND_102 = {1{`RANDOM}};
  dataBuffer_3_cf_intrVec_6 = _RAND_102[0:0];
  _RAND_103 = {1{`RANDOM}};
  dataBuffer_3_cf_intrVec_7 = _RAND_103[0:0];
  _RAND_104 = {1{`RANDOM}};
  dataBuffer_3_cf_intrVec_8 = _RAND_104[0:0];
  _RAND_105 = {1{`RANDOM}};
  dataBuffer_3_cf_intrVec_9 = _RAND_105[0:0];
  _RAND_106 = {1{`RANDOM}};
  dataBuffer_3_cf_intrVec_10 = _RAND_106[0:0];
  _RAND_107 = {1{`RANDOM}};
  dataBuffer_3_cf_intrVec_11 = _RAND_107[0:0];
  _RAND_108 = {1{`RANDOM}};
  dataBuffer_3_cf_brIdx = _RAND_108[3:0];
  _RAND_109 = {1{`RANDOM}};
  dataBuffer_3_cf_crossPageIPFFix = _RAND_109[0:0];
  _RAND_110 = {1{`RANDOM}};
  dataBuffer_3_ctrl_src1Type = _RAND_110[0:0];
  _RAND_111 = {1{`RANDOM}};
  dataBuffer_3_ctrl_src2Type = _RAND_111[0:0];
  _RAND_112 = {1{`RANDOM}};
  dataBuffer_3_ctrl_fuType = _RAND_112[2:0];
  _RAND_113 = {1{`RANDOM}};
  dataBuffer_3_ctrl_fuOpType = _RAND_113[6:0];
  _RAND_114 = {1{`RANDOM}};
  dataBuffer_3_ctrl_rfSrc1 = _RAND_114[4:0];
  _RAND_115 = {1{`RANDOM}};
  dataBuffer_3_ctrl_rfSrc2 = _RAND_115[4:0];
  _RAND_116 = {1{`RANDOM}};
  dataBuffer_3_ctrl_rfWen = _RAND_116[0:0];
  _RAND_117 = {1{`RANDOM}};
  dataBuffer_3_ctrl_rfDest = _RAND_117[4:0];
  _RAND_118 = {1{`RANDOM}};
  dataBuffer_3_ctrl_isNutCoreTrap = _RAND_118[0:0];
  _RAND_119 = {2{`RANDOM}};
  dataBuffer_3_data_imm = _RAND_119[63:0];
  _RAND_120 = {1{`RANDOM}};
  ringBufferHead = _RAND_120[1:0];
  _RAND_121 = {1{`RANDOM}};
  ringBufferTail = _RAND_121[1:0];
  _RAND_122 = {2{`RANDOM}};
  c = _RAND_122[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module CoherenceManager(
  input         clock,
  input         reset,
  output        io_in_req_ready, // @[src/main/scala/system/Coherence.scala 31:14]
  input         io_in_req_valid, // @[src/main/scala/system/Coherence.scala 31:14]
  input  [31:0] io_in_req_bits_addr, // @[src/main/scala/system/Coherence.scala 31:14]
  input  [3:0]  io_in_req_bits_cmd, // @[src/main/scala/system/Coherence.scala 31:14]
  input  [63:0] io_in_req_bits_wdata, // @[src/main/scala/system/Coherence.scala 31:14]
  output        io_in_resp_valid, // @[src/main/scala/system/Coherence.scala 31:14]
  output [3:0]  io_in_resp_bits_cmd, // @[src/main/scala/system/Coherence.scala 31:14]
  output [63:0] io_in_resp_bits_rdata, // @[src/main/scala/system/Coherence.scala 31:14]
  input         io_out_mem_req_ready, // @[src/main/scala/system/Coherence.scala 31:14]
  output        io_out_mem_req_valid, // @[src/main/scala/system/Coherence.scala 31:14]
  output [31:0] io_out_mem_req_bits_addr, // @[src/main/scala/system/Coherence.scala 31:14]
  output [3:0]  io_out_mem_req_bits_cmd, // @[src/main/scala/system/Coherence.scala 31:14]
  output [63:0] io_out_mem_req_bits_wdata, // @[src/main/scala/system/Coherence.scala 31:14]
  output        io_out_mem_resp_ready, // @[src/main/scala/system/Coherence.scala 31:14]
  input         io_out_mem_resp_valid, // @[src/main/scala/system/Coherence.scala 31:14]
  input  [3:0]  io_out_mem_resp_bits_cmd, // @[src/main/scala/system/Coherence.scala 31:14]
  input  [63:0] io_out_mem_resp_bits_rdata, // @[src/main/scala/system/Coherence.scala 31:14]
  input         io_out_coh_req_ready, // @[src/main/scala/system/Coherence.scala 31:14]
  output        io_out_coh_req_valid, // @[src/main/scala/system/Coherence.scala 31:14]
  output [31:0] io_out_coh_req_bits_addr, // @[src/main/scala/system/Coherence.scala 31:14]
  output [63:0] io_out_coh_req_bits_wdata, // @[src/main/scala/system/Coherence.scala 31:14]
  output        io_out_coh_resp_ready, // @[src/main/scala/system/Coherence.scala 31:14]
  input         io_out_coh_resp_valid, // @[src/main/scala/system/Coherence.scala 31:14]
  input  [3:0]  io_out_coh_resp_bits_cmd, // @[src/main/scala/system/Coherence.scala 31:14]
  input  [63:0] io_out_coh_resp_bits_rdata // @[src/main/scala/system/Coherence.scala 31:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [63:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  reg [2:0] state; // @[src/main/scala/system/Coherence.scala 45:22]
  wire  inflight = state != 3'h0; // @[src/main/scala/system/Coherence.scala 46:24]
  wire  _T_1 = ~io_in_req_bits_cmd[0]; // @[src/main/scala/bus/simplebus/SimpleBus.scala 73:18]
  wire  _T_4 = ~io_in_req_bits_cmd[0] & ~io_in_req_bits_cmd[3]; // @[src/main/scala/bus/simplebus/SimpleBus.scala 73:26]
  wire  _reqLatch_T = ~inflight; // @[src/main/scala/system/Coherence.scala 52:42]
  reg [31:0] reqLatch_addr; // @[src/main/scala/system/Coherence.scala 52:27]
  reg [3:0] reqLatch_cmd; // @[src/main/scala/system/Coherence.scala 52:27]
  reg [63:0] reqLatch_wdata; // @[src/main/scala/system/Coherence.scala 52:27]
  wire  _io_out_mem_req_valid_T_1 = io_in_req_valid & _reqLatch_T; // @[src/main/scala/system/Coherence.scala 65:43]
  wire  _GEN_5 = _T_4 & _io_out_mem_req_valid_T_1; // @[src/main/scala/system/Coherence.scala 63:24 67:39 68:26]
  wire  _GEN_6 = _T_4 & (io_out_coh_req_ready & _reqLatch_T); // @[src/main/scala/system/Coherence.scala 62:17 67:39 69:19]
  wire  _GEN_7 = io_in_req_bits_cmd[0] & (io_in_req_valid & _reqLatch_T); // @[src/main/scala/system/Coherence.scala 61:24 64:61 65:26]
  wire  _T_21 = io_in_req_ready & io_in_req_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  wire  _T_27 = io_in_req_bits_cmd == 4'h7; // @[src/main/scala/bus/simplebus/SimpleBus.scala 78:27]
  wire [2:0] _GEN_10 = _T_27 ? 3'h5 : state; // @[src/main/scala/system/Coherence.scala 45:22 78:{48,56}]
  wire  _T_29 = io_out_coh_resp_ready & io_out_coh_resp_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  wire  _state_T_1 = io_out_coh_resp_bits_cmd == 4'hc; // @[src/main/scala/bus/simplebus/SimpleBus.scala 92:24]
  wire [2:0] _state_T_2 = _state_T_1 ? 3'h2 : 3'h3; // @[src/main/scala/system/Coherence.scala 83:21]
  wire  _T_32 = io_in_resp_bits_cmd == 4'h6; // @[src/main/scala/bus/simplebus/SimpleBus.scala 91:24]
  wire [2:0] _GEN_14 = io_in_resp_valid & _T_32 ? 3'h0 : state; // @[src/main/scala/system/Coherence.scala 45:22 89:{56,64}]
  wire  _T_35 = io_out_mem_req_ready & io_out_mem_req_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  wire [2:0] _GEN_15 = _T_35 ? 3'h4 : state; // @[src/main/scala/system/Coherence.scala 45:22 94:{34,42}]
  wire  _T_37 = io_out_mem_resp_ready & io_out_mem_resp_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  wire  _T_38 = io_out_mem_resp_bits_cmd == 4'h6; // @[src/main/scala/bus/simplebus/SimpleBus.scala 91:24]
  wire [2:0] _GEN_16 = _T_37 & _T_38 ? 3'h0 : state; // @[src/main/scala/system/Coherence.scala 45:22 96:{89,97}]
  wire [2:0] _GEN_17 = _T_37 ? 3'h0 : state; // @[src/main/scala/system/Coherence.scala 45:22 97:{55,63}]
  wire [2:0] _GEN_18 = 3'h5 == state ? _GEN_17 : state; // @[src/main/scala/system/Coherence.scala 74:18 45:22]
  wire [2:0] _GEN_19 = 3'h4 == state ? _GEN_16 : _GEN_18; // @[src/main/scala/system/Coherence.scala 74:18]
  wire [31:0] _GEN_20 = 3'h3 == state ? reqLatch_addr : io_in_req_bits_addr; // @[src/main/scala/system/Coherence.scala 74:18 59:23 92:27]
  wire [3:0] _GEN_22 = 3'h3 == state ? reqLatch_cmd : io_in_req_bits_cmd; // @[src/main/scala/system/Coherence.scala 74:18 59:23 92:27]
  wire [63:0] _GEN_24 = 3'h3 == state ? reqLatch_wdata : io_in_req_bits_wdata; // @[src/main/scala/system/Coherence.scala 74:18 59:23 92:27]
  wire  _GEN_25 = 3'h3 == state | _GEN_7; // @[src/main/scala/system/Coherence.scala 74:18 93:28]
  wire [2:0] _GEN_26 = 3'h3 == state ? _GEN_15 : _GEN_19; // @[src/main/scala/system/Coherence.scala 74:18]
  wire  _GEN_28 = 3'h2 == state ? io_out_coh_resp_valid : io_out_mem_resp_valid; // @[src/main/scala/system/Coherence.scala 72:14 74:18 88:16]
  wire [3:0] _GEN_29 = 3'h2 == state ? io_out_coh_resp_bits_cmd : io_out_mem_resp_bits_cmd; // @[src/main/scala/system/Coherence.scala 72:14 74:18 88:16]
  wire [63:0] _GEN_30 = 3'h2 == state ? io_out_coh_resp_bits_rdata : io_out_mem_resp_bits_rdata; // @[src/main/scala/system/Coherence.scala 72:14 74:18 88:16]
  wire [31:0] _GEN_32 = 3'h2 == state ? io_in_req_bits_addr : _GEN_20; // @[src/main/scala/system/Coherence.scala 74:18 59:23]
  wire [3:0] _GEN_34 = 3'h2 == state ? io_in_req_bits_cmd : _GEN_22; // @[src/main/scala/system/Coherence.scala 74:18 59:23]
  wire [63:0] _GEN_36 = 3'h2 == state ? io_in_req_bits_wdata : _GEN_24; // @[src/main/scala/system/Coherence.scala 74:18 59:23]
  wire  _GEN_37 = 3'h2 == state ? _GEN_7 : _GEN_25; // @[src/main/scala/system/Coherence.scala 74:18]
  wire  _GEN_40 = 3'h1 == state ? io_out_mem_resp_valid : _GEN_28; // @[src/main/scala/system/Coherence.scala 72:14 74:18]
  wire [3:0] _GEN_41 = 3'h1 == state ? io_out_mem_resp_bits_cmd : _GEN_29; // @[src/main/scala/system/Coherence.scala 72:14 74:18]
  wire [63:0] _GEN_42 = 3'h1 == state ? io_out_mem_resp_bits_rdata : _GEN_30; // @[src/main/scala/system/Coherence.scala 72:14 74:18]
  wire [31:0] _GEN_43 = 3'h1 == state ? io_in_req_bits_addr : _GEN_32; // @[src/main/scala/system/Coherence.scala 74:18 59:23]
  wire [3:0] _GEN_45 = 3'h1 == state ? io_in_req_bits_cmd : _GEN_34; // @[src/main/scala/system/Coherence.scala 74:18 59:23]
  wire [63:0] _GEN_47 = 3'h1 == state ? io_in_req_bits_wdata : _GEN_36; // @[src/main/scala/system/Coherence.scala 74:18 59:23]
  wire  _GEN_48 = 3'h1 == state ? _GEN_7 : _GEN_37; // @[src/main/scala/system/Coherence.scala 74:18]
  assign io_in_req_ready = io_in_req_bits_cmd[0] ? io_out_mem_req_ready & _reqLatch_T : _GEN_6; // @[src/main/scala/system/Coherence.scala 64:61 66:19]
  assign io_in_resp_valid = 3'h0 == state ? io_out_mem_resp_valid : _GEN_40; // @[src/main/scala/system/Coherence.scala 72:14 74:18]
  assign io_in_resp_bits_cmd = 3'h0 == state ? io_out_mem_resp_bits_cmd : _GEN_41; // @[src/main/scala/system/Coherence.scala 72:14 74:18]
  assign io_in_resp_bits_rdata = 3'h0 == state ? io_out_mem_resp_bits_rdata : _GEN_42; // @[src/main/scala/system/Coherence.scala 72:14 74:18]
  assign io_out_mem_req_valid = 3'h0 == state ? _GEN_7 : _GEN_48; // @[src/main/scala/system/Coherence.scala 74:18]
  assign io_out_mem_req_bits_addr = 3'h0 == state ? io_in_req_bits_addr : _GEN_43; // @[src/main/scala/system/Coherence.scala 74:18 59:23]
  assign io_out_mem_req_bits_cmd = 3'h0 == state ? io_in_req_bits_cmd : _GEN_45; // @[src/main/scala/system/Coherence.scala 74:18 59:23]
  assign io_out_mem_req_bits_wdata = 3'h0 == state ? io_in_req_bits_wdata : _GEN_47; // @[src/main/scala/system/Coherence.scala 74:18 59:23]
  assign io_out_mem_resp_ready = 1'h1; // @[src/main/scala/system/Coherence.scala 72:14]
  assign io_out_coh_req_valid = io_in_req_bits_cmd[0] ? 1'h0 : _GEN_5; // @[src/main/scala/system/Coherence.scala 63:24 64:61]
  assign io_out_coh_req_bits_addr = io_in_req_bits_addr; // @[src/main/scala/system/Coherence.scala 54:16]
  assign io_out_coh_req_bits_wdata = io_in_req_bits_wdata; // @[src/main/scala/system/Coherence.scala 54:16]
  assign io_out_coh_resp_ready = 1'h1; // @[src/main/scala/system/Coherence.scala 56:18 74:18]
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/system/Coherence.scala 45:22]
      state <= 3'h0; // @[src/main/scala/system/Coherence.scala 45:22]
    end else if (3'h0 == state) begin // @[src/main/scala/system/Coherence.scala 74:18]
      if (_T_21) begin // @[src/main/scala/system/Coherence.scala 76:27]
        if (_T_4) begin // @[src/main/scala/system/Coherence.scala 77:38]
          state <= 3'h1; // @[src/main/scala/system/Coherence.scala 77:46]
        end else begin
          state <= _GEN_10;
        end
      end
    end else if (3'h1 == state) begin // @[src/main/scala/system/Coherence.scala 74:18]
      if (_T_29) begin // @[src/main/scala/system/Coherence.scala 82:35]
        state <= _state_T_2; // @[src/main/scala/system/Coherence.scala 83:15]
      end
    end else if (3'h2 == state) begin // @[src/main/scala/system/Coherence.scala 74:18]
      state <= _GEN_14;
    end else begin
      state <= _GEN_26;
    end
    if (~inflight & _T_4) begin // @[src/main/scala/system/Coherence.scala 52:27]
      reqLatch_addr <= io_in_req_bits_addr; // @[src/main/scala/system/Coherence.scala 52:27]
    end
    if (~inflight & _T_4) begin // @[src/main/scala/system/Coherence.scala 52:27]
      reqLatch_cmd <= io_in_req_bits_cmd; // @[src/main/scala/system/Coherence.scala 52:27]
    end
    if (~inflight & _T_4) begin // @[src/main/scala/system/Coherence.scala 52:27]
      reqLatch_wdata <= io_in_req_bits_wdata; // @[src/main/scala/system/Coherence.scala 52:27]
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~(io_in_req_valid & ~_T_4 & _T_1))) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Coherence.scala:49 assert(!(thisReq.valid && !thisReq.bits.isRead() && !thisReq.bits.isWrite()))\n"
            ); // @[src/main/scala/system/Coherence.scala 49:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~(io_in_req_valid & ~_T_4 & _T_1)) & ~reset) begin
          $fatal; // @[src/main/scala/system/Coherence.scala 49:9]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  reqLatch_addr = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  reqLatch_cmd = _RAND_2[3:0];
  _RAND_3 = {2{`RANDOM}};
  reqLatch_wdata = _RAND_3[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module AXI42SimpleBusConverter(
  input         clock,
  input         reset,
  output        io_in_aw_ready, // @[src/main/scala/bus/simplebus/ToAXI4.scala 27:14]
  input         io_in_aw_valid, // @[src/main/scala/bus/simplebus/ToAXI4.scala 27:14]
  input  [31:0] io_in_aw_bits_addr, // @[src/main/scala/bus/simplebus/ToAXI4.scala 27:14]
  input  [7:0]  io_in_aw_bits_len, // @[src/main/scala/bus/simplebus/ToAXI4.scala 27:14]
  input  [2:0]  io_in_aw_bits_size, // @[src/main/scala/bus/simplebus/ToAXI4.scala 27:14]
  output        io_in_w_ready, // @[src/main/scala/bus/simplebus/ToAXI4.scala 27:14]
  input         io_in_w_valid, // @[src/main/scala/bus/simplebus/ToAXI4.scala 27:14]
  input  [63:0] io_in_w_bits_data, // @[src/main/scala/bus/simplebus/ToAXI4.scala 27:14]
  input  [7:0]  io_in_w_bits_strb, // @[src/main/scala/bus/simplebus/ToAXI4.scala 27:14]
  input         io_in_b_ready, // @[src/main/scala/bus/simplebus/ToAXI4.scala 27:14]
  output        io_in_b_valid, // @[src/main/scala/bus/simplebus/ToAXI4.scala 27:14]
  output        io_in_ar_ready, // @[src/main/scala/bus/simplebus/ToAXI4.scala 27:14]
  input         io_in_ar_valid, // @[src/main/scala/bus/simplebus/ToAXI4.scala 27:14]
  input  [31:0] io_in_ar_bits_addr, // @[src/main/scala/bus/simplebus/ToAXI4.scala 27:14]
  input         io_in_r_ready, // @[src/main/scala/bus/simplebus/ToAXI4.scala 27:14]
  output        io_in_r_valid, // @[src/main/scala/bus/simplebus/ToAXI4.scala 27:14]
  output [63:0] io_in_r_bits_data, // @[src/main/scala/bus/simplebus/ToAXI4.scala 27:14]
  input         io_out_req_ready, // @[src/main/scala/bus/simplebus/ToAXI4.scala 27:14]
  output        io_out_req_valid, // @[src/main/scala/bus/simplebus/ToAXI4.scala 27:14]
  output [31:0] io_out_req_bits_addr, // @[src/main/scala/bus/simplebus/ToAXI4.scala 27:14]
  output [2:0]  io_out_req_bits_size, // @[src/main/scala/bus/simplebus/ToAXI4.scala 27:14]
  output [3:0]  io_out_req_bits_cmd, // @[src/main/scala/bus/simplebus/ToAXI4.scala 27:14]
  output [7:0]  io_out_req_bits_wmask, // @[src/main/scala/bus/simplebus/ToAXI4.scala 27:14]
  output [63:0] io_out_req_bits_wdata, // @[src/main/scala/bus/simplebus/ToAXI4.scala 27:14]
  output        io_out_resp_ready, // @[src/main/scala/bus/simplebus/ToAXI4.scala 27:14]
  input         io_out_resp_valid, // @[src/main/scala/bus/simplebus/ToAXI4.scala 27:14]
  input  [3:0]  io_out_resp_bits_cmd, // @[src/main/scala/bus/simplebus/ToAXI4.scala 27:14]
  input  [63:0] io_out_resp_bits_rdata // @[src/main/scala/bus/simplebus/ToAXI4.scala 27:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  reg [1:0] inflight_type; // @[src/main/scala/bus/simplebus/ToAXI4.scala 40:30]
  wire  _T = inflight_type == 2'h0; // @[src/main/scala/bus/simplebus/ToAXI4.scala 50:19]
  wire  _T_1 = ~_T; // @[src/main/scala/bus/simplebus/ToAXI4.scala 53:5]
  wire  _T_2 = ~_T_1; // @[src/main/scala/bus/simplebus/ToAXI4.scala 64:9]
  wire  _T_3 = ~_T_1 & io_in_ar_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 64:23]
  wire  _T_4 = io_out_req_ready & io_out_req_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  wire [1:0] _GEN_1 = _T_4 ? 2'h1 : inflight_type; // @[src/main/scala/bus/simplebus/ToAXI4.scala 43:19 74:25 40:30]
  wire [31:0] _GEN_2 = ~_T_1 & io_in_ar_valid ? io_in_ar_bits_addr : 32'h0; // @[src/main/scala/bus/simplebus/ToAXI4.scala 64:40 66:14 59:7]
  wire [2:0] _GEN_4 = ~_T_1 & io_in_ar_valid ? 3'h2 : 3'h0; // @[src/main/scala/bus/simplebus/ToAXI4.scala 64:40 69:14 59:7]
  wire [1:0] _GEN_8 = ~_T_1 & io_in_ar_valid ? _GEN_1 : inflight_type; // @[src/main/scala/bus/simplebus/ToAXI4.scala 40:30 64:40]
  wire  _T_5 = inflight_type == 2'h1; // @[src/main/scala/bus/simplebus/ToAXI4.scala 50:19]
  wire  _io_in_r_bits_last_T = io_out_resp_bits_cmd == 4'h6; // @[src/main/scala/bus/simplebus/SimpleBus.scala 91:24]
  wire  _T_7 = io_in_r_ready & io_in_r_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  wire [1:0] _GEN_9 = _T_7 & _io_in_r_bits_last_T ? 2'h0 : _GEN_8; // @[src/main/scala/bus/simplebus/ToAXI4.scala 46:19 88:42]
  wire [1:0] _GEN_15 = _T_5 & io_out_resp_valid ? _GEN_9 : _GEN_8; // @[src/main/scala/bus/simplebus/ToAXI4.scala 79:46]
  reg [31:0] aw_reg_addr; // @[src/main/scala/bus/simplebus/ToAXI4.scala 94:19]
  reg [7:0] aw_reg_len; // @[src/main/scala/bus/simplebus/ToAXI4.scala 94:19]
  reg [2:0] aw_reg_size; // @[src/main/scala/bus/simplebus/ToAXI4.scala 94:19]
  reg  bresp_en; // @[src/main/scala/bus/simplebus/ToAXI4.scala 95:25]
  wire  _T_14 = ~io_in_ar_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 97:42]
  wire  _T_16 = io_in_aw_ready & io_in_aw_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  wire  _T_17 = inflight_type == 2'h2; // @[src/main/scala/bus/simplebus/ToAXI4.scala 50:19]
  wire  _T_18 = io_in_w_ready & io_in_w_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  wire [2:0] _io_out_req_bits_cmd_T_4 = aw_reg_len == 8'h0 ? 3'h1 : 3'h7; // @[src/main/scala/bus/simplebus/ToAXI4.scala 107:19]
  wire  _GEN_37 = _T_17 & _T_18 | bresp_en; // @[src/main/scala/bus/simplebus/ToAXI4.scala 105:43 95:25]
  wire  _T_20 = io_in_b_ready & io_in_b_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  wire  _T_21 = io_in_ar_ready & io_in_ar_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  wire  _T_28 = ~reset; // @[src/main/scala/bus/simplebus/ToAXI4.scala 137:30]
  wire  _T_45 = io_out_resp_ready & io_out_resp_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  assign io_in_aw_ready = _T_2 & _T_14; // @[src/main/scala/bus/simplebus/ToAXI4.scala 132:33]
  assign io_in_w_ready = _T_17 & io_out_req_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 133:38]
  assign io_in_b_valid = bresp_en & io_out_resp_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 134:27]
  assign io_in_ar_ready = _T_2 & io_out_req_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 129:33]
  assign io_in_r_valid = _T_5 & io_out_resp_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 130:36]
  assign io_in_r_bits_data = _T_5 & io_out_resp_valid ? io_out_resp_bits_rdata : 64'h0; // @[src/main/scala/bus/simplebus/ToAXI4.scala 79:46 81:12 60:5]
  assign io_out_req_valid = _T_3 | _T_17 & io_in_w_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 127:52]
  assign io_out_req_bits_addr = _T_17 & _T_18 ? aw_reg_addr : _GEN_2; // @[src/main/scala/bus/simplebus/ToAXI4.scala 105:43 109:14]
  assign io_out_req_bits_size = _T_17 & _T_18 ? aw_reg_size : _GEN_4; // @[src/main/scala/bus/simplebus/ToAXI4.scala 105:43 110:14]
  assign io_out_req_bits_cmd = _T_17 & _T_18 ? {{1'd0}, _io_out_req_bits_cmd_T_4} : 4'h0; // @[src/main/scala/bus/simplebus/ToAXI4.scala 105:43 107:13]
  assign io_out_req_bits_wmask = _T_17 & _T_18 ? io_in_w_bits_strb : 8'h0; // @[src/main/scala/bus/simplebus/ToAXI4.scala 105:43 111:15]
  assign io_out_req_bits_wdata = _T_17 & _T_18 ? io_in_w_bits_data : 64'h0; // @[src/main/scala/bus/simplebus/ToAXI4.scala 105:43 112:15]
  assign io_out_resp_ready = _T_2 | _T_5 & io_in_r_ready | _T_17 & io_in_b_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 128:73]
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/bus/simplebus/ToAXI4.scala 40:30]
      inflight_type <= 2'h0; // @[src/main/scala/bus/simplebus/ToAXI4.scala 40:30]
    end else if (_T_20) begin // @[src/main/scala/bus/simplebus/ToAXI4.scala 120:21]
      inflight_type <= 2'h0; // @[src/main/scala/bus/simplebus/ToAXI4.scala 46:19]
    end else if (_T_2 & io_in_aw_valid & ~io_in_ar_valid) begin // @[src/main/scala/bus/simplebus/ToAXI4.scala 97:57]
      if (_T_16) begin // @[src/main/scala/bus/simplebus/ToAXI4.scala 100:24]
        inflight_type <= 2'h2; // @[src/main/scala/bus/simplebus/ToAXI4.scala 43:19]
      end else begin
        inflight_type <= _GEN_15;
      end
    end else begin
      inflight_type <= _GEN_15;
    end
    if (_T_2 & io_in_aw_valid & ~io_in_ar_valid) begin // @[src/main/scala/bus/simplebus/ToAXI4.scala 97:57]
      aw_reg_addr <= io_in_aw_bits_addr; // @[src/main/scala/bus/simplebus/ToAXI4.scala 98:12]
    end
    if (_T_2 & io_in_aw_valid & ~io_in_ar_valid) begin // @[src/main/scala/bus/simplebus/ToAXI4.scala 97:57]
      aw_reg_len <= io_in_aw_bits_len; // @[src/main/scala/bus/simplebus/ToAXI4.scala 98:12]
    end
    if (_T_2 & io_in_aw_valid & ~io_in_ar_valid) begin // @[src/main/scala/bus/simplebus/ToAXI4.scala 97:57]
      aw_reg_size <= io_in_aw_bits_size; // @[src/main/scala/bus/simplebus/ToAXI4.scala 98:12]
    end
    if (reset) begin // @[src/main/scala/bus/simplebus/ToAXI4.scala 95:25]
      bresp_en <= 1'h0; // @[src/main/scala/bus/simplebus/ToAXI4.scala 95:25]
    end else if (_T_20) begin // @[src/main/scala/bus/simplebus/ToAXI4.scala 120:21]
      bresp_en <= 1'h0; // @[src/main/scala/bus/simplebus/ToAXI4.scala 121:14]
    end else begin
      bresp_en <= _GEN_37;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_21 & ~reset & ~(_T_4 & _T_2)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:137 when (axi.ar.fire) { assert(mem.req.fire && !isInflight()); }\n"
            ); // @[src/main/scala/bus/simplebus/ToAXI4.scala 137:30]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(_T_4 & _T_2) & (_T_21 & ~reset)) begin
          $fatal; // @[src/main/scala/bus/simplebus/ToAXI4.scala 137:30]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_16 & _T_28 & ~_T_2) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:138 when (axi.aw.fire) { assert(!isInflight()); }\n"); // @[src/main/scala/bus/simplebus/ToAXI4.scala 138:30]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~_T_2 & (_T_16 & _T_28)) begin
          $fatal; // @[src/main/scala/bus/simplebus/ToAXI4.scala 138:30]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_18 & _T_28 & ~(_T_4 & _T_17)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:139 when (axi.w.fire) { assert(mem.req .fire && isState(axi_write)); }\n"
            ); // @[src/main/scala/bus/simplebus/ToAXI4.scala 139:29]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(_T_4 & _T_17) & (_T_18 & _T_28)) begin
          $fatal; // @[src/main/scala/bus/simplebus/ToAXI4.scala 139:29]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_20 & _T_28 & ~(_T_45 & _T_17)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:140 when (axi.b.fire) { assert(mem.resp.fire && isState(axi_write)); }\n"
            ); // @[src/main/scala/bus/simplebus/ToAXI4.scala 140:29]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(_T_45 & _T_17) & (_T_20 & _T_28)) begin
          $fatal; // @[src/main/scala/bus/simplebus/ToAXI4.scala 140:29]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_7 & _T_28 & ~(_T_45 & _T_5)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:141 when (axi.r.fire) { assert(mem.resp.fire && isState(axi_read)); }\n"
            ); // @[src/main/scala/bus/simplebus/ToAXI4.scala 141:29]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(_T_45 & _T_5) & (_T_7 & _T_28)) begin
          $fatal; // @[src/main/scala/bus/simplebus/ToAXI4.scala 141:29]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  inflight_type = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  aw_reg_addr = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  aw_reg_len = _RAND_2[7:0];
  _RAND_3 = {1{`RANDOM}};
  aw_reg_size = _RAND_3[2:0];
  _RAND_4 = {1{`RANDOM}};
  bresp_en = _RAND_4[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Prefetcher(
  input         clock,
  input         reset,
  output        io_in_ready, // @[src/main/scala/system/Prefetcher.scala 33:20]
  input         io_in_valid, // @[src/main/scala/system/Prefetcher.scala 33:20]
  input  [31:0] io_in_bits_addr, // @[src/main/scala/system/Prefetcher.scala 33:20]
  input  [2:0]  io_in_bits_size, // @[src/main/scala/system/Prefetcher.scala 33:20]
  input  [3:0]  io_in_bits_cmd, // @[src/main/scala/system/Prefetcher.scala 33:20]
  input  [7:0]  io_in_bits_wmask, // @[src/main/scala/system/Prefetcher.scala 33:20]
  input  [63:0] io_in_bits_wdata, // @[src/main/scala/system/Prefetcher.scala 33:20]
  input         io_out_ready, // @[src/main/scala/system/Prefetcher.scala 33:20]
  output        io_out_valid, // @[src/main/scala/system/Prefetcher.scala 33:20]
  output [31:0] io_out_bits_addr, // @[src/main/scala/system/Prefetcher.scala 33:20]
  output [2:0]  io_out_bits_size, // @[src/main/scala/system/Prefetcher.scala 33:20]
  output [3:0]  io_out_bits_cmd, // @[src/main/scala/system/Prefetcher.scala 33:20]
  output [7:0]  io_out_bits_wmask, // @[src/main/scala/system/Prefetcher.scala 33:20]
  output [63:0] io_out_bits_wdata, // @[src/main/scala/system/Prefetcher.scala 33:20]
  input         DISPLAY_ENABLE
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
`endif // RANDOMIZE_REG_INIT
  reg  getNewReq; // @[src/main/scala/system/Prefetcher.scala 37:26]
  reg [31:0] prefetchReq_addr; // @[src/main/scala/system/Prefetcher.scala 38:28]
  reg [2:0] prefetchReq_size; // @[src/main/scala/system/Prefetcher.scala 38:28]
  reg [7:0] prefetchReq_wmask; // @[src/main/scala/system/Prefetcher.scala 38:28]
  reg [63:0] prefetchReq_wdata; // @[src/main/scala/system/Prefetcher.scala 38:28]
  reg [63:0] lastReqAddr; // @[src/main/scala/system/Prefetcher.scala 44:28]
  wire  _T = io_in_ready & io_in_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  wire [63:0] _GEN_9 = {{32'd0}, io_in_bits_addr}; // @[src/main/scala/system/Prefetcher.scala 50:30]
  wire [63:0] _neqAddr_T = _GEN_9 & 64'hffffffffffffffc0; // @[src/main/scala/system/Prefetcher.scala 50:30]
  wire [63:0] _neqAddr_T_1 = lastReqAddr & 64'hffffffffffffffc0; // @[src/main/scala/system/Prefetcher.scala 50:59]
  wire  neqAddr = _neqAddr_T != _neqAddr_T_1; // @[src/main/scala/system/Prefetcher.scala 50:42]
  wire  _io_in_ready_T_1 = io_out_ready & io_out_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  wire [31:0] _io_out_valid_T = prefetchReq_addr ^ 32'h30000000; // @[src/main/scala/nutcore/NutCore.scala 87:11]
  wire  _io_out_valid_T_2 = _io_out_valid_T[31:28] == 4'h0; // @[src/main/scala/nutcore/NutCore.scala 87:44]
  wire [31:0] _io_out_valid_T_3 = prefetchReq_addr ^ 32'h40000000; // @[src/main/scala/nutcore/NutCore.scala 87:11]
  wire  _io_out_valid_T_5 = _io_out_valid_T_3[31:30] == 2'h0; // @[src/main/scala/nutcore/NutCore.scala 87:44]
  wire  _io_out_valid_T_6 = _io_out_valid_T_2 | _io_out_valid_T_5; // @[src/main/scala/nutcore/NutCore.scala 88:15]
  reg [63:0] c; // @[src/main/scala/utils/GTimer.scala 24:20]
  wire [63:0] _c_T_1 = c + 64'h1; // @[src/main/scala/utils/GTimer.scala 25:12]
  assign io_in_ready = ~getNewReq & (~io_in_valid | _io_in_ready_T_1); // @[src/main/scala/system/Prefetcher.scala 52:21 55:17 60:17]
  assign io_out_valid = ~getNewReq ? io_in_valid : ~_io_out_valid_T_6; // @[src/main/scala/system/Prefetcher.scala 52:21 54:18 59:18]
  assign io_out_bits_addr = ~getNewReq ? io_in_bits_addr : prefetchReq_addr; // @[src/main/scala/system/Prefetcher.scala 52:21 53:17 58:17]
  assign io_out_bits_size = ~getNewReq ? io_in_bits_size : prefetchReq_size; // @[src/main/scala/system/Prefetcher.scala 52:21 53:17 58:17]
  assign io_out_bits_cmd = ~getNewReq ? io_in_bits_cmd : 4'h4; // @[src/main/scala/system/Prefetcher.scala 52:21 53:17 58:17]
  assign io_out_bits_wmask = ~getNewReq ? io_in_bits_wmask : prefetchReq_wmask; // @[src/main/scala/system/Prefetcher.scala 52:21 53:17 58:17]
  assign io_out_bits_wdata = ~getNewReq ? io_in_bits_wdata : prefetchReq_wdata; // @[src/main/scala/system/Prefetcher.scala 52:21 53:17 58:17]
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/system/Prefetcher.scala 37:26]
      getNewReq <= 1'h0; // @[src/main/scala/system/Prefetcher.scala 37:26]
    end else if (~getNewReq) begin // @[src/main/scala/system/Prefetcher.scala 52:21]
      getNewReq <= _T & io_in_bits_cmd[1] & neqAddr; // @[src/main/scala/system/Prefetcher.scala 56:15]
    end else begin
      getNewReq <= ~(_io_in_ready_T_1 | _io_out_valid_T_6); // @[src/main/scala/system/Prefetcher.scala 61:15]
    end
    prefetchReq_addr <= io_in_bits_addr + 32'h40; // @[src/main/scala/system/Prefetcher.scala 40:39]
    prefetchReq_size <= io_in_bits_size; // @[src/main/scala/system/Prefetcher.scala 38:28]
    prefetchReq_wmask <= io_in_bits_wmask; // @[src/main/scala/system/Prefetcher.scala 38:28]
    prefetchReq_wdata <= io_in_bits_wdata; // @[src/main/scala/system/Prefetcher.scala 38:28]
    if (reset) begin // @[src/main/scala/system/Prefetcher.scala 44:28]
      lastReqAddr <= 64'h0; // @[src/main/scala/system/Prefetcher.scala 44:28]
    end else if (_T) begin // @[src/main/scala/system/Prefetcher.scala 45:21]
      lastReqAddr <= {{32'd0}, io_in_bits_addr}; // @[src/main/scala/system/Prefetcher.scala 46:18]
    end
    if (reset) begin // @[src/main/scala/utils/GTimer.scala 24:20]
      c <= 64'h0; // @[src/main/scala/utils/GTimer.scala 24:20]
    end else begin
      c <= _c_T_1; // @[src/main/scala/utils/GTimer.scala 25:7]
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & ~reset) begin
          $fwrite(32'h80000002,"%d: [Prefetcher]: in(%d,%d), out(%d,%d), in.bits.addr = %x\n",c,io_in_valid,io_in_ready,
            io_out_valid,io_out_ready,io_in_bits_addr); // @[src/main/scala/system/Prefetcher.scala 65:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  getNewReq = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  prefetchReq_addr = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  prefetchReq_size = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  prefetchReq_wmask = _RAND_3[7:0];
  _RAND_4 = {2{`RANDOM}};
  prefetchReq_wdata = _RAND_4[63:0];
  _RAND_5 = {2{`RANDOM}};
  lastReqAddr = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  c = _RAND_6[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module CacheStage1_2(
  input         clock,
  input         reset,
  output        io_in_ready, // @[src/main/scala/nutcore/mem/Cache.scala 133:14]
  input         io_in_valid, // @[src/main/scala/nutcore/mem/Cache.scala 133:14]
  input  [31:0] io_in_bits_addr, // @[src/main/scala/nutcore/mem/Cache.scala 133:14]
  input  [2:0]  io_in_bits_size, // @[src/main/scala/nutcore/mem/Cache.scala 133:14]
  input  [3:0]  io_in_bits_cmd, // @[src/main/scala/nutcore/mem/Cache.scala 133:14]
  input  [7:0]  io_in_bits_wmask, // @[src/main/scala/nutcore/mem/Cache.scala 133:14]
  input  [63:0] io_in_bits_wdata, // @[src/main/scala/nutcore/mem/Cache.scala 133:14]
  input         io_out_ready, // @[src/main/scala/nutcore/mem/Cache.scala 133:14]
  output        io_out_valid, // @[src/main/scala/nutcore/mem/Cache.scala 133:14]
  output [31:0] io_out_bits_req_addr, // @[src/main/scala/nutcore/mem/Cache.scala 133:14]
  output [2:0]  io_out_bits_req_size, // @[src/main/scala/nutcore/mem/Cache.scala 133:14]
  output [3:0]  io_out_bits_req_cmd, // @[src/main/scala/nutcore/mem/Cache.scala 133:14]
  output [7:0]  io_out_bits_req_wmask, // @[src/main/scala/nutcore/mem/Cache.scala 133:14]
  output [63:0] io_out_bits_req_wdata, // @[src/main/scala/nutcore/mem/Cache.scala 133:14]
  input         io_metaReadBus_req_ready, // @[src/main/scala/nutcore/mem/Cache.scala 133:14]
  output        io_metaReadBus_req_valid, // @[src/main/scala/nutcore/mem/Cache.scala 133:14]
  output [8:0]  io_metaReadBus_req_bits_setIdx, // @[src/main/scala/nutcore/mem/Cache.scala 133:14]
  input  [16:0] io_metaReadBus_resp_data_0_tag, // @[src/main/scala/nutcore/mem/Cache.scala 133:14]
  input         io_metaReadBus_resp_data_0_valid, // @[src/main/scala/nutcore/mem/Cache.scala 133:14]
  input         io_metaReadBus_resp_data_0_dirty, // @[src/main/scala/nutcore/mem/Cache.scala 133:14]
  input  [16:0] io_metaReadBus_resp_data_1_tag, // @[src/main/scala/nutcore/mem/Cache.scala 133:14]
  input         io_metaReadBus_resp_data_1_valid, // @[src/main/scala/nutcore/mem/Cache.scala 133:14]
  input         io_metaReadBus_resp_data_1_dirty, // @[src/main/scala/nutcore/mem/Cache.scala 133:14]
  input  [16:0] io_metaReadBus_resp_data_2_tag, // @[src/main/scala/nutcore/mem/Cache.scala 133:14]
  input         io_metaReadBus_resp_data_2_valid, // @[src/main/scala/nutcore/mem/Cache.scala 133:14]
  input         io_metaReadBus_resp_data_2_dirty, // @[src/main/scala/nutcore/mem/Cache.scala 133:14]
  input  [16:0] io_metaReadBus_resp_data_3_tag, // @[src/main/scala/nutcore/mem/Cache.scala 133:14]
  input         io_metaReadBus_resp_data_3_valid, // @[src/main/scala/nutcore/mem/Cache.scala 133:14]
  input         io_metaReadBus_resp_data_3_dirty, // @[src/main/scala/nutcore/mem/Cache.scala 133:14]
  input         io_dataReadBus_req_ready, // @[src/main/scala/nutcore/mem/Cache.scala 133:14]
  output        io_dataReadBus_req_valid, // @[src/main/scala/nutcore/mem/Cache.scala 133:14]
  output [11:0] io_dataReadBus_req_bits_setIdx, // @[src/main/scala/nutcore/mem/Cache.scala 133:14]
  input  [63:0] io_dataReadBus_resp_data_0_data, // @[src/main/scala/nutcore/mem/Cache.scala 133:14]
  input  [63:0] io_dataReadBus_resp_data_1_data, // @[src/main/scala/nutcore/mem/Cache.scala 133:14]
  input  [63:0] io_dataReadBus_resp_data_2_data, // @[src/main/scala/nutcore/mem/Cache.scala 133:14]
  input  [63:0] io_dataReadBus_resp_data_3_data, // @[src/main/scala/nutcore/mem/Cache.scala 133:14]
  input         DISPLAY_ENABLE
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  wire  _T = io_in_ready & io_in_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  reg [63:0] c; // @[src/main/scala/utils/GTimer.scala 24:20]
  wire [63:0] _c_T_1 = c + 64'h1; // @[src/main/scala/utils/GTimer.scala 25:12]
  wire  _T_1 = _T & DISPLAY_ENABLE; // @[src/main/scala/utils/Debug.scala 55:16]
  wire  _T_3 = ~reset; // @[src/main/scala/utils/Debug.scala 56:24]
  wire  _io_in_ready_T_1 = io_out_ready & io_out_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  reg [63:0] c_1; // @[src/main/scala/utils/GTimer.scala 24:20]
  wire [63:0] _c_T_3 = c_1 + 64'h1; // @[src/main/scala/utils/GTimer.scala 25:12]
  assign io_in_ready = (~io_in_valid | _io_in_ready_T_1) & io_metaReadBus_req_ready & io_dataReadBus_req_ready; // @[src/main/scala/nutcore/mem/Cache.scala 145:76]
  assign io_out_valid = io_in_valid & io_metaReadBus_req_ready & io_dataReadBus_req_ready; // @[src/main/scala/nutcore/mem/Cache.scala 144:59]
  assign io_out_bits_req_addr = io_in_bits_addr; // @[src/main/scala/nutcore/mem/Cache.scala 143:19]
  assign io_out_bits_req_size = io_in_bits_size; // @[src/main/scala/nutcore/mem/Cache.scala 143:19]
  assign io_out_bits_req_cmd = io_in_bits_cmd; // @[src/main/scala/nutcore/mem/Cache.scala 143:19]
  assign io_out_bits_req_wmask = io_in_bits_wmask; // @[src/main/scala/nutcore/mem/Cache.scala 143:19]
  assign io_out_bits_req_wdata = io_in_bits_wdata; // @[src/main/scala/nutcore/mem/Cache.scala 143:19]
  assign io_metaReadBus_req_valid = io_in_valid & io_out_ready; // @[src/main/scala/nutcore/mem/Cache.scala 139:34]
  assign io_metaReadBus_req_bits_setIdx = io_in_bits_addr[14:6]; // @[src/main/scala/nutcore/mem/Cache.scala 77:45]
  assign io_dataReadBus_req_valid = io_in_valid & io_out_ready; // @[src/main/scala/nutcore/mem/Cache.scala 139:34]
  assign io_dataReadBus_req_bits_setIdx = {io_in_bits_addr[14:6],io_in_bits_addr[5:3]}; // @[src/main/scala/nutcore/mem/Cache.scala 78:35]
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/utils/GTimer.scala 24:20]
      c <= 64'h0; // @[src/main/scala/utils/GTimer.scala 24:20]
    end else begin
      c <= _c_T_1; // @[src/main/scala/utils/GTimer.scala 25:7]
    end
    if (reset) begin // @[src/main/scala/utils/GTimer.scala 24:20]
      c_1 <= 64'h0; // @[src/main/scala/utils/GTimer.scala 24:20]
    end else begin
      c_1 <= _c_T_3; // @[src/main/scala/utils/GTimer.scala 25:7]
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1 & ~reset) begin
          $fwrite(32'h80000002,"[%d] CacheStage1_2: ",c); // @[src/main/scala/utils/Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1 & _T_3) begin
          $fwrite(32'h80000002,"[L1$] cache stage1, addr in: %x, user: %x id: %x\n",io_in_bits_addr,1'h0,1'h0); // @[src/main/scala/utils/Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & ~reset) begin
          $fwrite(32'h80000002,"[%d] CacheStage1_2: ",c_1); // @[src/main/scala/utils/Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_3) begin
          $fwrite(32'h80000002,
            "in.ready = %d, in.valid = %d, out.valid = %d, out.ready = %d, addr = %x, cmd = %x, dataReadBus.req.valid = %d\n"
            ,io_in_ready,io_in_valid,io_out_valid,io_out_ready,io_in_bits_addr,io_in_bits_cmd,io_dataReadBus_req_valid); // @[src/main/scala/utils/Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  c = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  c_1 = _RAND_1[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module CacheStage2_2(
  input         clock,
  input         reset,
  output        io_in_ready, // @[src/main/scala/nutcore/mem/Cache.scala 171:14]
  input         io_in_valid, // @[src/main/scala/nutcore/mem/Cache.scala 171:14]
  input  [31:0] io_in_bits_req_addr, // @[src/main/scala/nutcore/mem/Cache.scala 171:14]
  input  [2:0]  io_in_bits_req_size, // @[src/main/scala/nutcore/mem/Cache.scala 171:14]
  input  [3:0]  io_in_bits_req_cmd, // @[src/main/scala/nutcore/mem/Cache.scala 171:14]
  input  [7:0]  io_in_bits_req_wmask, // @[src/main/scala/nutcore/mem/Cache.scala 171:14]
  input  [63:0] io_in_bits_req_wdata, // @[src/main/scala/nutcore/mem/Cache.scala 171:14]
  input         io_out_ready, // @[src/main/scala/nutcore/mem/Cache.scala 171:14]
  output        io_out_valid, // @[src/main/scala/nutcore/mem/Cache.scala 171:14]
  output [31:0] io_out_bits_req_addr, // @[src/main/scala/nutcore/mem/Cache.scala 171:14]
  output [2:0]  io_out_bits_req_size, // @[src/main/scala/nutcore/mem/Cache.scala 171:14]
  output [3:0]  io_out_bits_req_cmd, // @[src/main/scala/nutcore/mem/Cache.scala 171:14]
  output [7:0]  io_out_bits_req_wmask, // @[src/main/scala/nutcore/mem/Cache.scala 171:14]
  output [63:0] io_out_bits_req_wdata, // @[src/main/scala/nutcore/mem/Cache.scala 171:14]
  output [16:0] io_out_bits_metas_0_tag, // @[src/main/scala/nutcore/mem/Cache.scala 171:14]
  output        io_out_bits_metas_0_valid, // @[src/main/scala/nutcore/mem/Cache.scala 171:14]
  output        io_out_bits_metas_0_dirty, // @[src/main/scala/nutcore/mem/Cache.scala 171:14]
  output [16:0] io_out_bits_metas_1_tag, // @[src/main/scala/nutcore/mem/Cache.scala 171:14]
  output        io_out_bits_metas_1_valid, // @[src/main/scala/nutcore/mem/Cache.scala 171:14]
  output        io_out_bits_metas_1_dirty, // @[src/main/scala/nutcore/mem/Cache.scala 171:14]
  output [16:0] io_out_bits_metas_2_tag, // @[src/main/scala/nutcore/mem/Cache.scala 171:14]
  output        io_out_bits_metas_2_valid, // @[src/main/scala/nutcore/mem/Cache.scala 171:14]
  output        io_out_bits_metas_2_dirty, // @[src/main/scala/nutcore/mem/Cache.scala 171:14]
  output [16:0] io_out_bits_metas_3_tag, // @[src/main/scala/nutcore/mem/Cache.scala 171:14]
  output        io_out_bits_metas_3_valid, // @[src/main/scala/nutcore/mem/Cache.scala 171:14]
  output        io_out_bits_metas_3_dirty, // @[src/main/scala/nutcore/mem/Cache.scala 171:14]
  output [63:0] io_out_bits_datas_0_data, // @[src/main/scala/nutcore/mem/Cache.scala 171:14]
  output [63:0] io_out_bits_datas_1_data, // @[src/main/scala/nutcore/mem/Cache.scala 171:14]
  output [63:0] io_out_bits_datas_2_data, // @[src/main/scala/nutcore/mem/Cache.scala 171:14]
  output [63:0] io_out_bits_datas_3_data, // @[src/main/scala/nutcore/mem/Cache.scala 171:14]
  output        io_out_bits_hit, // @[src/main/scala/nutcore/mem/Cache.scala 171:14]
  output [3:0]  io_out_bits_waymask, // @[src/main/scala/nutcore/mem/Cache.scala 171:14]
  output        io_out_bits_mmio, // @[src/main/scala/nutcore/mem/Cache.scala 171:14]
  output        io_out_bits_isForwardData, // @[src/main/scala/nutcore/mem/Cache.scala 171:14]
  output [63:0] io_out_bits_forwardData_data_data, // @[src/main/scala/nutcore/mem/Cache.scala 171:14]
  output [3:0]  io_out_bits_forwardData_waymask, // @[src/main/scala/nutcore/mem/Cache.scala 171:14]
  input  [16:0] io_metaReadResp_0_tag, // @[src/main/scala/nutcore/mem/Cache.scala 171:14]
  input         io_metaReadResp_0_valid, // @[src/main/scala/nutcore/mem/Cache.scala 171:14]
  input         io_metaReadResp_0_dirty, // @[src/main/scala/nutcore/mem/Cache.scala 171:14]
  input  [16:0] io_metaReadResp_1_tag, // @[src/main/scala/nutcore/mem/Cache.scala 171:14]
  input         io_metaReadResp_1_valid, // @[src/main/scala/nutcore/mem/Cache.scala 171:14]
  input         io_metaReadResp_1_dirty, // @[src/main/scala/nutcore/mem/Cache.scala 171:14]
  input  [16:0] io_metaReadResp_2_tag, // @[src/main/scala/nutcore/mem/Cache.scala 171:14]
  input         io_metaReadResp_2_valid, // @[src/main/scala/nutcore/mem/Cache.scala 171:14]
  input         io_metaReadResp_2_dirty, // @[src/main/scala/nutcore/mem/Cache.scala 171:14]
  input  [16:0] io_metaReadResp_3_tag, // @[src/main/scala/nutcore/mem/Cache.scala 171:14]
  input         io_metaReadResp_3_valid, // @[src/main/scala/nutcore/mem/Cache.scala 171:14]
  input         io_metaReadResp_3_dirty, // @[src/main/scala/nutcore/mem/Cache.scala 171:14]
  input  [63:0] io_dataReadResp_0_data, // @[src/main/scala/nutcore/mem/Cache.scala 171:14]
  input  [63:0] io_dataReadResp_1_data, // @[src/main/scala/nutcore/mem/Cache.scala 171:14]
  input  [63:0] io_dataReadResp_2_data, // @[src/main/scala/nutcore/mem/Cache.scala 171:14]
  input  [63:0] io_dataReadResp_3_data, // @[src/main/scala/nutcore/mem/Cache.scala 171:14]
  input         io_metaWriteBus_req_valid, // @[src/main/scala/nutcore/mem/Cache.scala 171:14]
  input  [8:0]  io_metaWriteBus_req_bits_setIdx, // @[src/main/scala/nutcore/mem/Cache.scala 171:14]
  input  [16:0] io_metaWriteBus_req_bits_data_tag, // @[src/main/scala/nutcore/mem/Cache.scala 171:14]
  input         io_metaWriteBus_req_bits_data_dirty, // @[src/main/scala/nutcore/mem/Cache.scala 171:14]
  input  [3:0]  io_metaWriteBus_req_bits_waymask, // @[src/main/scala/nutcore/mem/Cache.scala 171:14]
  input         io_dataWriteBus_req_valid, // @[src/main/scala/nutcore/mem/Cache.scala 171:14]
  input  [11:0] io_dataWriteBus_req_bits_setIdx, // @[src/main/scala/nutcore/mem/Cache.scala 171:14]
  input  [63:0] io_dataWriteBus_req_bits_data_data, // @[src/main/scala/nutcore/mem/Cache.scala 171:14]
  input  [3:0]  io_dataWriteBus_req_bits_waymask, // @[src/main/scala/nutcore/mem/Cache.scala 171:14]
  input         DISPLAY_ENABLE
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [63:0] _RAND_12;
  reg [63:0] _RAND_13;
  reg [63:0] _RAND_14;
  reg [63:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [63:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [63:0] _RAND_19;
  reg [63:0] _RAND_20;
`endif // RANDOMIZE_REG_INIT
  wire [2:0] addr_wordIndex = io_in_bits_req_addr[5:3]; // @[src/main/scala/nutcore/mem/Cache.scala 174:31]
  wire [8:0] addr_index = io_in_bits_req_addr[14:6]; // @[src/main/scala/nutcore/mem/Cache.scala 174:31]
  wire [16:0] addr_tag = io_in_bits_req_addr[31:15]; // @[src/main/scala/nutcore/mem/Cache.scala 174:31]
  wire  isForwardMeta = io_in_valid & io_metaWriteBus_req_valid & io_metaWriteBus_req_bits_setIdx == addr_index; // @[src/main/scala/nutcore/mem/Cache.scala 176:64]
  reg  isForwardMetaReg; // @[src/main/scala/nutcore/mem/Cache.scala 177:33]
  wire  _GEN_0 = isForwardMeta | isForwardMetaReg; // @[src/main/scala/nutcore/mem/Cache.scala 178:24 177:33 178:43]
  wire  _T = io_in_ready & io_in_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  wire  _T_1 = ~io_in_valid; // @[src/main/scala/nutcore/mem/Cache.scala 179:23]
  wire  _T_2 = _T | ~io_in_valid; // @[src/main/scala/nutcore/mem/Cache.scala 179:20]
  reg [16:0] forwardMetaReg_data_tag; // @[src/main/scala/nutcore/mem/Cache.scala 180:33]
  reg  forwardMetaReg_data_dirty; // @[src/main/scala/nutcore/mem/Cache.scala 180:33]
  reg [3:0] forwardMetaReg_waymask; // @[src/main/scala/nutcore/mem/Cache.scala 180:33]
  wire [16:0] _GEN_3 = isForwardMeta ? io_metaWriteBus_req_bits_data_tag : forwardMetaReg_data_tag; // @[src/main/scala/nutcore/mem/Cache.scala 180:{33,33,33}]
  wire  _GEN_5 = isForwardMeta ? io_metaWriteBus_req_bits_data_dirty : forwardMetaReg_data_dirty; // @[src/main/scala/nutcore/mem/Cache.scala 180:{33,33,33}]
  wire [3:0] _GEN_6 = isForwardMeta ? io_metaWriteBus_req_bits_waymask : forwardMetaReg_waymask; // @[src/main/scala/nutcore/mem/Cache.scala 180:{33,33,33}]
  wire  pickForwardMeta = isForwardMetaReg | isForwardMeta; // @[src/main/scala/nutcore/mem/Cache.scala 183:42]
  wire  forwardWaymask_0 = _GEN_6[0]; // @[src/main/scala/nutcore/mem/Cache.scala 185:61]
  wire  forwardWaymask_1 = _GEN_6[1]; // @[src/main/scala/nutcore/mem/Cache.scala 185:61]
  wire  forwardWaymask_2 = _GEN_6[2]; // @[src/main/scala/nutcore/mem/Cache.scala 185:61]
  wire  forwardWaymask_3 = _GEN_6[3]; // @[src/main/scala/nutcore/mem/Cache.scala 185:61]
  wire [16:0] metaWay_0_tag = pickForwardMeta & forwardWaymask_0 ? _GEN_3 : io_metaReadResp_0_tag; // @[src/main/scala/nutcore/mem/Cache.scala 187:22]
  wire  metaWay_0_valid = pickForwardMeta & forwardWaymask_0 | io_metaReadResp_0_valid; // @[src/main/scala/nutcore/mem/Cache.scala 187:22]
  wire [16:0] metaWay_1_tag = pickForwardMeta & forwardWaymask_1 ? _GEN_3 : io_metaReadResp_1_tag; // @[src/main/scala/nutcore/mem/Cache.scala 187:22]
  wire  metaWay_1_valid = pickForwardMeta & forwardWaymask_1 | io_metaReadResp_1_valid; // @[src/main/scala/nutcore/mem/Cache.scala 187:22]
  wire [16:0] metaWay_2_tag = pickForwardMeta & forwardWaymask_2 ? _GEN_3 : io_metaReadResp_2_tag; // @[src/main/scala/nutcore/mem/Cache.scala 187:22]
  wire  metaWay_2_valid = pickForwardMeta & forwardWaymask_2 | io_metaReadResp_2_valid; // @[src/main/scala/nutcore/mem/Cache.scala 187:22]
  wire [16:0] metaWay_3_tag = pickForwardMeta & forwardWaymask_3 ? _GEN_3 : io_metaReadResp_3_tag; // @[src/main/scala/nutcore/mem/Cache.scala 187:22]
  wire  metaWay_3_valid = pickForwardMeta & forwardWaymask_3 | io_metaReadResp_3_valid; // @[src/main/scala/nutcore/mem/Cache.scala 187:22]
  wire  _hitVec_T_2 = metaWay_0_valid & metaWay_0_tag == addr_tag & io_in_valid; // @[src/main/scala/nutcore/mem/Cache.scala 190:73]
  wire  _hitVec_T_5 = metaWay_1_valid & metaWay_1_tag == addr_tag & io_in_valid; // @[src/main/scala/nutcore/mem/Cache.scala 190:73]
  wire  _hitVec_T_8 = metaWay_2_valid & metaWay_2_tag == addr_tag & io_in_valid; // @[src/main/scala/nutcore/mem/Cache.scala 190:73]
  wire  _hitVec_T_11 = metaWay_3_valid & metaWay_3_tag == addr_tag & io_in_valid; // @[src/main/scala/nutcore/mem/Cache.scala 190:73]
  wire [3:0] hitVec = {_hitVec_T_11,_hitVec_T_8,_hitVec_T_5,_hitVec_T_2}; // @[src/main/scala/nutcore/mem/Cache.scala 190:90]
  reg [63:0] victimWaymask_lfsr; // @[src/main/scala/utils/LFSR64.scala 25:23]
  wire  victimWaymask_xor = victimWaymask_lfsr[0] ^ victimWaymask_lfsr[1] ^ victimWaymask_lfsr[3] ^ victimWaymask_lfsr[4
    ]; // @[src/main/scala/utils/LFSR64.scala 26:43]
  wire [63:0] _victimWaymask_lfsr_T_2 = {victimWaymask_xor,victimWaymask_lfsr[63:1]}; // @[src/main/scala/utils/LFSR64.scala 28:41]
  wire [3:0] victimWaymask = 4'h1 << victimWaymask_lfsr[1:0]; // @[src/main/scala/nutcore/mem/Cache.scala 191:42]
  wire  _invalidVec_T = ~metaWay_0_valid; // @[src/main/scala/nutcore/mem/Cache.scala 193:45]
  wire  _invalidVec_T_1 = ~metaWay_1_valid; // @[src/main/scala/nutcore/mem/Cache.scala 193:45]
  wire  _invalidVec_T_2 = ~metaWay_2_valid; // @[src/main/scala/nutcore/mem/Cache.scala 193:45]
  wire  _invalidVec_T_3 = ~metaWay_3_valid; // @[src/main/scala/nutcore/mem/Cache.scala 193:45]
  wire [3:0] invalidVec = {_invalidVec_T_3,_invalidVec_T_2,_invalidVec_T_1,_invalidVec_T}; // @[src/main/scala/nutcore/mem/Cache.scala 193:56]
  wire  hasInvalidWay = |invalidVec; // @[src/main/scala/nutcore/mem/Cache.scala 194:34]
  wire [1:0] _refillInvalidWaymask_T_3 = invalidVec >= 4'h2 ? 2'h2 : 2'h1; // @[src/main/scala/nutcore/mem/Cache.scala 197:8]
  wire [2:0] _refillInvalidWaymask_T_4 = invalidVec >= 4'h4 ? 3'h4 : {{1'd0}, _refillInvalidWaymask_T_3}; // @[src/main/scala/nutcore/mem/Cache.scala 196:8]
  wire [3:0] refillInvalidWaymask = invalidVec >= 4'h8 ? 4'h8 : {{1'd0}, _refillInvalidWaymask_T_4}; // @[src/main/scala/nutcore/mem/Cache.scala 195:33]
  wire [3:0] _waymask_T = hasInvalidWay ? refillInvalidWaymask : victimWaymask; // @[src/main/scala/nutcore/mem/Cache.scala 200:49]
  wire [3:0] waymask = io_out_bits_hit ? hitVec : _waymask_T; // @[src/main/scala/nutcore/mem/Cache.scala 200:20]
  wire [1:0] _T_7 = waymask[0] + waymask[1]; // @[src/main/scala/nutcore/mem/Cache.scala 201:16]
  wire [1:0] _T_9 = waymask[2] + waymask[3]; // @[src/main/scala/nutcore/mem/Cache.scala 201:16]
  wire [2:0] _T_11 = _T_7 + _T_9; // @[src/main/scala/nutcore/mem/Cache.scala 201:16]
  wire  _T_13 = _T_11 > 3'h1; // @[src/main/scala/nutcore/mem/Cache.scala 201:26]
  reg [63:0] c; // @[src/main/scala/utils/GTimer.scala 24:20]
  wire [63:0] _c_T_1 = c + 64'h1; // @[src/main/scala/utils/GTimer.scala 25:12]
  wire  _T_16 = ~reset; // @[src/main/scala/utils/Debug.scala 56:24]
  reg [63:0] c_1; // @[src/main/scala/utils/GTimer.scala 24:20]
  wire [63:0] _c_T_3 = c_1 + 64'h1; // @[src/main/scala/utils/GTimer.scala 25:12]
  reg [63:0] c_2; // @[src/main/scala/utils/GTimer.scala 24:20]
  wire [63:0] _c_T_5 = c_2 + 64'h1; // @[src/main/scala/utils/GTimer.scala 25:12]
  reg [63:0] c_3; // @[src/main/scala/utils/GTimer.scala 24:20]
  wire [63:0] _c_T_7 = c_3 + 64'h1; // @[src/main/scala/utils/GTimer.scala 25:12]
  reg [63:0] c_4; // @[src/main/scala/utils/GTimer.scala 24:20]
  wire [63:0] _c_T_9 = c_4 + 64'h1; // @[src/main/scala/utils/GTimer.scala 25:12]
  reg [63:0] c_5; // @[src/main/scala/utils/GTimer.scala 24:20]
  wire [63:0] _c_T_11 = c_5 + 64'h1; // @[src/main/scala/utils/GTimer.scala 25:12]
  reg [63:0] c_6; // @[src/main/scala/utils/GTimer.scala 24:20]
  wire [63:0] _c_T_13 = c_6 + 64'h1; // @[src/main/scala/utils/GTimer.scala 25:12]
  reg [63:0] c_7; // @[src/main/scala/utils/GTimer.scala 24:20]
  wire [63:0] _c_T_15 = c_7 + 64'h1; // @[src/main/scala/utils/GTimer.scala 25:12]
  reg [63:0] c_8; // @[src/main/scala/utils/GTimer.scala 24:20]
  wire [63:0] _c_T_17 = c_8 + 64'h1; // @[src/main/scala/utils/GTimer.scala 25:12]
  reg [63:0] c_9; // @[src/main/scala/utils/GTimer.scala 24:20]
  wire [63:0] _c_T_19 = c_9 + 64'h1; // @[src/main/scala/utils/GTimer.scala 25:12]
  reg [63:0] c_10; // @[src/main/scala/utils/GTimer.scala 24:20]
  wire [63:0] _c_T_21 = c_10 + 64'h1; // @[src/main/scala/utils/GTimer.scala 25:12]
  wire [31:0] _io_out_bits_mmio_T = io_in_bits_req_addr ^ 32'h30000000; // @[src/main/scala/nutcore/NutCore.scala 87:11]
  wire  _io_out_bits_mmio_T_2 = _io_out_bits_mmio_T[31:28] == 4'h0; // @[src/main/scala/nutcore/NutCore.scala 87:44]
  wire [31:0] _io_out_bits_mmio_T_3 = io_in_bits_req_addr ^ 32'h40000000; // @[src/main/scala/nutcore/NutCore.scala 87:11]
  wire  _io_out_bits_mmio_T_5 = _io_out_bits_mmio_T_3[31:30] == 2'h0; // @[src/main/scala/nutcore/NutCore.scala 87:44]
  wire [11:0] _isForwardData_T_8 = {addr_index,addr_wordIndex}; // @[src/main/scala/nutcore/mem/Cache.scala 78:35]
  wire  _isForwardData_T_10 = io_dataWriteBus_req_valid & io_dataWriteBus_req_bits_setIdx == _isForwardData_T_8; // @[src/main/scala/nutcore/mem/Cache.scala 217:13]
  wire  isForwardData = io_in_valid & _isForwardData_T_10; // @[src/main/scala/nutcore/mem/Cache.scala 216:35]
  reg  isForwardDataReg; // @[src/main/scala/nutcore/mem/Cache.scala 219:33]
  wire  _GEN_8 = isForwardData | isForwardDataReg; // @[src/main/scala/nutcore/mem/Cache.scala 220:24 219:33 220:43]
  reg [63:0] forwardDataReg_data_data; // @[src/main/scala/nutcore/mem/Cache.scala 222:33]
  reg [3:0] forwardDataReg_waymask; // @[src/main/scala/nutcore/mem/Cache.scala 222:33]
  wire  _io_in_ready_T_1 = io_out_ready & io_out_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  reg [63:0] c_11; // @[src/main/scala/utils/GTimer.scala 24:20]
  wire [63:0] _c_T_23 = c_11 + 64'h1; // @[src/main/scala/utils/GTimer.scala 25:12]
  reg [63:0] c_12; // @[src/main/scala/utils/GTimer.scala 24:20]
  wire [63:0] _c_T_25 = c_12 + 64'h1; // @[src/main/scala/utils/GTimer.scala 25:12]
  wire  _GEN_13 = _T_13 & DISPLAY_ENABLE; // @[src/main/scala/utils/Debug.scala 56:24]
  assign io_in_ready = _T_1 | _io_in_ready_T_1; // @[src/main/scala/nutcore/mem/Cache.scala 228:31]
  assign io_out_valid = io_in_valid; // @[src/main/scala/nutcore/mem/Cache.scala 227:16]
  assign io_out_bits_req_addr = io_in_bits_req_addr; // @[src/main/scala/nutcore/mem/Cache.scala 226:19]
  assign io_out_bits_req_size = io_in_bits_req_size; // @[src/main/scala/nutcore/mem/Cache.scala 226:19]
  assign io_out_bits_req_cmd = io_in_bits_req_cmd; // @[src/main/scala/nutcore/mem/Cache.scala 226:19]
  assign io_out_bits_req_wmask = io_in_bits_req_wmask; // @[src/main/scala/nutcore/mem/Cache.scala 226:19]
  assign io_out_bits_req_wdata = io_in_bits_req_wdata; // @[src/main/scala/nutcore/mem/Cache.scala 226:19]
  assign io_out_bits_metas_0_tag = pickForwardMeta & forwardWaymask_0 ? _GEN_3 : io_metaReadResp_0_tag; // @[src/main/scala/nutcore/mem/Cache.scala 187:22]
  assign io_out_bits_metas_0_valid = pickForwardMeta & forwardWaymask_0 | io_metaReadResp_0_valid; // @[src/main/scala/nutcore/mem/Cache.scala 187:22]
  assign io_out_bits_metas_0_dirty = pickForwardMeta & forwardWaymask_0 ? _GEN_5 : io_metaReadResp_0_dirty; // @[src/main/scala/nutcore/mem/Cache.scala 187:22]
  assign io_out_bits_metas_1_tag = pickForwardMeta & forwardWaymask_1 ? _GEN_3 : io_metaReadResp_1_tag; // @[src/main/scala/nutcore/mem/Cache.scala 187:22]
  assign io_out_bits_metas_1_valid = pickForwardMeta & forwardWaymask_1 | io_metaReadResp_1_valid; // @[src/main/scala/nutcore/mem/Cache.scala 187:22]
  assign io_out_bits_metas_1_dirty = pickForwardMeta & forwardWaymask_1 ? _GEN_5 : io_metaReadResp_1_dirty; // @[src/main/scala/nutcore/mem/Cache.scala 187:22]
  assign io_out_bits_metas_2_tag = pickForwardMeta & forwardWaymask_2 ? _GEN_3 : io_metaReadResp_2_tag; // @[src/main/scala/nutcore/mem/Cache.scala 187:22]
  assign io_out_bits_metas_2_valid = pickForwardMeta & forwardWaymask_2 | io_metaReadResp_2_valid; // @[src/main/scala/nutcore/mem/Cache.scala 187:22]
  assign io_out_bits_metas_2_dirty = pickForwardMeta & forwardWaymask_2 ? _GEN_5 : io_metaReadResp_2_dirty; // @[src/main/scala/nutcore/mem/Cache.scala 187:22]
  assign io_out_bits_metas_3_tag = pickForwardMeta & forwardWaymask_3 ? _GEN_3 : io_metaReadResp_3_tag; // @[src/main/scala/nutcore/mem/Cache.scala 187:22]
  assign io_out_bits_metas_3_valid = pickForwardMeta & forwardWaymask_3 | io_metaReadResp_3_valid; // @[src/main/scala/nutcore/mem/Cache.scala 187:22]
  assign io_out_bits_metas_3_dirty = pickForwardMeta & forwardWaymask_3 ? _GEN_5 : io_metaReadResp_3_dirty; // @[src/main/scala/nutcore/mem/Cache.scala 187:22]
  assign io_out_bits_datas_0_data = io_dataReadResp_0_data; // @[src/main/scala/nutcore/mem/Cache.scala 213:21]
  assign io_out_bits_datas_1_data = io_dataReadResp_1_data; // @[src/main/scala/nutcore/mem/Cache.scala 213:21]
  assign io_out_bits_datas_2_data = io_dataReadResp_2_data; // @[src/main/scala/nutcore/mem/Cache.scala 213:21]
  assign io_out_bits_datas_3_data = io_dataReadResp_3_data; // @[src/main/scala/nutcore/mem/Cache.scala 213:21]
  assign io_out_bits_hit = io_in_valid & |hitVec; // @[src/main/scala/nutcore/mem/Cache.scala 211:34]
  assign io_out_bits_waymask = io_out_bits_hit ? hitVec : _waymask_T; // @[src/main/scala/nutcore/mem/Cache.scala 200:20]
  assign io_out_bits_mmio = _io_out_bits_mmio_T_2 | _io_out_bits_mmio_T_5; // @[src/main/scala/nutcore/NutCore.scala 88:15]
  assign io_out_bits_isForwardData = isForwardDataReg | isForwardData; // @[src/main/scala/nutcore/mem/Cache.scala 223:49]
  assign io_out_bits_forwardData_data_data = isForwardData ? io_dataWriteBus_req_bits_data_data :
    forwardDataReg_data_data; // @[src/main/scala/nutcore/mem/Cache.scala 224:33]
  assign io_out_bits_forwardData_waymask = isForwardData ? io_dataWriteBus_req_bits_waymask : forwardDataReg_waymask; // @[src/main/scala/nutcore/mem/Cache.scala 224:33]
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/nutcore/mem/Cache.scala 177:33]
      isForwardMetaReg <= 1'h0; // @[src/main/scala/nutcore/mem/Cache.scala 177:33]
    end else if (_T | ~io_in_valid) begin // @[src/main/scala/nutcore/mem/Cache.scala 179:37]
      isForwardMetaReg <= 1'h0; // @[src/main/scala/nutcore/mem/Cache.scala 179:56]
    end else begin
      isForwardMetaReg <= _GEN_0;
    end
    if (isForwardMeta) begin // @[src/main/scala/nutcore/mem/Cache.scala 180:33]
      forwardMetaReg_data_tag <= io_metaWriteBus_req_bits_data_tag; // @[src/main/scala/nutcore/mem/Cache.scala 180:33]
    end
    if (isForwardMeta) begin // @[src/main/scala/nutcore/mem/Cache.scala 180:33]
      forwardMetaReg_data_dirty <= io_metaWriteBus_req_bits_data_dirty; // @[src/main/scala/nutcore/mem/Cache.scala 180:33]
    end
    if (isForwardMeta) begin // @[src/main/scala/nutcore/mem/Cache.scala 180:33]
      forwardMetaReg_waymask <= io_metaWriteBus_req_bits_waymask; // @[src/main/scala/nutcore/mem/Cache.scala 180:33]
    end
    if (reset) begin // @[src/main/scala/utils/LFSR64.scala 25:23]
      victimWaymask_lfsr <= 64'h1234567887654321; // @[src/main/scala/utils/LFSR64.scala 25:23]
    end else if (victimWaymask_lfsr == 64'h0) begin // @[src/main/scala/utils/LFSR64.scala 28:18]
      victimWaymask_lfsr <= 64'h1;
    end else begin
      victimWaymask_lfsr <= _victimWaymask_lfsr_T_2;
    end
    if (reset) begin // @[src/main/scala/utils/GTimer.scala 24:20]
      c <= 64'h0; // @[src/main/scala/utils/GTimer.scala 24:20]
    end else begin
      c <= _c_T_1; // @[src/main/scala/utils/GTimer.scala 25:7]
    end
    if (reset) begin // @[src/main/scala/utils/GTimer.scala 24:20]
      c_1 <= 64'h0; // @[src/main/scala/utils/GTimer.scala 24:20]
    end else begin
      c_1 <= _c_T_3; // @[src/main/scala/utils/GTimer.scala 25:7]
    end
    if (reset) begin // @[src/main/scala/utils/GTimer.scala 24:20]
      c_2 <= 64'h0; // @[src/main/scala/utils/GTimer.scala 24:20]
    end else begin
      c_2 <= _c_T_5; // @[src/main/scala/utils/GTimer.scala 25:7]
    end
    if (reset) begin // @[src/main/scala/utils/GTimer.scala 24:20]
      c_3 <= 64'h0; // @[src/main/scala/utils/GTimer.scala 24:20]
    end else begin
      c_3 <= _c_T_7; // @[src/main/scala/utils/GTimer.scala 25:7]
    end
    if (reset) begin // @[src/main/scala/utils/GTimer.scala 24:20]
      c_4 <= 64'h0; // @[src/main/scala/utils/GTimer.scala 24:20]
    end else begin
      c_4 <= _c_T_9; // @[src/main/scala/utils/GTimer.scala 25:7]
    end
    if (reset) begin // @[src/main/scala/utils/GTimer.scala 24:20]
      c_5 <= 64'h0; // @[src/main/scala/utils/GTimer.scala 24:20]
    end else begin
      c_5 <= _c_T_11; // @[src/main/scala/utils/GTimer.scala 25:7]
    end
    if (reset) begin // @[src/main/scala/utils/GTimer.scala 24:20]
      c_6 <= 64'h0; // @[src/main/scala/utils/GTimer.scala 24:20]
    end else begin
      c_6 <= _c_T_13; // @[src/main/scala/utils/GTimer.scala 25:7]
    end
    if (reset) begin // @[src/main/scala/utils/GTimer.scala 24:20]
      c_7 <= 64'h0; // @[src/main/scala/utils/GTimer.scala 24:20]
    end else begin
      c_7 <= _c_T_15; // @[src/main/scala/utils/GTimer.scala 25:7]
    end
    if (reset) begin // @[src/main/scala/utils/GTimer.scala 24:20]
      c_8 <= 64'h0; // @[src/main/scala/utils/GTimer.scala 24:20]
    end else begin
      c_8 <= _c_T_17; // @[src/main/scala/utils/GTimer.scala 25:7]
    end
    if (reset) begin // @[src/main/scala/utils/GTimer.scala 24:20]
      c_9 <= 64'h0; // @[src/main/scala/utils/GTimer.scala 24:20]
    end else begin
      c_9 <= _c_T_19; // @[src/main/scala/utils/GTimer.scala 25:7]
    end
    if (reset) begin // @[src/main/scala/utils/GTimer.scala 24:20]
      c_10 <= 64'h0; // @[src/main/scala/utils/GTimer.scala 24:20]
    end else begin
      c_10 <= _c_T_21; // @[src/main/scala/utils/GTimer.scala 25:7]
    end
    if (reset) begin // @[src/main/scala/nutcore/mem/Cache.scala 219:33]
      isForwardDataReg <= 1'h0; // @[src/main/scala/nutcore/mem/Cache.scala 219:33]
    end else if (_T_2) begin // @[src/main/scala/nutcore/mem/Cache.scala 221:37]
      isForwardDataReg <= 1'h0; // @[src/main/scala/nutcore/mem/Cache.scala 221:56]
    end else begin
      isForwardDataReg <= _GEN_8;
    end
    if (isForwardData) begin // @[src/main/scala/nutcore/mem/Cache.scala 222:33]
      forwardDataReg_data_data <= io_dataWriteBus_req_bits_data_data; // @[src/main/scala/nutcore/mem/Cache.scala 222:33]
    end
    if (isForwardData) begin // @[src/main/scala/nutcore/mem/Cache.scala 222:33]
      forwardDataReg_waymask <= io_dataWriteBus_req_bits_waymask; // @[src/main/scala/nutcore/mem/Cache.scala 222:33]
    end
    if (reset) begin // @[src/main/scala/utils/GTimer.scala 24:20]
      c_11 <= 64'h0; // @[src/main/scala/utils/GTimer.scala 24:20]
    end else begin
      c_11 <= _c_T_23; // @[src/main/scala/utils/GTimer.scala 25:7]
    end
    if (reset) begin // @[src/main/scala/utils/GTimer.scala 24:20]
      c_12 <= 64'h0; // @[src/main/scala/utils/GTimer.scala 24:20]
    end else begin
      c_12 <= _c_T_25; // @[src/main/scala/utils/GTimer.scala 25:7]
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_13 & DISPLAY_ENABLE & ~reset) begin
          $fwrite(32'h80000002,"[%d] CacheStage2_2: ",c); // @[src/main/scala/utils/Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_13 & _T_16) begin
          $fwrite(32'h80000002,"[ERROR] metaWay %x metat %x reqt %x\n",metaWay_0_valid,metaWay_0_tag,addr_tag); // @[src/main/scala/utils/Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_13 & DISPLAY_ENABLE & ~reset) begin
          $fwrite(32'h80000002,"[%d] CacheStage2_2: ",c_1); // @[src/main/scala/utils/Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_13 & _T_16) begin
          $fwrite(32'h80000002,"[ERROR] metaWay %x metat %x reqt %x\n",metaWay_1_valid,metaWay_1_tag,addr_tag); // @[src/main/scala/utils/Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_13 & DISPLAY_ENABLE & ~reset) begin
          $fwrite(32'h80000002,"[%d] CacheStage2_2: ",c_2); // @[src/main/scala/utils/Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_13 & _T_16) begin
          $fwrite(32'h80000002,"[ERROR] metaWay %x metat %x reqt %x\n",metaWay_2_valid,metaWay_2_tag,addr_tag); // @[src/main/scala/utils/Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_13 & DISPLAY_ENABLE & ~reset) begin
          $fwrite(32'h80000002,"[%d] CacheStage2_2: ",c_3); // @[src/main/scala/utils/Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_13 & _T_16) begin
          $fwrite(32'h80000002,"[ERROR] metaWay %x metat %x reqt %x\n",metaWay_3_valid,metaWay_3_tag,addr_tag); // @[src/main/scala/utils/Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_13 & DISPLAY_ENABLE & ~reset) begin
          $fwrite(32'h80000002,"[%d] CacheStage2_2: ",c_4); // @[src/main/scala/utils/Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_13 & _T_16) begin
          $fwrite(32'h80000002,"[ERROR] metaReadResp %x metat %x reqt %x\n",io_metaReadResp_0_valid,
            io_metaReadResp_0_tag,addr_tag); // @[src/main/scala/utils/Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_13 & DISPLAY_ENABLE & ~reset) begin
          $fwrite(32'h80000002,"[%d] CacheStage2_2: ",c_5); // @[src/main/scala/utils/Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_13 & _T_16) begin
          $fwrite(32'h80000002,"[ERROR] metaReadResp %x metat %x reqt %x\n",io_metaReadResp_1_valid,
            io_metaReadResp_1_tag,addr_tag); // @[src/main/scala/utils/Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_13 & DISPLAY_ENABLE & ~reset) begin
          $fwrite(32'h80000002,"[%d] CacheStage2_2: ",c_6); // @[src/main/scala/utils/Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_13 & _T_16) begin
          $fwrite(32'h80000002,"[ERROR] metaReadResp %x metat %x reqt %x\n",io_metaReadResp_2_valid,
            io_metaReadResp_2_tag,addr_tag); // @[src/main/scala/utils/Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_13 & DISPLAY_ENABLE & ~reset) begin
          $fwrite(32'h80000002,"[%d] CacheStage2_2: ",c_7); // @[src/main/scala/utils/Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_13 & _T_16) begin
          $fwrite(32'h80000002,"[ERROR] metaReadResp %x metat %x reqt %x\n",io_metaReadResp_3_valid,
            io_metaReadResp_3_tag,addr_tag); // @[src/main/scala/utils/Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_13 & DISPLAY_ENABLE & ~reset) begin
          $fwrite(32'h80000002,"[%d] CacheStage2_2: ",c_8); // @[src/main/scala/utils/Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_13 & _T_16) begin
          $fwrite(32'h80000002,"[ERROR] forwardMetaReg isForwardMetaReg %x %x metat %x wm %b\n",isForwardMetaReg,1'h1,
            forwardMetaReg_data_tag,forwardMetaReg_waymask); // @[src/main/scala/utils/Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_13 & DISPLAY_ENABLE & ~reset) begin
          $fwrite(32'h80000002,"[%d] CacheStage2_2: ",c_9); // @[src/main/scala/utils/Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_13 & _T_16) begin
          $fwrite(32'h80000002,"[ERROR] forwardMeta isForwardMeta %x %x metat %x wm %b\n",isForwardMeta,1'h1,
            io_metaWriteBus_req_bits_data_tag,io_metaWriteBus_req_bits_waymask); // @[src/main/scala/utils/Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_13 & DISPLAY_ENABLE & ~reset) begin
          $fwrite(32'h80000002,"[%d] CacheStage2_2: ",c_10); // @[src/main/scala/utils/Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_13 & _T_16) begin
          $fwrite(32'h80000002,"[ERROR] hit %b wmask %b hitvec %b\n",io_out_bits_hit,_GEN_6,hitVec); // @[src/main/scala/utils/Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_16 & ~(~(io_in_valid & _T_13))) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Cache.scala:208 assert(!(io.in.valid && PopCount(waymask) > 1.U))\n"); // @[src/main/scala/nutcore/mem/Cache.scala 208:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~(io_in_valid & _T_13)) & _T_16) begin
          $fatal; // @[src/main/scala/nutcore/mem/Cache.scala 208:9]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & ~reset) begin
          $fwrite(32'h80000002,"[%d] CacheStage2_2: ",c_11); // @[src/main/scala/utils/Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_16) begin
          $fwrite(32'h80000002,"[isFD:%d isFDreg:%d inFire:%d invalid:%d \n",isForwardData,isForwardDataReg,_T,
            io_in_valid); // @[src/main/scala/utils/Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & ~reset) begin
          $fwrite(32'h80000002,"[%d] CacheStage2_2: ",c_12); // @[src/main/scala/utils/Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_16) begin
          $fwrite(32'h80000002,"[isFM:%d isFMreg:%d metawreq:%x widx:%x ridx:%x \n",isForwardMeta,isForwardMetaReg,
            io_metaWriteBus_req_valid,io_metaWriteBus_req_bits_setIdx,addr_index); // @[src/main/scala/utils/Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  isForwardMetaReg = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  forwardMetaReg_data_tag = _RAND_1[16:0];
  _RAND_2 = {1{`RANDOM}};
  forwardMetaReg_data_dirty = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  forwardMetaReg_waymask = _RAND_3[3:0];
  _RAND_4 = {2{`RANDOM}};
  victimWaymask_lfsr = _RAND_4[63:0];
  _RAND_5 = {2{`RANDOM}};
  c = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  c_1 = _RAND_6[63:0];
  _RAND_7 = {2{`RANDOM}};
  c_2 = _RAND_7[63:0];
  _RAND_8 = {2{`RANDOM}};
  c_3 = _RAND_8[63:0];
  _RAND_9 = {2{`RANDOM}};
  c_4 = _RAND_9[63:0];
  _RAND_10 = {2{`RANDOM}};
  c_5 = _RAND_10[63:0];
  _RAND_11 = {2{`RANDOM}};
  c_6 = _RAND_11[63:0];
  _RAND_12 = {2{`RANDOM}};
  c_7 = _RAND_12[63:0];
  _RAND_13 = {2{`RANDOM}};
  c_8 = _RAND_13[63:0];
  _RAND_14 = {2{`RANDOM}};
  c_9 = _RAND_14[63:0];
  _RAND_15 = {2{`RANDOM}};
  c_10 = _RAND_15[63:0];
  _RAND_16 = {1{`RANDOM}};
  isForwardDataReg = _RAND_16[0:0];
  _RAND_17 = {2{`RANDOM}};
  forwardDataReg_data_data = _RAND_17[63:0];
  _RAND_18 = {1{`RANDOM}};
  forwardDataReg_waymask = _RAND_18[3:0];
  _RAND_19 = {2{`RANDOM}};
  c_11 = _RAND_19[63:0];
  _RAND_20 = {2{`RANDOM}};
  c_12 = _RAND_20[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Arbiter_10(
  input         io_in_0_valid, // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
  input  [8:0]  io_in_0_bits_setIdx, // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
  input  [16:0] io_in_0_bits_data_tag, // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
  input  [3:0]  io_in_0_bits_waymask, // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
  input         io_in_1_valid, // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
  input  [8:0]  io_in_1_bits_setIdx, // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
  input  [16:0] io_in_1_bits_data_tag, // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
  input         io_in_1_bits_data_dirty, // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
  input  [3:0]  io_in_1_bits_waymask, // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
  output        io_out_valid, // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
  output [8:0]  io_out_bits_setIdx, // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
  output [16:0] io_out_bits_data_tag, // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
  output        io_out_bits_data_dirty, // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
  output [3:0]  io_out_bits_waymask // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
);
  wire  grant_1 = ~io_in_0_valid; // @[src/main/scala/chisel3/util/Arbiter.scala 45:78]
  assign io_out_valid = ~grant_1 | io_in_1_valid; // @[src/main/scala/chisel3/util/Arbiter.scala 148:31]
  assign io_out_bits_setIdx = io_in_0_valid ? io_in_0_bits_setIdx : io_in_1_bits_setIdx; // @[src/main/scala/chisel3/util/Arbiter.scala 137:15 139:26 141:19]
  assign io_out_bits_data_tag = io_in_0_valid ? io_in_0_bits_data_tag : io_in_1_bits_data_tag; // @[src/main/scala/chisel3/util/Arbiter.scala 137:15 139:26 141:19]
  assign io_out_bits_data_dirty = io_in_0_valid | io_in_1_bits_data_dirty; // @[src/main/scala/chisel3/util/Arbiter.scala 137:15 139:26 141:19]
  assign io_out_bits_waymask = io_in_0_valid ? io_in_0_bits_waymask : io_in_1_bits_waymask; // @[src/main/scala/chisel3/util/Arbiter.scala 137:15 139:26 141:19]
endmodule
module Arbiter_11(
  input         io_in_0_valid, // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
  input  [11:0] io_in_0_bits_setIdx, // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
  input  [63:0] io_in_0_bits_data_data, // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
  input  [3:0]  io_in_0_bits_waymask, // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
  input         io_in_1_valid, // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
  input  [11:0] io_in_1_bits_setIdx, // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
  input  [63:0] io_in_1_bits_data_data, // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
  input  [3:0]  io_in_1_bits_waymask, // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
  output        io_out_valid, // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
  output [11:0] io_out_bits_setIdx, // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
  output [63:0] io_out_bits_data_data, // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
  output [3:0]  io_out_bits_waymask // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
);
  wire  grant_1 = ~io_in_0_valid; // @[src/main/scala/chisel3/util/Arbiter.scala 45:78]
  assign io_out_valid = ~grant_1 | io_in_1_valid; // @[src/main/scala/chisel3/util/Arbiter.scala 148:31]
  assign io_out_bits_setIdx = io_in_0_valid ? io_in_0_bits_setIdx : io_in_1_bits_setIdx; // @[src/main/scala/chisel3/util/Arbiter.scala 137:15 139:26 141:19]
  assign io_out_bits_data_data = io_in_0_valid ? io_in_0_bits_data_data : io_in_1_bits_data_data; // @[src/main/scala/chisel3/util/Arbiter.scala 137:15 139:26 141:19]
  assign io_out_bits_waymask = io_in_0_valid ? io_in_0_bits_waymask : io_in_1_bits_waymask; // @[src/main/scala/chisel3/util/Arbiter.scala 137:15 139:26 141:19]
endmodule
module CacheStage3_2(
  input         clock,
  input         reset,
  output        io_in_ready, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  input         io_in_valid, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  input  [31:0] io_in_bits_req_addr, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  input  [2:0]  io_in_bits_req_size, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  input  [3:0]  io_in_bits_req_cmd, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  input  [7:0]  io_in_bits_req_wmask, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  input  [63:0] io_in_bits_req_wdata, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  input  [16:0] io_in_bits_metas_0_tag, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  input         io_in_bits_metas_0_valid, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  input         io_in_bits_metas_0_dirty, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  input  [16:0] io_in_bits_metas_1_tag, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  input         io_in_bits_metas_1_valid, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  input         io_in_bits_metas_1_dirty, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  input  [16:0] io_in_bits_metas_2_tag, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  input         io_in_bits_metas_2_valid, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  input         io_in_bits_metas_2_dirty, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  input  [16:0] io_in_bits_metas_3_tag, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  input         io_in_bits_metas_3_valid, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  input         io_in_bits_metas_3_dirty, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  input  [63:0] io_in_bits_datas_0_data, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  input  [63:0] io_in_bits_datas_1_data, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  input  [63:0] io_in_bits_datas_2_data, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  input  [63:0] io_in_bits_datas_3_data, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  input         io_in_bits_hit, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  input  [3:0]  io_in_bits_waymask, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  input         io_in_bits_mmio, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  input         io_in_bits_isForwardData, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  input  [63:0] io_in_bits_forwardData_data_data, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  input  [3:0]  io_in_bits_forwardData_waymask, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  input         io_out_ready, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  output        io_out_valid, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  output [3:0]  io_out_bits_cmd, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  output [63:0] io_out_bits_rdata, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  output        io_isFinish, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  input         io_dataReadBus_req_ready, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  output        io_dataReadBus_req_valid, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  output [11:0] io_dataReadBus_req_bits_setIdx, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  input  [63:0] io_dataReadBus_resp_data_0_data, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  input  [63:0] io_dataReadBus_resp_data_1_data, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  input  [63:0] io_dataReadBus_resp_data_2_data, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  input  [63:0] io_dataReadBus_resp_data_3_data, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  output        io_dataWriteBus_req_valid, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  output [11:0] io_dataWriteBus_req_bits_setIdx, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  output [63:0] io_dataWriteBus_req_bits_data_data, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  output [3:0]  io_dataWriteBus_req_bits_waymask, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  output        io_metaWriteBus_req_valid, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  output [8:0]  io_metaWriteBus_req_bits_setIdx, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  output [16:0] io_metaWriteBus_req_bits_data_tag, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  output        io_metaWriteBus_req_bits_data_valid, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  output        io_metaWriteBus_req_bits_data_dirty, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  output [3:0]  io_metaWriteBus_req_bits_waymask, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  input         io_mem_req_ready, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  output        io_mem_req_valid, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  output [31:0] io_mem_req_bits_addr, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  output [2:0]  io_mem_req_bits_size, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  output [3:0]  io_mem_req_bits_cmd, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  output [7:0]  io_mem_req_bits_wmask, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  output [63:0] io_mem_req_bits_wdata, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  output        io_mem_resp_ready, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  input         io_mem_resp_valid, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  input  [3:0]  io_mem_resp_bits_cmd, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  input  [63:0] io_mem_resp_bits_rdata, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  output        io_cohResp_valid, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  output        io_dataReadRespToL1, // @[src/main/scala/nutcore/mem/Cache.scala 252:14]
  input         DISPLAY_ENABLE
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [63:0] _RAND_14;
  reg [63:0] _RAND_15;
  reg [63:0] _RAND_16;
  reg [63:0] _RAND_17;
  reg [63:0] _RAND_18;
  reg [63:0] _RAND_19;
  reg [63:0] _RAND_20;
  reg [63:0] _RAND_21;
  reg [63:0] _RAND_22;
  reg [63:0] _RAND_23;
  reg [63:0] _RAND_24;
  reg [63:0] _RAND_25;
`endif // RANDOMIZE_REG_INIT
  wire  metaWriteArb_io_in_0_valid; // @[src/main/scala/nutcore/mem/Cache.scala 254:28]
  wire [8:0] metaWriteArb_io_in_0_bits_setIdx; // @[src/main/scala/nutcore/mem/Cache.scala 254:28]
  wire [16:0] metaWriteArb_io_in_0_bits_data_tag; // @[src/main/scala/nutcore/mem/Cache.scala 254:28]
  wire [3:0] metaWriteArb_io_in_0_bits_waymask; // @[src/main/scala/nutcore/mem/Cache.scala 254:28]
  wire  metaWriteArb_io_in_1_valid; // @[src/main/scala/nutcore/mem/Cache.scala 254:28]
  wire [8:0] metaWriteArb_io_in_1_bits_setIdx; // @[src/main/scala/nutcore/mem/Cache.scala 254:28]
  wire [16:0] metaWriteArb_io_in_1_bits_data_tag; // @[src/main/scala/nutcore/mem/Cache.scala 254:28]
  wire  metaWriteArb_io_in_1_bits_data_dirty; // @[src/main/scala/nutcore/mem/Cache.scala 254:28]
  wire [3:0] metaWriteArb_io_in_1_bits_waymask; // @[src/main/scala/nutcore/mem/Cache.scala 254:28]
  wire  metaWriteArb_io_out_valid; // @[src/main/scala/nutcore/mem/Cache.scala 254:28]
  wire [8:0] metaWriteArb_io_out_bits_setIdx; // @[src/main/scala/nutcore/mem/Cache.scala 254:28]
  wire [16:0] metaWriteArb_io_out_bits_data_tag; // @[src/main/scala/nutcore/mem/Cache.scala 254:28]
  wire  metaWriteArb_io_out_bits_data_dirty; // @[src/main/scala/nutcore/mem/Cache.scala 254:28]
  wire [3:0] metaWriteArb_io_out_bits_waymask; // @[src/main/scala/nutcore/mem/Cache.scala 254:28]
  wire  dataWriteArb_io_in_0_valid; // @[src/main/scala/nutcore/mem/Cache.scala 255:28]
  wire [11:0] dataWriteArb_io_in_0_bits_setIdx; // @[src/main/scala/nutcore/mem/Cache.scala 255:28]
  wire [63:0] dataWriteArb_io_in_0_bits_data_data; // @[src/main/scala/nutcore/mem/Cache.scala 255:28]
  wire [3:0] dataWriteArb_io_in_0_bits_waymask; // @[src/main/scala/nutcore/mem/Cache.scala 255:28]
  wire  dataWriteArb_io_in_1_valid; // @[src/main/scala/nutcore/mem/Cache.scala 255:28]
  wire [11:0] dataWriteArb_io_in_1_bits_setIdx; // @[src/main/scala/nutcore/mem/Cache.scala 255:28]
  wire [63:0] dataWriteArb_io_in_1_bits_data_data; // @[src/main/scala/nutcore/mem/Cache.scala 255:28]
  wire [3:0] dataWriteArb_io_in_1_bits_waymask; // @[src/main/scala/nutcore/mem/Cache.scala 255:28]
  wire  dataWriteArb_io_out_valid; // @[src/main/scala/nutcore/mem/Cache.scala 255:28]
  wire [11:0] dataWriteArb_io_out_bits_setIdx; // @[src/main/scala/nutcore/mem/Cache.scala 255:28]
  wire [63:0] dataWriteArb_io_out_bits_data_data; // @[src/main/scala/nutcore/mem/Cache.scala 255:28]
  wire [3:0] dataWriteArb_io_out_bits_waymask; // @[src/main/scala/nutcore/mem/Cache.scala 255:28]
  wire [2:0] addr_wordIndex = io_in_bits_req_addr[5:3]; // @[src/main/scala/nutcore/mem/Cache.scala 258:31]
  wire [8:0] addr_index = io_in_bits_req_addr[14:6]; // @[src/main/scala/nutcore/mem/Cache.scala 258:31]
  wire [16:0] addr_tag = io_in_bits_req_addr[31:15]; // @[src/main/scala/nutcore/mem/Cache.scala 258:31]
  wire  mmio = io_in_valid & io_in_bits_mmio; // @[src/main/scala/nutcore/mem/Cache.scala 259:26]
  wire  hit = io_in_valid & io_in_bits_hit; // @[src/main/scala/nutcore/mem/Cache.scala 260:25]
  wire  miss = io_in_valid & ~io_in_bits_hit; // @[src/main/scala/nutcore/mem/Cache.scala 261:26]
  wire  _probe_T_1 = io_in_bits_req_cmd == 4'h8; // @[src/main/scala/bus/simplebus/SimpleBus.scala 79:23]
  wire  probe = io_in_valid & _probe_T_1; // @[src/main/scala/nutcore/mem/Cache.scala 262:39]
  wire  _hitReadBurst_T = io_in_bits_req_cmd == 4'h2; // @[src/main/scala/bus/simplebus/SimpleBus.scala 76:27]
  wire  hitReadBurst = hit & _hitReadBurst_T; // @[src/main/scala/nutcore/mem/Cache.scala 263:26]
  wire  meta_dirty = io_in_bits_waymask[0] & io_in_bits_metas_0_dirty | io_in_bits_waymask[1] & io_in_bits_metas_1_dirty
     | io_in_bits_waymask[2] & io_in_bits_metas_2_dirty | io_in_bits_waymask[3] & io_in_bits_metas_3_dirty; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [16:0] _meta_T_18 = io_in_bits_waymask[0] ? io_in_bits_metas_0_tag : 17'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [16:0] _meta_T_19 = io_in_bits_waymask[1] ? io_in_bits_metas_1_tag : 17'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [16:0] _meta_T_20 = io_in_bits_waymask[2] ? io_in_bits_metas_2_tag : 17'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [16:0] _meta_T_21 = io_in_bits_waymask[3] ? io_in_bits_metas_3_tag : 17'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [16:0] _meta_T_22 = _meta_T_18 | _meta_T_19; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [16:0] _meta_T_23 = _meta_T_22 | _meta_T_20; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [16:0] meta_tag = _meta_T_23 | _meta_T_21; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _T_3 = ~reset; // @[src/main/scala/nutcore/mem/Cache.scala 265:9]
  wire  useForwardData = io_in_bits_isForwardData & io_in_bits_waymask == io_in_bits_forwardData_waymask; // @[src/main/scala/nutcore/mem/Cache.scala 273:49]
  wire [63:0] _dataReadArray_T_4 = io_in_bits_waymask[0] ? io_in_bits_datas_0_data : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _dataReadArray_T_5 = io_in_bits_waymask[1] ? io_in_bits_datas_1_data : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _dataReadArray_T_6 = io_in_bits_waymask[2] ? io_in_bits_datas_2_data : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _dataReadArray_T_7 = io_in_bits_waymask[3] ? io_in_bits_datas_3_data : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _dataReadArray_T_8 = _dataReadArray_T_4 | _dataReadArray_T_5; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _dataReadArray_T_9 = _dataReadArray_T_8 | _dataReadArray_T_6; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _dataReadArray_T_10 = _dataReadArray_T_9 | _dataReadArray_T_7; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] dataRead = useForwardData ? io_in_bits_forwardData_data_data : _dataReadArray_T_10; // @[src/main/scala/nutcore/mem/Cache.scala 275:21]
  wire [7:0] _wordMask_T_12 = io_in_bits_req_wmask[0] ? 8'hff : 8'h0; // @[src/main/scala/utils/BitUtils.scala 27:45]
  wire [7:0] _wordMask_T_14 = io_in_bits_req_wmask[1] ? 8'hff : 8'h0; // @[src/main/scala/utils/BitUtils.scala 27:45]
  wire [7:0] _wordMask_T_16 = io_in_bits_req_wmask[2] ? 8'hff : 8'h0; // @[src/main/scala/utils/BitUtils.scala 27:45]
  wire [7:0] _wordMask_T_18 = io_in_bits_req_wmask[3] ? 8'hff : 8'h0; // @[src/main/scala/utils/BitUtils.scala 27:45]
  wire [7:0] _wordMask_T_20 = io_in_bits_req_wmask[4] ? 8'hff : 8'h0; // @[src/main/scala/utils/BitUtils.scala 27:45]
  wire [7:0] _wordMask_T_22 = io_in_bits_req_wmask[5] ? 8'hff : 8'h0; // @[src/main/scala/utils/BitUtils.scala 27:45]
  wire [7:0] _wordMask_T_24 = io_in_bits_req_wmask[6] ? 8'hff : 8'h0; // @[src/main/scala/utils/BitUtils.scala 27:45]
  wire [7:0] _wordMask_T_26 = io_in_bits_req_wmask[7] ? 8'hff : 8'h0; // @[src/main/scala/utils/BitUtils.scala 27:45]
  wire [63:0] _wordMask_T_27 = {_wordMask_T_26,_wordMask_T_24,_wordMask_T_22,_wordMask_T_20,_wordMask_T_18,
    _wordMask_T_16,_wordMask_T_14,_wordMask_T_12}; // @[src/main/scala/utils/BitUtils.scala 27:26]
  wire [63:0] wordMask = io_in_bits_req_cmd[0] ? _wordMask_T_27 : 64'h0; // @[src/main/scala/nutcore/mem/Cache.scala 276:21]
  reg [2:0] writeL2BeatCnt_value; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
  wire  _T_6 = io_in_bits_req_cmd == 4'h3; // @[src/main/scala/nutcore/mem/Cache.scala 279:32]
  wire  _T_7 = io_in_bits_req_cmd == 4'h7; // @[src/main/scala/bus/simplebus/SimpleBus.scala 78:27]
  wire  _T_8 = io_in_bits_req_cmd == 4'h3 | _T_7; // @[src/main/scala/nutcore/mem/Cache.scala 279:60]
  wire [2:0] _value_T_1 = writeL2BeatCnt_value + 3'h1; // @[src/main/scala/chisel3/util/Counter.scala 77:24]
  wire [2:0] _GEN_0 = io_out_valid & (io_in_bits_req_cmd == 4'h3 | _T_7) ? _value_T_1 : writeL2BeatCnt_value; // @[src/main/scala/nutcore/mem/Cache.scala 279:83 src/main/scala/chisel3/util/Counter.scala 77:15 61:40]
  wire  hitWrite = hit & io_in_bits_req_cmd[0]; // @[src/main/scala/nutcore/mem/Cache.scala 283:22]
  wire [63:0] _dataHitWriteBus_x1_T = io_in_bits_req_wdata & wordMask; // @[src/main/scala/utils/BitUtils.scala 34:14]
  wire [63:0] _dataHitWriteBus_x1_T_1 = ~wordMask; // @[src/main/scala/utils/BitUtils.scala 34:39]
  wire [63:0] _dataHitWriteBus_x1_T_2 = dataRead & _dataHitWriteBus_x1_T_1; // @[src/main/scala/utils/BitUtils.scala 34:37]
  wire [63:0] dataHitWriteBus_x1_data = _dataHitWriteBus_x1_T | _dataHitWriteBus_x1_T_2; // @[src/main/scala/utils/BitUtils.scala 34:26]
  wire [2:0] _dataHitWriteBus_x3_T_3 = _T_8 ? writeL2BeatCnt_value : addr_wordIndex; // @[src/main/scala/nutcore/mem/Cache.scala 286:51]
  wire [11:0] dataHitWriteBus_x3 = {addr_index,_dataHitWriteBus_x3_T_3}; // @[src/main/scala/nutcore/mem/Cache.scala 286:35]
  wire  metaHitWriteBus_x5 = hitWrite & ~meta_dirty; // @[src/main/scala/nutcore/mem/Cache.scala 289:22]
  reg [3:0] state; // @[src/main/scala/nutcore/mem/Cache.scala 294:22]
  reg [2:0] readBeatCnt_value; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
  reg [2:0] writeBeatCnt_value; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
  reg [1:0] state2; // @[src/main/scala/nutcore/mem/Cache.scala 304:23]
  wire  _T_14 = state == 4'h3; // @[src/main/scala/nutcore/mem/Cache.scala 306:39]
  wire  _T_15 = state == 4'h8; // @[src/main/scala/nutcore/mem/Cache.scala 306:66]
  wire [2:0] _T_20 = _T_15 ? readBeatCnt_value : writeBeatCnt_value; // @[src/main/scala/nutcore/mem/Cache.scala 307:33]
  reg [63:0] dataWay_0_data; // @[src/main/scala/nutcore/mem/Cache.scala 308:26]
  reg [63:0] dataWay_1_data; // @[src/main/scala/nutcore/mem/Cache.scala 308:26]
  reg [63:0] dataWay_2_data; // @[src/main/scala/nutcore/mem/Cache.scala 308:26]
  reg [63:0] dataWay_3_data; // @[src/main/scala/nutcore/mem/Cache.scala 308:26]
  wire [63:0] _dataHitWay_T_4 = io_in_bits_waymask[0] ? dataWay_0_data : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _dataHitWay_T_5 = io_in_bits_waymask[1] ? dataWay_1_data : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _dataHitWay_T_6 = io_in_bits_waymask[2] ? dataWay_2_data : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _dataHitWay_T_7 = io_in_bits_waymask[3] ? dataWay_3_data : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _dataHitWay_T_8 = _dataHitWay_T_4 | _dataHitWay_T_5; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _dataHitWay_T_9 = _dataHitWay_T_8 | _dataHitWay_T_6; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _dataHitWay_T_10 = _dataHitWay_T_9 | _dataHitWay_T_7; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _T_23 = io_dataReadBus_req_ready & io_dataReadBus_req_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  wire  _T_26 = io_mem_req_ready & io_mem_req_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  wire [1:0] _GEN_8 = _T_26 | io_cohResp_valid | hitReadBurst ? 2'h0 : state2; // @[src/main/scala/nutcore/mem/Cache.scala 314:105 304:23 314:96]
  wire [31:0] raddr = {io_in_bits_req_addr[31:3],3'h0}; // @[src/main/scala/nutcore/mem/Cache.scala 318:35]
  wire [31:0] waddr = {meta_tag,addr_index,6'h0}; // @[src/main/scala/nutcore/mem/Cache.scala 321:18]
  wire  _cmd_T = state == 4'h1; // @[src/main/scala/nutcore/mem/Cache.scala 322:23]
  wire [2:0] _cmd_T_2 = writeBeatCnt_value == 3'h7 ? 3'h7 : 3'h3; // @[src/main/scala/nutcore/mem/Cache.scala 323:8]
  wire [2:0] cmd = state == 4'h1 ? 3'h2 : _cmd_T_2; // @[src/main/scala/nutcore/mem/Cache.scala 322:16]
  wire  _io_mem_req_valid_T_2 = state2 == 2'h2; // @[src/main/scala/nutcore/mem/Cache.scala 329:89]
  reg  afterFirstRead; // @[src/main/scala/nutcore/mem/Cache.scala 336:31]
  reg  alreadyOutFire; // @[src/main/scala/nutcore/mem/Cache.scala 337:33]
  wire  _GEN_12 = io_out_valid | alreadyOutFire; // @[src/main/scala/nutcore/mem/Cache.scala 337:{33,33,33}]
  wire  _readingFirst_T_1 = io_mem_resp_ready & io_mem_resp_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  wire  _readingFirst_T_3 = state == 4'h2; // @[src/main/scala/nutcore/mem/Cache.scala 338:68]
  wire  readingFirst = ~afterFirstRead & _readingFirst_T_1 & state == 4'h2; // @[src/main/scala/nutcore/mem/Cache.scala 338:58]
  wire  _inRdataRegDemand_T_2 = mmio ? state == 4'h6 : readingFirst; // @[src/main/scala/nutcore/mem/Cache.scala 340:39]
  reg [63:0] inRdataRegDemand; // @[src/main/scala/nutcore/mem/Cache.scala 339:35]
  wire  _io_cohResp_valid_T = state == 4'h0; // @[src/main/scala/nutcore/mem/Cache.scala 343:31]
  wire  _io_cohResp_valid_T_4 = _T_15 & _io_mem_req_valid_T_2; // @[src/main/scala/nutcore/mem/Cache.scala 344:46]
  wire  _releaseLast_T_2 = _T_15 & io_cohResp_valid; // @[src/main/scala/nutcore/mem/Cache.scala 346:49]
  reg [2:0] releaseLast_c_value; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
  wire  releaseLast_wrap_wrap = releaseLast_c_value == 3'h7; // @[src/main/scala/chisel3/util/Counter.scala 73:24]
  wire [2:0] _releaseLast_wrap_value_T_1 = releaseLast_c_value + 3'h1; // @[src/main/scala/chisel3/util/Counter.scala 77:24]
  wire  releaseLast = _releaseLast_T_2 & releaseLast_wrap_wrap; // @[src/main/scala/chisel3/util/Counter.scala 118:{16,23} 117:24]
  wire  respToL1Fire = hitReadBurst & _io_mem_req_valid_T_2; // @[src/main/scala/nutcore/mem/Cache.scala 350:51]
  wire  _respToL1Last_T_4 = _io_cohResp_valid_T | _io_cohResp_valid_T_4; // @[src/main/scala/nutcore/mem/Cache.scala 351:48]
  wire  _respToL1Last_T_5 = (_io_cohResp_valid_T | _io_cohResp_valid_T_4) & hitReadBurst; // @[src/main/scala/nutcore/mem/Cache.scala 351:96]
  reg [2:0] respToL1Last_c_value; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
  wire  respToL1Last_wrap_wrap = respToL1Last_c_value == 3'h7; // @[src/main/scala/chisel3/util/Counter.scala 73:24]
  wire [2:0] _respToL1Last_wrap_value_T_1 = respToL1Last_c_value + 3'h1; // @[src/main/scala/chisel3/util/Counter.scala 77:24]
  wire  respToL1Last = _respToL1Last_T_5 & respToL1Last_wrap_wrap; // @[src/main/scala/chisel3/util/Counter.scala 118:{16,23} 117:24]
  wire [3:0] _state_T = hit ? 4'h8 : 4'h0; // @[src/main/scala/nutcore/mem/Cache.scala 360:23]
  wire [2:0] _value_T_4 = addr_wordIndex + 3'h1; // @[src/main/scala/nutcore/mem/Cache.scala 365:93]
  wire [2:0] _value_T_5 = addr_wordIndex == 3'h7 ? 3'h0 : _value_T_4; // @[src/main/scala/nutcore/mem/Cache.scala 365:33]
  wire [3:0] _state_T_3 = meta_dirty ? 4'h3 : 4'h1; // @[src/main/scala/nutcore/mem/Cache.scala 367:42]
  wire [3:0] _state_T_4 = mmio ? 4'h5 : _state_T_3; // @[src/main/scala/nutcore/mem/Cache.scala 367:21]
  wire [3:0] _GEN_20 = miss | mmio ? _state_T_4 : state; // @[src/main/scala/nutcore/mem/Cache.scala 366:49 367:15 294:22]
  wire [2:0] _value_T_7 = readBeatCnt_value + 3'h1; // @[src/main/scala/chisel3/util/Counter.scala 77:24]
  wire [2:0] _GEN_27 = io_cohResp_valid | respToL1Fire ? _value_T_7 : readBeatCnt_value; // @[src/main/scala/nutcore/mem/Cache.scala 375:46 src/main/scala/chisel3/util/Counter.scala 77:15 61:40]
  wire  _T_50 = respToL1Fire & respToL1Last; // @[src/main/scala/nutcore/mem/Cache.scala 376:69]
  wire [3:0] _GEN_28 = probe & io_cohResp_valid & releaseLast | respToL1Fire & respToL1Last ? 4'h0 : state; // @[src/main/scala/nutcore/mem/Cache.scala 294:22 376:{86,94}]
  wire [3:0] _GEN_29 = _T_26 ? 4'h2 : state; // @[src/main/scala/nutcore/mem/Cache.scala 379:48 380:13 294:22]
  wire [2:0] _GEN_30 = _T_26 ? addr_wordIndex : readBeatCnt_value; // @[src/main/scala/nutcore/mem/Cache.scala 379:48 381:25 src/main/scala/chisel3/util/Counter.scala 61:40]
  wire [2:0] _GEN_31 = _T_6 ? 3'h0 : _GEN_0; // @[src/main/scala/nutcore/mem/Cache.scala 388:{52,75}]
  wire  _T_57 = io_mem_resp_bits_cmd == 4'h6; // @[src/main/scala/bus/simplebus/SimpleBus.scala 91:24]
  wire [3:0] _GEN_32 = _T_57 ? 4'h7 : state; // @[src/main/scala/nutcore/mem/Cache.scala 294:22 389:{44,52}]
  wire  _GEN_33 = _readingFirst_T_1 | afterFirstRead; // @[src/main/scala/nutcore/mem/Cache.scala 385:31 386:24 336:31]
  wire [2:0] _GEN_34 = _readingFirst_T_1 ? _value_T_7 : readBeatCnt_value; // @[src/main/scala/nutcore/mem/Cache.scala 385:31 src/main/scala/chisel3/util/Counter.scala 77:15 61:40]
  wire [2:0] _GEN_35 = _readingFirst_T_1 ? _GEN_31 : _GEN_0; // @[src/main/scala/nutcore/mem/Cache.scala 385:31]
  wire [3:0] _GEN_36 = _readingFirst_T_1 ? _GEN_32 : state; // @[src/main/scala/nutcore/mem/Cache.scala 294:22 385:31]
  wire [2:0] _value_T_11 = writeBeatCnt_value + 3'h1; // @[src/main/scala/chisel3/util/Counter.scala 77:24]
  wire [2:0] _GEN_37 = _T_26 ? _value_T_11 : writeBeatCnt_value; // @[src/main/scala/nutcore/mem/Cache.scala 394:30 src/main/scala/chisel3/util/Counter.scala 77:15 61:40]
  wire  _T_60 = io_mem_req_bits_cmd == 4'h7; // @[src/main/scala/bus/simplebus/SimpleBus.scala 78:27]
  wire [3:0] _GEN_38 = _T_60 & _T_26 ? 4'h4 : state; // @[src/main/scala/nutcore/mem/Cache.scala 294:22 395:{63,71}]
  wire [3:0] _GEN_39 = _readingFirst_T_1 ? 4'h1 : state; // @[src/main/scala/nutcore/mem/Cache.scala 294:22 398:{51,59}]
  wire [3:0] _GEN_40 = _GEN_12 ? 4'h0 : state; // @[src/main/scala/nutcore/mem/Cache.scala 294:22 399:{74,82}]
  wire [3:0] _GEN_41 = 4'h7 == state ? _GEN_40 : state; // @[src/main/scala/nutcore/mem/Cache.scala 353:18 294:22]
  wire [3:0] _GEN_42 = 4'h4 == state ? _GEN_39 : _GEN_41; // @[src/main/scala/nutcore/mem/Cache.scala 353:18]
  wire [2:0] _GEN_43 = 4'h3 == state ? _GEN_37 : writeBeatCnt_value; // @[src/main/scala/nutcore/mem/Cache.scala 353:18 src/main/scala/chisel3/util/Counter.scala 61:40]
  wire [3:0] _GEN_44 = 4'h3 == state ? _GEN_38 : _GEN_42; // @[src/main/scala/nutcore/mem/Cache.scala 353:18]
  wire  _GEN_45 = 4'h2 == state ? _GEN_33 : afterFirstRead; // @[src/main/scala/nutcore/mem/Cache.scala 353:18 336:31]
  wire [2:0] _GEN_46 = 4'h2 == state ? _GEN_34 : readBeatCnt_value; // @[src/main/scala/nutcore/mem/Cache.scala 353:18 src/main/scala/chisel3/util/Counter.scala 61:40]
  wire [2:0] _GEN_47 = 4'h2 == state ? _GEN_35 : _GEN_0; // @[src/main/scala/nutcore/mem/Cache.scala 353:18]
  wire [3:0] _GEN_48 = 4'h2 == state ? _GEN_36 : _GEN_44; // @[src/main/scala/nutcore/mem/Cache.scala 353:18]
  wire [2:0] _GEN_49 = 4'h2 == state ? writeBeatCnt_value : _GEN_43; // @[src/main/scala/nutcore/mem/Cache.scala 353:18 src/main/scala/chisel3/util/Counter.scala 61:40]
  wire [3:0] _GEN_50 = 4'h1 == state ? _GEN_29 : _GEN_48; // @[src/main/scala/nutcore/mem/Cache.scala 353:18]
  wire [2:0] _GEN_51 = 4'h1 == state ? _GEN_30 : _GEN_46; // @[src/main/scala/nutcore/mem/Cache.scala 353:18]
  wire  _GEN_52 = 4'h1 == state ? afterFirstRead : _GEN_45; // @[src/main/scala/nutcore/mem/Cache.scala 353:18 336:31]
  wire [2:0] _GEN_53 = 4'h1 == state ? _GEN_0 : _GEN_47; // @[src/main/scala/nutcore/mem/Cache.scala 353:18]
  wire [2:0] _GEN_54 = 4'h1 == state ? writeBeatCnt_value : _GEN_49; // @[src/main/scala/nutcore/mem/Cache.scala 353:18 src/main/scala/chisel3/util/Counter.scala 61:40]
  wire [2:0] _GEN_55 = 4'h8 == state ? _GEN_27 : _GEN_51; // @[src/main/scala/nutcore/mem/Cache.scala 353:18]
  wire [3:0] _GEN_56 = 4'h8 == state ? _GEN_28 : _GEN_50; // @[src/main/scala/nutcore/mem/Cache.scala 353:18]
  wire  _GEN_57 = 4'h8 == state ? afterFirstRead : _GEN_52; // @[src/main/scala/nutcore/mem/Cache.scala 353:18 336:31]
  wire [2:0] _GEN_58 = 4'h8 == state ? _GEN_0 : _GEN_53; // @[src/main/scala/nutcore/mem/Cache.scala 353:18]
  wire [2:0] _GEN_59 = 4'h8 == state ? writeBeatCnt_value : _GEN_54; // @[src/main/scala/nutcore/mem/Cache.scala 353:18 src/main/scala/chisel3/util/Counter.scala 61:40]
  wire [63:0] _dataRefill_T = readingFirst ? wordMask : 64'h0; // @[src/main/scala/nutcore/mem/Cache.scala 402:67]
  wire [63:0] _dataRefill_T_1 = io_in_bits_req_wdata & _dataRefill_T; // @[src/main/scala/utils/BitUtils.scala 34:14]
  wire [63:0] _dataRefill_T_2 = ~_dataRefill_T; // @[src/main/scala/utils/BitUtils.scala 34:39]
  wire [63:0] _dataRefill_T_3 = io_mem_resp_bits_rdata & _dataRefill_T_2; // @[src/main/scala/utils/BitUtils.scala 34:37]
  wire [63:0] dataRefill = _dataRefill_T_1 | _dataRefill_T_3; // @[src/main/scala/utils/BitUtils.scala 34:26]
  wire  dataRefillWriteBus_x9 = _readingFirst_T_3 & _readingFirst_T_1; // @[src/main/scala/nutcore/mem/Cache.scala 404:39]
  wire  metaRefillWriteBus_req_valid = dataRefillWriteBus_x9 & _T_57; // @[src/main/scala/nutcore/mem/Cache.scala 412:59]
  wire  _T_73 = dataRefillWriteBus_x9 & _hitReadBurst_T; // @[src/main/scala/nutcore/mem/Cache.scala 422:57]
  wire [2:0] _io_out_bits_cmd_T_1 = _T_57 ? 3'h6 : 3'h2; // @[src/main/scala/nutcore/mem/Cache.scala 425:29]
  wire [63:0] _io_out_bits_rdata_T = hit ? dataRead : inRdataRegDemand; // @[src/main/scala/nutcore/mem/Cache.scala 428:31]
  wire [2:0] _io_out_bits_cmd_T_2 = respToL1Last ? 3'h6 : 3'h2; // @[src/main/scala/nutcore/mem/Cache.scala 433:29]
  wire [63:0] _GEN_76 = hitReadBurst & _T_15 ? _dataHitWay_T_10 : _io_out_bits_rdata_T; // @[src/main/scala/nutcore/mem/Cache.scala 430:54 432:25 435:25]
  wire [3:0] _GEN_77 = hitReadBurst & _T_15 ? {{1'd0}, _io_out_bits_cmd_T_2} : io_in_bits_req_cmd; // @[src/main/scala/nutcore/mem/Cache.scala 430:54 433:23 436:23]
  wire [63:0] _GEN_78 = _T_7 | _T_6 ? _io_out_bits_rdata_T : _GEN_76; // @[src/main/scala/nutcore/mem/Cache.scala 426:75 428:25]
  wire  _io_out_valid_T_4 = state == 4'h7; // @[src/main/scala/nutcore/mem/Cache.scala 446:48]
  wire  _io_out_valid_T_17 = io_in_bits_req_cmd[0] & (hit | ~hit & state == 4'h7) | _T_73 | _T_50 & _T_15; // @[src/main/scala/nutcore/mem/Cache.scala 446:159]
  wire  _io_out_valid_T_23 = io_in_bits_req_cmd[0] | mmio ? _io_out_valid_T_4 : afterFirstRead & ~alreadyOutFire; // @[src/main/scala/nutcore/mem/Cache.scala 447:45]
  wire  _io_out_valid_T_25 = probe ? 1'h0 : hit | _io_out_valid_T_23; // @[src/main/scala/nutcore/mem/Cache.scala 447:8]
  wire  _io_out_valid_T_26 = io_in_bits_req_cmd[1] ? _io_out_valid_T_17 : _io_out_valid_T_25; // @[src/main/scala/nutcore/mem/Cache.scala 445:37]
  wire  _io_isFinish_T_4 = miss ? _io_cohResp_valid_T : _T_15 & releaseLast; // @[src/main/scala/nutcore/mem/Cache.scala 454:51]
  wire  _io_isFinish_T_13 = hit | io_in_bits_req_cmd[0] ? io_out_valid : _io_out_valid_T_4 & _GEN_12; // @[src/main/scala/nutcore/mem/Cache.scala 455:8]
  wire [255:0] _T_99 = {io_in_bits_datas_3_data,io_in_bits_datas_2_data,io_in_bits_datas_1_data,io_in_bits_datas_0_data}
    ; // @[src/main/scala/nutcore/mem/Cache.scala 464:465]
  reg [63:0] c; // @[src/main/scala/utils/GTimer.scala 24:20]
  wire [63:0] _c_T_1 = c + 64'h1; // @[src/main/scala/utils/GTimer.scala 25:12]
  reg [63:0] c_1; // @[src/main/scala/utils/GTimer.scala 24:20]
  wire [63:0] _c_T_3 = c_1 + 64'h1; // @[src/main/scala/utils/GTimer.scala 25:12]
  reg [63:0] c_2; // @[src/main/scala/utils/GTimer.scala 24:20]
  wire [63:0] _c_T_5 = c_2 + 64'h1; // @[src/main/scala/utils/GTimer.scala 25:12]
  wire  _T_106 = io_metaWriteBus_req_valid & DISPLAY_ENABLE; // @[src/main/scala/utils/Debug.scala 55:16]
  reg [63:0] c_3; // @[src/main/scala/utils/GTimer.scala 24:20]
  wire [63:0] _c_T_7 = c_3 + 64'h1; // @[src/main/scala/utils/GTimer.scala 25:12]
  reg [63:0] c_4; // @[src/main/scala/utils/GTimer.scala 24:20]
  wire [63:0] _c_T_9 = c_4 + 64'h1; // @[src/main/scala/utils/GTimer.scala 25:12]
  reg [63:0] c_5; // @[src/main/scala/utils/GTimer.scala 24:20]
  wire [63:0] _c_T_11 = c_5 + 64'h1; // @[src/main/scala/utils/GTimer.scala 25:12]
  reg [63:0] c_6; // @[src/main/scala/utils/GTimer.scala 24:20]
  wire [63:0] _c_T_13 = c_6 + 64'h1; // @[src/main/scala/utils/GTimer.scala 25:12]
  reg [63:0] c_7; // @[src/main/scala/utils/GTimer.scala 24:20]
  wire [63:0] _c_T_15 = c_7 + 64'h1; // @[src/main/scala/utils/GTimer.scala 25:12]
  reg [63:0] c_8; // @[src/main/scala/utils/GTimer.scala 24:20]
  wire [63:0] _c_T_17 = c_8 + 64'h1; // @[src/main/scala/utils/GTimer.scala 25:12]
  wire  _T_138 = io_dataWriteBus_req_valid & DISPLAY_ENABLE; // @[src/main/scala/utils/Debug.scala 55:16]
  wire  _T_145 = _T_14 & _T_26; // @[src/main/scala/nutcore/mem/Cache.scala 473:35]
  reg [63:0] c_9; // @[src/main/scala/utils/GTimer.scala 24:20]
  wire [63:0] _c_T_19 = c_9 + 64'h1; // @[src/main/scala/utils/GTimer.scala 25:12]
  wire  _T_150 = _T_145 & DISPLAY_ENABLE; // @[src/main/scala/utils/Debug.scala 55:16]
  wire  _T_157 = _cmd_T & _T_26; // @[src/main/scala/nutcore/mem/Cache.scala 474:34]
  reg [63:0] c_10; // @[src/main/scala/utils/GTimer.scala 24:20]
  wire [63:0] _c_T_21 = c_10 + 64'h1; // @[src/main/scala/utils/GTimer.scala 25:12]
  wire  _T_162 = _T_157 & DISPLAY_ENABLE; // @[src/main/scala/utils/Debug.scala 55:16]
  reg [63:0] c_11; // @[src/main/scala/utils/GTimer.scala 24:20]
  wire [63:0] _c_T_23 = c_11 + 64'h1; // @[src/main/scala/utils/GTimer.scala 25:12]
  wire  _T_174 = dataRefillWriteBus_x9 & DISPLAY_ENABLE; // @[src/main/scala/utils/Debug.scala 55:16]
  Arbiter_10 metaWriteArb ( // @[src/main/scala/nutcore/mem/Cache.scala 254:28]
    .io_in_0_valid(metaWriteArb_io_in_0_valid),
    .io_in_0_bits_setIdx(metaWriteArb_io_in_0_bits_setIdx),
    .io_in_0_bits_data_tag(metaWriteArb_io_in_0_bits_data_tag),
    .io_in_0_bits_waymask(metaWriteArb_io_in_0_bits_waymask),
    .io_in_1_valid(metaWriteArb_io_in_1_valid),
    .io_in_1_bits_setIdx(metaWriteArb_io_in_1_bits_setIdx),
    .io_in_1_bits_data_tag(metaWriteArb_io_in_1_bits_data_tag),
    .io_in_1_bits_data_dirty(metaWriteArb_io_in_1_bits_data_dirty),
    .io_in_1_bits_waymask(metaWriteArb_io_in_1_bits_waymask),
    .io_out_valid(metaWriteArb_io_out_valid),
    .io_out_bits_setIdx(metaWriteArb_io_out_bits_setIdx),
    .io_out_bits_data_tag(metaWriteArb_io_out_bits_data_tag),
    .io_out_bits_data_dirty(metaWriteArb_io_out_bits_data_dirty),
    .io_out_bits_waymask(metaWriteArb_io_out_bits_waymask)
  );
  Arbiter_11 dataWriteArb ( // @[src/main/scala/nutcore/mem/Cache.scala 255:28]
    .io_in_0_valid(dataWriteArb_io_in_0_valid),
    .io_in_0_bits_setIdx(dataWriteArb_io_in_0_bits_setIdx),
    .io_in_0_bits_data_data(dataWriteArb_io_in_0_bits_data_data),
    .io_in_0_bits_waymask(dataWriteArb_io_in_0_bits_waymask),
    .io_in_1_valid(dataWriteArb_io_in_1_valid),
    .io_in_1_bits_setIdx(dataWriteArb_io_in_1_bits_setIdx),
    .io_in_1_bits_data_data(dataWriteArb_io_in_1_bits_data_data),
    .io_in_1_bits_waymask(dataWriteArb_io_in_1_bits_waymask),
    .io_out_valid(dataWriteArb_io_out_valid),
    .io_out_bits_setIdx(dataWriteArb_io_out_bits_setIdx),
    .io_out_bits_data_data(dataWriteArb_io_out_bits_data_data),
    .io_out_bits_waymask(dataWriteArb_io_out_bits_waymask)
  );
  assign io_in_ready = _io_cohResp_valid_T & ~hitReadBurst & ~miss & ~probe; // @[src/main/scala/nutcore/mem/Cache.scala 458:79]
  assign io_out_valid = io_in_valid & _io_out_valid_T_26; // @[src/main/scala/nutcore/mem/Cache.scala 445:31]
  assign io_out_bits_cmd = dataRefillWriteBus_x9 & _hitReadBurst_T ? {{1'd0}, _io_out_bits_cmd_T_1} : _GEN_77; // @[src/main/scala/nutcore/mem/Cache.scala 422:79 425:23]
  assign io_out_bits_rdata = dataRefillWriteBus_x9 & _hitReadBurst_T ? dataRefill : _GEN_78; // @[src/main/scala/nutcore/mem/Cache.scala 422:79 424:25]
  assign io_isFinish = probe ? io_cohResp_valid & _io_isFinish_T_4 : _io_isFinish_T_13; // @[src/main/scala/nutcore/mem/Cache.scala 454:21]
  assign io_dataReadBus_req_valid = (state == 4'h3 | state == 4'h8) & state2 == 2'h0; // @[src/main/scala/nutcore/mem/Cache.scala 306:81]
  assign io_dataReadBus_req_bits_setIdx = {addr_index,_T_20}; // @[src/main/scala/nutcore/mem/Cache.scala 307:17]
  assign io_dataWriteBus_req_valid = dataWriteArb_io_out_valid; // @[src/main/scala/nutcore/mem/Cache.scala 409:23]
  assign io_dataWriteBus_req_bits_setIdx = dataWriteArb_io_out_bits_setIdx; // @[src/main/scala/nutcore/mem/Cache.scala 409:23]
  assign io_dataWriteBus_req_bits_data_data = dataWriteArb_io_out_bits_data_data; // @[src/main/scala/nutcore/mem/Cache.scala 409:23]
  assign io_dataWriteBus_req_bits_waymask = dataWriteArb_io_out_bits_waymask; // @[src/main/scala/nutcore/mem/Cache.scala 409:23]
  assign io_metaWriteBus_req_valid = metaWriteArb_io_out_valid; // @[src/main/scala/nutcore/mem/Cache.scala 419:23]
  assign io_metaWriteBus_req_bits_setIdx = metaWriteArb_io_out_bits_setIdx; // @[src/main/scala/nutcore/mem/Cache.scala 419:23]
  assign io_metaWriteBus_req_bits_data_tag = metaWriteArb_io_out_bits_data_tag; // @[src/main/scala/nutcore/mem/Cache.scala 419:23]
  assign io_metaWriteBus_req_bits_data_valid = 1'h1; // @[src/main/scala/nutcore/mem/Cache.scala 419:23]
  assign io_metaWriteBus_req_bits_data_dirty = metaWriteArb_io_out_bits_data_dirty; // @[src/main/scala/nutcore/mem/Cache.scala 419:23]
  assign io_metaWriteBus_req_bits_waymask = metaWriteArb_io_out_bits_waymask; // @[src/main/scala/nutcore/mem/Cache.scala 419:23]
  assign io_mem_req_valid = _cmd_T | _T_14 & state2 == 2'h2; // @[src/main/scala/nutcore/mem/Cache.scala 329:48]
  assign io_mem_req_bits_addr = _cmd_T ? raddr : waddr; // @[src/main/scala/nutcore/mem/Cache.scala 324:35]
  assign io_mem_req_bits_size = 3'h3; // @[src/main/scala/bus/simplebus/SimpleBus.scala 66:15]
  assign io_mem_req_bits_cmd = {{1'd0}, cmd}; // @[src/main/scala/bus/simplebus/SimpleBus.scala 65:14]
  assign io_mem_req_bits_wmask = 8'hff; // @[src/main/scala/nutcore/mem/Cache.scala 326:37]
  assign io_mem_req_bits_wdata = _dataHitWay_T_9 | _dataHitWay_T_7; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign io_mem_resp_ready = 1'h1; // @[src/main/scala/nutcore/mem/Cache.scala 328:21]
  assign io_cohResp_valid = state == 4'h0 & probe | _io_cohResp_valid_T_4; // @[src/main/scala/nutcore/mem/Cache.scala 343:53]
  assign io_dataReadRespToL1 = hitReadBurst & _respToL1Last_T_4; // @[src/main/scala/nutcore/mem/Cache.scala 459:39]
  assign metaWriteArb_io_in_0_valid = hitWrite & ~meta_dirty; // @[src/main/scala/nutcore/mem/Cache.scala 289:22]
  assign metaWriteArb_io_in_0_bits_setIdx = io_in_bits_req_addr[14:6]; // @[src/main/scala/nutcore/mem/Cache.scala 77:45]
  assign metaWriteArb_io_in_0_bits_data_tag = _meta_T_23 | _meta_T_21; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign metaWriteArb_io_in_0_bits_waymask = io_in_bits_waymask; // @[src/main/scala/nutcore/mem/Cache.scala 288:29 src/main/scala/utils/SRAMTemplate.scala 38:24]
  assign metaWriteArb_io_in_1_valid = dataRefillWriteBus_x9 & _T_57; // @[src/main/scala/nutcore/mem/Cache.scala 412:59]
  assign metaWriteArb_io_in_1_bits_setIdx = io_in_bits_req_addr[14:6]; // @[src/main/scala/nutcore/mem/Cache.scala 77:45]
  assign metaWriteArb_io_in_1_bits_data_tag = io_in_bits_req_addr[31:15]; // @[src/main/scala/nutcore/mem/Cache.scala 258:31]
  assign metaWriteArb_io_in_1_bits_data_dirty = io_in_bits_req_cmd[0]; // @[src/main/scala/bus/simplebus/SimpleBus.scala 74:22]
  assign metaWriteArb_io_in_1_bits_waymask = io_in_bits_waymask; // @[src/main/scala/nutcore/mem/Cache.scala 411:32 src/main/scala/utils/SRAMTemplate.scala 38:24]
  assign dataWriteArb_io_in_0_valid = hit & io_in_bits_req_cmd[0]; // @[src/main/scala/nutcore/mem/Cache.scala 283:22]
  assign dataWriteArb_io_in_0_bits_setIdx = {addr_index,_dataHitWriteBus_x3_T_3}; // @[src/main/scala/nutcore/mem/Cache.scala 286:35]
  assign dataWriteArb_io_in_0_bits_data_data = _dataHitWriteBus_x1_T | _dataHitWriteBus_x1_T_2; // @[src/main/scala/utils/BitUtils.scala 34:26]
  assign dataWriteArb_io_in_0_bits_waymask = io_in_bits_waymask; // @[src/main/scala/nutcore/mem/Cache.scala 284:29 src/main/scala/utils/SRAMTemplate.scala 38:24]
  assign dataWriteArb_io_in_1_valid = _readingFirst_T_3 & _readingFirst_T_1; // @[src/main/scala/nutcore/mem/Cache.scala 404:39]
  assign dataWriteArb_io_in_1_bits_setIdx = {addr_index,readBeatCnt_value}; // @[src/main/scala/nutcore/mem/Cache.scala 404:72]
  assign dataWriteArb_io_in_1_bits_data_data = _dataRefill_T_1 | _dataRefill_T_3; // @[src/main/scala/utils/BitUtils.scala 34:26]
  assign dataWriteArb_io_in_1_bits_waymask = io_in_bits_waymask; // @[src/main/scala/nutcore/mem/Cache.scala 403:32 src/main/scala/utils/SRAMTemplate.scala 38:24]
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/chisel3/util/Counter.scala 61:40]
      writeL2BeatCnt_value <= 3'h0; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end else if (4'h0 == state) begin // @[src/main/scala/nutcore/mem/Cache.scala 353:18]
      writeL2BeatCnt_value <= _GEN_0;
    end else if (4'h5 == state) begin // @[src/main/scala/nutcore/mem/Cache.scala 353:18]
      writeL2BeatCnt_value <= _GEN_0;
    end else if (4'h6 == state) begin // @[src/main/scala/nutcore/mem/Cache.scala 353:18]
      writeL2BeatCnt_value <= _GEN_0;
    end else begin
      writeL2BeatCnt_value <= _GEN_58;
    end
    if (reset) begin // @[src/main/scala/nutcore/mem/Cache.scala 294:22]
      state <= 4'h0; // @[src/main/scala/nutcore/mem/Cache.scala 294:22]
    end else if (4'h0 == state) begin // @[src/main/scala/nutcore/mem/Cache.scala 353:18]
      if (probe) begin // @[src/main/scala/nutcore/mem/Cache.scala 358:20]
        if (io_cohResp_valid) begin // @[src/main/scala/nutcore/mem/Cache.scala 359:32]
          state <= _state_T; // @[src/main/scala/nutcore/mem/Cache.scala 360:17]
        end
      end else if (hitReadBurst) begin // @[src/main/scala/nutcore/mem/Cache.scala 363:50]
        state <= 4'h8; // @[src/main/scala/nutcore/mem/Cache.scala 364:15]
      end else begin
        state <= _GEN_20;
      end
    end else if (!(4'h5 == state)) begin // @[src/main/scala/nutcore/mem/Cache.scala 353:18]
      if (!(4'h6 == state)) begin // @[src/main/scala/nutcore/mem/Cache.scala 353:18]
        state <= _GEN_56;
      end
    end
    if (reset) begin // @[src/main/scala/chisel3/util/Counter.scala 61:40]
      readBeatCnt_value <= 3'h0; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end else if (4'h0 == state) begin // @[src/main/scala/nutcore/mem/Cache.scala 353:18]
      if (probe) begin // @[src/main/scala/nutcore/mem/Cache.scala 358:20]
        if (io_cohResp_valid) begin // @[src/main/scala/nutcore/mem/Cache.scala 359:32]
          readBeatCnt_value <= addr_wordIndex; // @[src/main/scala/nutcore/mem/Cache.scala 361:29]
        end
      end else if (hitReadBurst) begin // @[src/main/scala/nutcore/mem/Cache.scala 363:50]
        readBeatCnt_value <= _value_T_5; // @[src/main/scala/nutcore/mem/Cache.scala 365:27]
      end
    end else if (!(4'h5 == state)) begin // @[src/main/scala/nutcore/mem/Cache.scala 353:18]
      if (!(4'h6 == state)) begin // @[src/main/scala/nutcore/mem/Cache.scala 353:18]
        readBeatCnt_value <= _GEN_55;
      end
    end
    if (reset) begin // @[src/main/scala/chisel3/util/Counter.scala 61:40]
      writeBeatCnt_value <= 3'h0; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end else if (!(4'h0 == state)) begin // @[src/main/scala/nutcore/mem/Cache.scala 353:18]
      if (!(4'h5 == state)) begin // @[src/main/scala/nutcore/mem/Cache.scala 353:18]
        if (!(4'h6 == state)) begin // @[src/main/scala/nutcore/mem/Cache.scala 353:18]
          writeBeatCnt_value <= _GEN_59;
        end
      end
    end
    if (reset) begin // @[src/main/scala/nutcore/mem/Cache.scala 304:23]
      state2 <= 2'h0; // @[src/main/scala/nutcore/mem/Cache.scala 304:23]
    end else if (2'h0 == state2) begin // @[src/main/scala/nutcore/mem/Cache.scala 311:19]
      if (_T_23) begin // @[src/main/scala/nutcore/mem/Cache.scala 312:51]
        state2 <= 2'h1; // @[src/main/scala/nutcore/mem/Cache.scala 312:60]
      end
    end else if (2'h1 == state2) begin // @[src/main/scala/nutcore/mem/Cache.scala 311:19]
      state2 <= 2'h2; // @[src/main/scala/nutcore/mem/Cache.scala 313:35]
    end else if (2'h2 == state2) begin // @[src/main/scala/nutcore/mem/Cache.scala 311:19]
      state2 <= _GEN_8;
    end
    if (state2 == 2'h1) begin // @[src/main/scala/nutcore/mem/Cache.scala 308:26]
      dataWay_0_data <= io_dataReadBus_resp_data_0_data; // @[src/main/scala/nutcore/mem/Cache.scala 308:26]
    end
    if (state2 == 2'h1) begin // @[src/main/scala/nutcore/mem/Cache.scala 308:26]
      dataWay_1_data <= io_dataReadBus_resp_data_1_data; // @[src/main/scala/nutcore/mem/Cache.scala 308:26]
    end
    if (state2 == 2'h1) begin // @[src/main/scala/nutcore/mem/Cache.scala 308:26]
      dataWay_2_data <= io_dataReadBus_resp_data_2_data; // @[src/main/scala/nutcore/mem/Cache.scala 308:26]
    end
    if (state2 == 2'h1) begin // @[src/main/scala/nutcore/mem/Cache.scala 308:26]
      dataWay_3_data <= io_dataReadBus_resp_data_3_data; // @[src/main/scala/nutcore/mem/Cache.scala 308:26]
    end
    if (reset) begin // @[src/main/scala/nutcore/mem/Cache.scala 336:31]
      afterFirstRead <= 1'h0; // @[src/main/scala/nutcore/mem/Cache.scala 336:31]
    end else if (4'h0 == state) begin // @[src/main/scala/nutcore/mem/Cache.scala 353:18]
      afterFirstRead <= 1'h0; // @[src/main/scala/nutcore/mem/Cache.scala 355:22]
    end else if (!(4'h5 == state)) begin // @[src/main/scala/nutcore/mem/Cache.scala 353:18]
      if (!(4'h6 == state)) begin // @[src/main/scala/nutcore/mem/Cache.scala 353:18]
        afterFirstRead <= _GEN_57;
      end
    end
    if (reset) begin // @[src/main/scala/nutcore/mem/Cache.scala 337:33]
      alreadyOutFire <= 1'h0; // @[src/main/scala/nutcore/mem/Cache.scala 337:33]
    end else if (4'h0 == state) begin // @[src/main/scala/nutcore/mem/Cache.scala 353:18]
      alreadyOutFire <= 1'h0; // @[src/main/scala/nutcore/mem/Cache.scala 356:22]
    end else begin
      alreadyOutFire <= _GEN_12;
    end
    if (_inRdataRegDemand_T_2) begin // @[src/main/scala/nutcore/mem/Cache.scala 339:35]
      if (mmio) begin // @[src/main/scala/nutcore/mem/Cache.scala 339:39]
        inRdataRegDemand <= 64'h0;
      end else begin
        inRdataRegDemand <= io_mem_resp_bits_rdata;
      end
    end
    if (reset) begin // @[src/main/scala/chisel3/util/Counter.scala 61:40]
      releaseLast_c_value <= 3'h0; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end else if (_releaseLast_T_2) begin // @[src/main/scala/chisel3/util/Counter.scala 118:16]
      releaseLast_c_value <= _releaseLast_wrap_value_T_1; // @[src/main/scala/chisel3/util/Counter.scala 77:15]
    end
    if (reset) begin // @[src/main/scala/chisel3/util/Counter.scala 61:40]
      respToL1Last_c_value <= 3'h0; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end else if (_respToL1Last_T_5) begin // @[src/main/scala/chisel3/util/Counter.scala 118:16]
      respToL1Last_c_value <= _respToL1Last_wrap_value_T_1; // @[src/main/scala/chisel3/util/Counter.scala 77:15]
    end
    if (reset) begin // @[src/main/scala/utils/GTimer.scala 24:20]
      c <= 64'h0; // @[src/main/scala/utils/GTimer.scala 24:20]
    end else begin
      c <= _c_T_1; // @[src/main/scala/utils/GTimer.scala 25:7]
    end
    if (reset) begin // @[src/main/scala/utils/GTimer.scala 24:20]
      c_1 <= 64'h0; // @[src/main/scala/utils/GTimer.scala 24:20]
    end else begin
      c_1 <= _c_T_3; // @[src/main/scala/utils/GTimer.scala 25:7]
    end
    if (reset) begin // @[src/main/scala/utils/GTimer.scala 24:20]
      c_2 <= 64'h0; // @[src/main/scala/utils/GTimer.scala 24:20]
    end else begin
      c_2 <= _c_T_5; // @[src/main/scala/utils/GTimer.scala 25:7]
    end
    if (reset) begin // @[src/main/scala/utils/GTimer.scala 24:20]
      c_3 <= 64'h0; // @[src/main/scala/utils/GTimer.scala 24:20]
    end else begin
      c_3 <= _c_T_7; // @[src/main/scala/utils/GTimer.scala 25:7]
    end
    if (reset) begin // @[src/main/scala/utils/GTimer.scala 24:20]
      c_4 <= 64'h0; // @[src/main/scala/utils/GTimer.scala 24:20]
    end else begin
      c_4 <= _c_T_9; // @[src/main/scala/utils/GTimer.scala 25:7]
    end
    if (reset) begin // @[src/main/scala/utils/GTimer.scala 24:20]
      c_5 <= 64'h0; // @[src/main/scala/utils/GTimer.scala 24:20]
    end else begin
      c_5 <= _c_T_11; // @[src/main/scala/utils/GTimer.scala 25:7]
    end
    if (reset) begin // @[src/main/scala/utils/GTimer.scala 24:20]
      c_6 <= 64'h0; // @[src/main/scala/utils/GTimer.scala 24:20]
    end else begin
      c_6 <= _c_T_13; // @[src/main/scala/utils/GTimer.scala 25:7]
    end
    if (reset) begin // @[src/main/scala/utils/GTimer.scala 24:20]
      c_7 <= 64'h0; // @[src/main/scala/utils/GTimer.scala 24:20]
    end else begin
      c_7 <= _c_T_15; // @[src/main/scala/utils/GTimer.scala 25:7]
    end
    if (reset) begin // @[src/main/scala/utils/GTimer.scala 24:20]
      c_8 <= 64'h0; // @[src/main/scala/utils/GTimer.scala 24:20]
    end else begin
      c_8 <= _c_T_17; // @[src/main/scala/utils/GTimer.scala 25:7]
    end
    if (reset) begin // @[src/main/scala/utils/GTimer.scala 24:20]
      c_9 <= 64'h0; // @[src/main/scala/utils/GTimer.scala 24:20]
    end else begin
      c_9 <= _c_T_19; // @[src/main/scala/utils/GTimer.scala 25:7]
    end
    if (reset) begin // @[src/main/scala/utils/GTimer.scala 24:20]
      c_10 <= 64'h0; // @[src/main/scala/utils/GTimer.scala 24:20]
    end else begin
      c_10 <= _c_T_21; // @[src/main/scala/utils/GTimer.scala 25:7]
    end
    if (reset) begin // @[src/main/scala/utils/GTimer.scala 24:20]
      c_11 <= 64'h0; // @[src/main/scala/utils/GTimer.scala 24:20]
    end else begin
      c_11 <= _c_T_23; // @[src/main/scala/utils/GTimer.scala 25:7]
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~(mmio & hit))) begin
          $fwrite(32'h80000002,
            "Assertion failed: MMIO request should not hit in cache\n    at Cache.scala:265 assert(!(mmio && hit), \"MMIO request should not hit in cache\")\n"
            ); // @[src/main/scala/nutcore/mem/Cache.scala 265:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~(mmio & hit)) & ~reset) begin
          $fatal; // @[src/main/scala/nutcore/mem/Cache.scala 265:9]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3 & ~(~(metaHitWriteBus_x5 & metaRefillWriteBus_req_valid))) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Cache.scala:461 assert(!(metaHitWriteBus.req.valid && metaRefillWriteBus.req.valid))\n"
            ); // @[src/main/scala/nutcore/mem/Cache.scala 461:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~(metaHitWriteBus_x5 & metaRefillWriteBus_req_valid)) & _T_3) begin
          $fatal; // @[src/main/scala/nutcore/mem/Cache.scala 461:9]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3 & ~(~(hitWrite & dataRefillWriteBus_x9))) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Cache.scala:462 assert(!(dataHitWriteBus.req.valid && dataRefillWriteBus.req.valid))\n"
            ); // @[src/main/scala/nutcore/mem/Cache.scala 462:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~(hitWrite & dataRefillWriteBus_x9)) & _T_3) begin
          $fatal; // @[src/main/scala/nutcore/mem/Cache.scala 462:9]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_3) begin
          $fwrite(32'h80000002,"[%d] CacheStage3_2: ",c); // @[src/main/scala/utils/Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_3) begin
          $fwrite(32'h80000002," metaread idx %x waymask %b metas %x%x:%x %x%x:%x %x%x:%x %x%x:%x %x\n",addr_index,
            io_in_bits_waymask,io_in_bits_metas_0_valid,io_in_bits_metas_0_dirty,io_in_bits_metas_0_tag,
            io_in_bits_metas_1_valid,io_in_bits_metas_1_dirty,io_in_bits_metas_1_tag,io_in_bits_metas_2_valid,
            io_in_bits_metas_2_dirty,io_in_bits_metas_2_tag,io_in_bits_metas_3_valid,io_in_bits_metas_3_dirty,
            io_in_bits_metas_3_tag,_T_99); // @[src/main/scala/utils/Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_106 & _T_3) begin
          $fwrite(32'h80000002,"[%d] CacheStage3_2: ",c_2); // @[src/main/scala/utils/Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_106 & _T_3) begin
          $fwrite(32'h80000002,"%d: [l2cache S3]: metawrite idx %x wmask %b meta %x%x:%x\n",c_1,
            io_metaWriteBus_req_bits_setIdx,io_metaWriteBus_req_bits_waymask,io_metaWriteBus_req_bits_data_valid,
            io_metaWriteBus_req_bits_data_dirty,io_metaWriteBus_req_bits_data_tag); // @[src/main/scala/utils/Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_3) begin
          $fwrite(32'h80000002,"[%d] CacheStage3_2: ",c_3); // @[src/main/scala/utils/Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_3) begin
          $fwrite(32'h80000002,
            " in.ready = %d, in.valid = %d, hit = %x, state = %d, addr = %x cmd:%d probe:%d isFinish:%d\n",io_in_ready,
            io_in_valid,hit,state,io_in_bits_req_addr,io_in_bits_req_cmd,probe,io_isFinish); // @[src/main/scala/utils/Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_3) begin
          $fwrite(32'h80000002,"[%d] CacheStage3_2: ",c_4); // @[src/main/scala/utils/Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_3) begin
          $fwrite(32'h80000002," out.valid:%d rdata:%x cmd:%d user:%x id:%x \n",io_out_valid,io_out_bits_rdata,
            io_out_bits_cmd,1'h0,1'h0); // @[src/main/scala/utils/Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_3) begin
          $fwrite(32'h80000002,"[%d] CacheStage3_2: ",c_5); // @[src/main/scala/utils/Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_3) begin
          $fwrite(32'h80000002," DHW: (%d, %d), data:%x setIdx:%x MHW:(%d, %d)\n",hitWrite,1'h1,dataHitWriteBus_x1_data,
            dataHitWriteBus_x3,metaHitWriteBus_x5,1'h1); // @[src/main/scala/utils/Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_3) begin
          $fwrite(32'h80000002,"[%d] CacheStage3_2: ",c_6); // @[src/main/scala/utils/Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_3) begin
          $fwrite(32'h80000002," DreadCache: %x \n",_T_99); // @[src/main/scala/utils/Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_3) begin
          $fwrite(32'h80000002,"[%d] CacheStage3_2: ",c_7); // @[src/main/scala/utils/Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_3) begin
          $fwrite(32'h80000002," useFD:%d isFD:%d FD:%x DreadArray:%x dataRead:%x inwaymask:%x FDwaymask:%x \n",
            useForwardData,io_in_bits_isForwardData,io_in_bits_forwardData_data_data,_dataReadArray_T_10,dataRead,
            io_in_bits_waymask,io_in_bits_forwardData_waymask); // @[src/main/scala/utils/Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_138 & _T_3) begin
          $fwrite(32'h80000002,"[%d] CacheStage3_2: ",c_8); // @[src/main/scala/utils/Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_138 & _T_3) begin
          $fwrite(32'h80000002,"[WB] waymask: %b data:%x setIdx:%x\n",io_dataWriteBus_req_bits_waymask,
            io_dataWriteBus_req_bits_data_data,io_dataWriteBus_req_bits_setIdx); // @[src/main/scala/utils/Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_150 & _T_3) begin
          $fwrite(32'h80000002,"[%d] CacheStage3_2: ",c_9); // @[src/main/scala/utils/Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_150 & _T_3) begin
          $fwrite(32'h80000002,"[COUTW] cnt %x addr %x data %x cmd %x size %x wmask %x tag %x idx %x waymask %b \n",
            writeBeatCnt_value,io_mem_req_bits_addr,io_mem_req_bits_wdata,io_mem_req_bits_cmd,io_mem_req_bits_size,
            io_mem_req_bits_wmask,addr_tag,addr_index,io_in_bits_waymask); // @[src/main/scala/utils/Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_162 & _T_3) begin
          $fwrite(32'h80000002,"[%d] CacheStage3_2: ",c_10); // @[src/main/scala/utils/Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_162 & _T_3) begin
          $fwrite(32'h80000002,"[COUTR] addr %x tag %x idx %x waymask %b \n",io_mem_req_bits_addr,addr_tag,addr_index,
            io_in_bits_waymask); // @[src/main/scala/utils/Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_174 & _T_3) begin
          $fwrite(32'h80000002,"[%d] CacheStage3_2: ",c_11); // @[src/main/scala/utils/Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_174 & _T_3) begin
          $fwrite(32'h80000002,"[COUTR] cnt %x data %x tag %x idx %x waymask %b \n",readBeatCnt_value,
            io_mem_resp_bits_rdata,addr_tag,addr_index,io_in_bits_waymask); // @[src/main/scala/utils/Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  writeL2BeatCnt_value = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  state = _RAND_1[3:0];
  _RAND_2 = {1{`RANDOM}};
  readBeatCnt_value = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  writeBeatCnt_value = _RAND_3[2:0];
  _RAND_4 = {1{`RANDOM}};
  state2 = _RAND_4[1:0];
  _RAND_5 = {2{`RANDOM}};
  dataWay_0_data = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  dataWay_1_data = _RAND_6[63:0];
  _RAND_7 = {2{`RANDOM}};
  dataWay_2_data = _RAND_7[63:0];
  _RAND_8 = {2{`RANDOM}};
  dataWay_3_data = _RAND_8[63:0];
  _RAND_9 = {1{`RANDOM}};
  afterFirstRead = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  alreadyOutFire = _RAND_10[0:0];
  _RAND_11 = {2{`RANDOM}};
  inRdataRegDemand = _RAND_11[63:0];
  _RAND_12 = {1{`RANDOM}};
  releaseLast_c_value = _RAND_12[2:0];
  _RAND_13 = {1{`RANDOM}};
  respToL1Last_c_value = _RAND_13[2:0];
  _RAND_14 = {2{`RANDOM}};
  c = _RAND_14[63:0];
  _RAND_15 = {2{`RANDOM}};
  c_1 = _RAND_15[63:0];
  _RAND_16 = {2{`RANDOM}};
  c_2 = _RAND_16[63:0];
  _RAND_17 = {2{`RANDOM}};
  c_3 = _RAND_17[63:0];
  _RAND_18 = {2{`RANDOM}};
  c_4 = _RAND_18[63:0];
  _RAND_19 = {2{`RANDOM}};
  c_5 = _RAND_19[63:0];
  _RAND_20 = {2{`RANDOM}};
  c_6 = _RAND_20[63:0];
  _RAND_21 = {2{`RANDOM}};
  c_7 = _RAND_21[63:0];
  _RAND_22 = {2{`RANDOM}};
  c_8 = _RAND_22[63:0];
  _RAND_23 = {2{`RANDOM}};
  c_9 = _RAND_23[63:0];
  _RAND_24 = {2{`RANDOM}};
  c_10 = _RAND_24[63:0];
  _RAND_25 = {2{`RANDOM}};
  c_11 = _RAND_25[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module SRAMTemplate_5(
  input         clock,
  input         reset,
  output        io_r_req_ready, // @[src/main/scala/utils/SRAMTemplate.scala 70:14]
  input         io_r_req_valid, // @[src/main/scala/utils/SRAMTemplate.scala 70:14]
  input  [8:0]  io_r_req_bits_setIdx, // @[src/main/scala/utils/SRAMTemplate.scala 70:14]
  output [16:0] io_r_resp_data_0_tag, // @[src/main/scala/utils/SRAMTemplate.scala 70:14]
  output        io_r_resp_data_0_valid, // @[src/main/scala/utils/SRAMTemplate.scala 70:14]
  output        io_r_resp_data_0_dirty, // @[src/main/scala/utils/SRAMTemplate.scala 70:14]
  output [16:0] io_r_resp_data_1_tag, // @[src/main/scala/utils/SRAMTemplate.scala 70:14]
  output        io_r_resp_data_1_valid, // @[src/main/scala/utils/SRAMTemplate.scala 70:14]
  output        io_r_resp_data_1_dirty, // @[src/main/scala/utils/SRAMTemplate.scala 70:14]
  output [16:0] io_r_resp_data_2_tag, // @[src/main/scala/utils/SRAMTemplate.scala 70:14]
  output        io_r_resp_data_2_valid, // @[src/main/scala/utils/SRAMTemplate.scala 70:14]
  output        io_r_resp_data_2_dirty, // @[src/main/scala/utils/SRAMTemplate.scala 70:14]
  output [16:0] io_r_resp_data_3_tag, // @[src/main/scala/utils/SRAMTemplate.scala 70:14]
  output        io_r_resp_data_3_valid, // @[src/main/scala/utils/SRAMTemplate.scala 70:14]
  output        io_r_resp_data_3_dirty, // @[src/main/scala/utils/SRAMTemplate.scala 70:14]
  input         io_w_req_valid, // @[src/main/scala/utils/SRAMTemplate.scala 70:14]
  input  [8:0]  io_w_req_bits_setIdx, // @[src/main/scala/utils/SRAMTemplate.scala 70:14]
  input  [16:0] io_w_req_bits_data_tag, // @[src/main/scala/utils/SRAMTemplate.scala 70:14]
  input         io_w_req_bits_data_dirty, // @[src/main/scala/utils/SRAMTemplate.scala 70:14]
  input  [3:0]  io_w_req_bits_waymask // @[src/main/scala/utils/SRAMTemplate.scala 70:14]
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_9;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
`endif // RANDOMIZE_REG_INIT
  reg [18:0] array_0 [0:511]; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
  wire  array_0_rdata_MPORT_en; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
  wire [8:0] array_0_rdata_MPORT_addr; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
  wire [18:0] array_0_rdata_MPORT_data; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
  wire [18:0] array_0_MPORT_data; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
  wire [8:0] array_0_MPORT_addr; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
  wire  array_0_MPORT_mask; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
  wire  array_0_MPORT_en; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
  reg  array_0_rdata_MPORT_en_pipe_0;
  reg [8:0] array_0_rdata_MPORT_addr_pipe_0;
  reg [18:0] array_1 [0:511]; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
  wire  array_1_rdata_MPORT_en; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
  wire [8:0] array_1_rdata_MPORT_addr; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
  wire [18:0] array_1_rdata_MPORT_data; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
  wire [18:0] array_1_MPORT_data; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
  wire [8:0] array_1_MPORT_addr; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
  wire  array_1_MPORT_mask; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
  wire  array_1_MPORT_en; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
  reg  array_1_rdata_MPORT_en_pipe_0;
  reg [8:0] array_1_rdata_MPORT_addr_pipe_0;
  reg [18:0] array_2 [0:511]; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
  wire  array_2_rdata_MPORT_en; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
  wire [8:0] array_2_rdata_MPORT_addr; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
  wire [18:0] array_2_rdata_MPORT_data; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
  wire [18:0] array_2_MPORT_data; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
  wire [8:0] array_2_MPORT_addr; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
  wire  array_2_MPORT_mask; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
  wire  array_2_MPORT_en; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
  reg  array_2_rdata_MPORT_en_pipe_0;
  reg [8:0] array_2_rdata_MPORT_addr_pipe_0;
  reg [18:0] array_3 [0:511]; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
  wire  array_3_rdata_MPORT_en; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
  wire [8:0] array_3_rdata_MPORT_addr; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
  wire [18:0] array_3_rdata_MPORT_data; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
  wire [18:0] array_3_MPORT_data; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
  wire [8:0] array_3_MPORT_addr; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
  wire  array_3_MPORT_mask; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
  wire  array_3_MPORT_en; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
  reg  array_3_rdata_MPORT_en_pipe_0;
  reg [8:0] array_3_rdata_MPORT_addr_pipe_0;
  reg  resetState; // @[src/main/scala/utils/SRAMTemplate.scala 80:30]
  reg [8:0] resetSet; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
  wire  wrap_wrap = resetSet == 9'h1ff; // @[src/main/scala/chisel3/util/Counter.scala 73:24]
  wire [8:0] _wrap_value_T_1 = resetSet + 9'h1; // @[src/main/scala/chisel3/util/Counter.scala 77:24]
  wire  resetFinish = resetState & wrap_wrap; // @[src/main/scala/chisel3/util/Counter.scala 118:{16,23} 117:24]
  wire  _GEN_2 = resetFinish ? 1'h0 : resetState; // @[src/main/scala/utils/SRAMTemplate.scala 82:24 80:30 82:38]
  wire  wen = io_w_req_valid | resetState; // @[src/main/scala/utils/SRAMTemplate.scala 88:52]
  wire  _realRen_T = ~wen; // @[src/main/scala/utils/SRAMTemplate.scala 89:41]
  wire [18:0] _wdataword_T = {io_w_req_bits_data_tag,1'h1,io_w_req_bits_data_dirty}; // @[src/main/scala/utils/SRAMTemplate.scala 92:78]
  wire [3:0] waymask = resetState ? 4'hf : io_w_req_bits_waymask; // @[src/main/scala/utils/SRAMTemplate.scala 93:20]
  wire [18:0] _rdata_WIRE_1 = array_0_rdata_MPORT_data; // @[src/main/scala/utils/SRAMTemplate.scala 98:{78,78}]
  wire [18:0] _rdata_WIRE_2 = array_1_rdata_MPORT_data; // @[src/main/scala/utils/SRAMTemplate.scala 98:{78,78}]
  wire [18:0] _rdata_WIRE_3 = array_2_rdata_MPORT_data; // @[src/main/scala/utils/SRAMTemplate.scala 98:{78,78}]
  wire [18:0] _rdata_WIRE_4 = array_3_rdata_MPORT_data; // @[src/main/scala/utils/SRAMTemplate.scala 98:{78,78}]
  assign array_0_rdata_MPORT_en = array_0_rdata_MPORT_en_pipe_0;
  assign array_0_rdata_MPORT_addr = array_0_rdata_MPORT_addr_pipe_0;
  assign array_0_rdata_MPORT_data = array_0[array_0_rdata_MPORT_addr]; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
  assign array_0_MPORT_data = resetState ? 19'h0 : _wdataword_T;
  assign array_0_MPORT_addr = resetState ? resetSet : io_w_req_bits_setIdx;
  assign array_0_MPORT_mask = waymask[0];
  assign array_0_MPORT_en = io_w_req_valid | resetState;
  assign array_1_rdata_MPORT_en = array_1_rdata_MPORT_en_pipe_0;
  assign array_1_rdata_MPORT_addr = array_1_rdata_MPORT_addr_pipe_0;
  assign array_1_rdata_MPORT_data = array_1[array_1_rdata_MPORT_addr]; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
  assign array_1_MPORT_data = resetState ? 19'h0 : _wdataword_T;
  assign array_1_MPORT_addr = resetState ? resetSet : io_w_req_bits_setIdx;
  assign array_1_MPORT_mask = waymask[1];
  assign array_1_MPORT_en = io_w_req_valid | resetState;
  assign array_2_rdata_MPORT_en = array_2_rdata_MPORT_en_pipe_0;
  assign array_2_rdata_MPORT_addr = array_2_rdata_MPORT_addr_pipe_0;
  assign array_2_rdata_MPORT_data = array_2[array_2_rdata_MPORT_addr]; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
  assign array_2_MPORT_data = resetState ? 19'h0 : _wdataword_T;
  assign array_2_MPORT_addr = resetState ? resetSet : io_w_req_bits_setIdx;
  assign array_2_MPORT_mask = waymask[2];
  assign array_2_MPORT_en = io_w_req_valid | resetState;
  assign array_3_rdata_MPORT_en = array_3_rdata_MPORT_en_pipe_0;
  assign array_3_rdata_MPORT_addr = array_3_rdata_MPORT_addr_pipe_0;
  assign array_3_rdata_MPORT_data = array_3[array_3_rdata_MPORT_addr]; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
  assign array_3_MPORT_data = resetState ? 19'h0 : _wdataword_T;
  assign array_3_MPORT_addr = resetState ? resetSet : io_w_req_bits_setIdx;
  assign array_3_MPORT_mask = waymask[3];
  assign array_3_MPORT_en = io_w_req_valid | resetState;
  assign io_r_req_ready = ~resetState & _realRen_T; // @[src/main/scala/utils/SRAMTemplate.scala 101:33]
  assign io_r_resp_data_0_tag = _rdata_WIRE_1[18:2]; // @[src/main/scala/utils/SRAMTemplate.scala 98:78]
  assign io_r_resp_data_0_valid = _rdata_WIRE_1[1]; // @[src/main/scala/utils/SRAMTemplate.scala 98:78]
  assign io_r_resp_data_0_dirty = _rdata_WIRE_1[0]; // @[src/main/scala/utils/SRAMTemplate.scala 98:78]
  assign io_r_resp_data_1_tag = _rdata_WIRE_2[18:2]; // @[src/main/scala/utils/SRAMTemplate.scala 98:78]
  assign io_r_resp_data_1_valid = _rdata_WIRE_2[1]; // @[src/main/scala/utils/SRAMTemplate.scala 98:78]
  assign io_r_resp_data_1_dirty = _rdata_WIRE_2[0]; // @[src/main/scala/utils/SRAMTemplate.scala 98:78]
  assign io_r_resp_data_2_tag = _rdata_WIRE_3[18:2]; // @[src/main/scala/utils/SRAMTemplate.scala 98:78]
  assign io_r_resp_data_2_valid = _rdata_WIRE_3[1]; // @[src/main/scala/utils/SRAMTemplate.scala 98:78]
  assign io_r_resp_data_2_dirty = _rdata_WIRE_3[0]; // @[src/main/scala/utils/SRAMTemplate.scala 98:78]
  assign io_r_resp_data_3_tag = _rdata_WIRE_4[18:2]; // @[src/main/scala/utils/SRAMTemplate.scala 98:78]
  assign io_r_resp_data_3_valid = _rdata_WIRE_4[1]; // @[src/main/scala/utils/SRAMTemplate.scala 98:78]
  assign io_r_resp_data_3_dirty = _rdata_WIRE_4[0]; // @[src/main/scala/utils/SRAMTemplate.scala 98:78]
  always @(posedge clock) begin
    if (array_0_MPORT_en & array_0_MPORT_mask) begin
      array_0[array_0_MPORT_addr] <= array_0_MPORT_data; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
    end
    array_0_rdata_MPORT_en_pipe_0 <= io_r_req_valid & _realRen_T;
    if (io_r_req_valid & _realRen_T) begin
      array_0_rdata_MPORT_addr_pipe_0 <= io_r_req_bits_setIdx;
    end
    if (array_1_MPORT_en & array_1_MPORT_mask) begin
      array_1[array_1_MPORT_addr] <= array_1_MPORT_data; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
    end
    array_1_rdata_MPORT_en_pipe_0 <= io_r_req_valid & _realRen_T;
    if (io_r_req_valid & _realRen_T) begin
      array_1_rdata_MPORT_addr_pipe_0 <= io_r_req_bits_setIdx;
    end
    if (array_2_MPORT_en & array_2_MPORT_mask) begin
      array_2[array_2_MPORT_addr] <= array_2_MPORT_data; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
    end
    array_2_rdata_MPORT_en_pipe_0 <= io_r_req_valid & _realRen_T;
    if (io_r_req_valid & _realRen_T) begin
      array_2_rdata_MPORT_addr_pipe_0 <= io_r_req_bits_setIdx;
    end
    if (array_3_MPORT_en & array_3_MPORT_mask) begin
      array_3[array_3_MPORT_addr] <= array_3_MPORT_data; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
    end
    array_3_rdata_MPORT_en_pipe_0 <= io_r_req_valid & _realRen_T;
    if (io_r_req_valid & _realRen_T) begin
      array_3_rdata_MPORT_addr_pipe_0 <= io_r_req_bits_setIdx;
    end
    resetState <= reset | _GEN_2; // @[src/main/scala/utils/SRAMTemplate.scala 80:{30,30}]
    if (reset) begin // @[src/main/scala/chisel3/util/Counter.scala 61:40]
      resetSet <= 9'h0; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end else if (resetState) begin // @[src/main/scala/chisel3/util/Counter.scala 118:16]
      resetSet <= _wrap_value_T_1; // @[src/main/scala/chisel3/util/Counter.scala 77:15]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    array_0[initvar] = _RAND_0[18:0];
  _RAND_3 = {1{`RANDOM}};
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    array_1[initvar] = _RAND_3[18:0];
  _RAND_6 = {1{`RANDOM}};
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    array_2[initvar] = _RAND_6[18:0];
  _RAND_9 = {1{`RANDOM}};
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    array_3[initvar] = _RAND_9[18:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  array_0_rdata_MPORT_en_pipe_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  array_0_rdata_MPORT_addr_pipe_0 = _RAND_2[8:0];
  _RAND_4 = {1{`RANDOM}};
  array_1_rdata_MPORT_en_pipe_0 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  array_1_rdata_MPORT_addr_pipe_0 = _RAND_5[8:0];
  _RAND_7 = {1{`RANDOM}};
  array_2_rdata_MPORT_en_pipe_0 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  array_2_rdata_MPORT_addr_pipe_0 = _RAND_8[8:0];
  _RAND_10 = {1{`RANDOM}};
  array_3_rdata_MPORT_en_pipe_0 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  array_3_rdata_MPORT_addr_pipe_0 = _RAND_11[8:0];
  _RAND_12 = {1{`RANDOM}};
  resetState = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  resetSet = _RAND_13[8:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Arbiter_12(
  output       io_in_0_ready, // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
  input        io_in_0_valid, // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
  input  [8:0] io_in_0_bits_setIdx, // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
  input        io_out_ready, // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
  output       io_out_valid, // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
  output [8:0] io_out_bits_setIdx // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
);
  assign io_in_0_ready = io_out_ready; // @[src/main/scala/chisel3/util/Arbiter.scala 147:19]
  assign io_out_valid = io_in_0_valid; // @[src/main/scala/chisel3/util/Arbiter.scala 148:31]
  assign io_out_bits_setIdx = io_in_0_bits_setIdx; // @[src/main/scala/chisel3/util/Arbiter.scala 137:15]
endmodule
module SRAMTemplateWithArbiter_4(
  input         clock,
  input         reset,
  output        io_r_0_req_ready, // @[src/main/scala/utils/SRAMTemplate.scala 116:14]
  input         io_r_0_req_valid, // @[src/main/scala/utils/SRAMTemplate.scala 116:14]
  input  [8:0]  io_r_0_req_bits_setIdx, // @[src/main/scala/utils/SRAMTemplate.scala 116:14]
  output [16:0] io_r_0_resp_data_0_tag, // @[src/main/scala/utils/SRAMTemplate.scala 116:14]
  output        io_r_0_resp_data_0_valid, // @[src/main/scala/utils/SRAMTemplate.scala 116:14]
  output        io_r_0_resp_data_0_dirty, // @[src/main/scala/utils/SRAMTemplate.scala 116:14]
  output [16:0] io_r_0_resp_data_1_tag, // @[src/main/scala/utils/SRAMTemplate.scala 116:14]
  output        io_r_0_resp_data_1_valid, // @[src/main/scala/utils/SRAMTemplate.scala 116:14]
  output        io_r_0_resp_data_1_dirty, // @[src/main/scala/utils/SRAMTemplate.scala 116:14]
  output [16:0] io_r_0_resp_data_2_tag, // @[src/main/scala/utils/SRAMTemplate.scala 116:14]
  output        io_r_0_resp_data_2_valid, // @[src/main/scala/utils/SRAMTemplate.scala 116:14]
  output        io_r_0_resp_data_2_dirty, // @[src/main/scala/utils/SRAMTemplate.scala 116:14]
  output [16:0] io_r_0_resp_data_3_tag, // @[src/main/scala/utils/SRAMTemplate.scala 116:14]
  output        io_r_0_resp_data_3_valid, // @[src/main/scala/utils/SRAMTemplate.scala 116:14]
  output        io_r_0_resp_data_3_dirty, // @[src/main/scala/utils/SRAMTemplate.scala 116:14]
  input         io_w_req_valid, // @[src/main/scala/utils/SRAMTemplate.scala 116:14]
  input  [8:0]  io_w_req_bits_setIdx, // @[src/main/scala/utils/SRAMTemplate.scala 116:14]
  input  [16:0] io_w_req_bits_data_tag, // @[src/main/scala/utils/SRAMTemplate.scala 116:14]
  input         io_w_req_bits_data_dirty, // @[src/main/scala/utils/SRAMTemplate.scala 116:14]
  input  [3:0]  io_w_req_bits_waymask // @[src/main/scala/utils/SRAMTemplate.scala 116:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
`endif // RANDOMIZE_REG_INIT
  wire  ram_clock; // @[src/main/scala/utils/SRAMTemplate.scala 121:19]
  wire  ram_reset; // @[src/main/scala/utils/SRAMTemplate.scala 121:19]
  wire  ram_io_r_req_ready; // @[src/main/scala/utils/SRAMTemplate.scala 121:19]
  wire  ram_io_r_req_valid; // @[src/main/scala/utils/SRAMTemplate.scala 121:19]
  wire [8:0] ram_io_r_req_bits_setIdx; // @[src/main/scala/utils/SRAMTemplate.scala 121:19]
  wire [16:0] ram_io_r_resp_data_0_tag; // @[src/main/scala/utils/SRAMTemplate.scala 121:19]
  wire  ram_io_r_resp_data_0_valid; // @[src/main/scala/utils/SRAMTemplate.scala 121:19]
  wire  ram_io_r_resp_data_0_dirty; // @[src/main/scala/utils/SRAMTemplate.scala 121:19]
  wire [16:0] ram_io_r_resp_data_1_tag; // @[src/main/scala/utils/SRAMTemplate.scala 121:19]
  wire  ram_io_r_resp_data_1_valid; // @[src/main/scala/utils/SRAMTemplate.scala 121:19]
  wire  ram_io_r_resp_data_1_dirty; // @[src/main/scala/utils/SRAMTemplate.scala 121:19]
  wire [16:0] ram_io_r_resp_data_2_tag; // @[src/main/scala/utils/SRAMTemplate.scala 121:19]
  wire  ram_io_r_resp_data_2_valid; // @[src/main/scala/utils/SRAMTemplate.scala 121:19]
  wire  ram_io_r_resp_data_2_dirty; // @[src/main/scala/utils/SRAMTemplate.scala 121:19]
  wire [16:0] ram_io_r_resp_data_3_tag; // @[src/main/scala/utils/SRAMTemplate.scala 121:19]
  wire  ram_io_r_resp_data_3_valid; // @[src/main/scala/utils/SRAMTemplate.scala 121:19]
  wire  ram_io_r_resp_data_3_dirty; // @[src/main/scala/utils/SRAMTemplate.scala 121:19]
  wire  ram_io_w_req_valid; // @[src/main/scala/utils/SRAMTemplate.scala 121:19]
  wire [8:0] ram_io_w_req_bits_setIdx; // @[src/main/scala/utils/SRAMTemplate.scala 121:19]
  wire [16:0] ram_io_w_req_bits_data_tag; // @[src/main/scala/utils/SRAMTemplate.scala 121:19]
  wire  ram_io_w_req_bits_data_dirty; // @[src/main/scala/utils/SRAMTemplate.scala 121:19]
  wire [3:0] ram_io_w_req_bits_waymask; // @[src/main/scala/utils/SRAMTemplate.scala 121:19]
  wire  readArb_io_in_0_ready; // @[src/main/scala/utils/SRAMTemplate.scala 124:23]
  wire  readArb_io_in_0_valid; // @[src/main/scala/utils/SRAMTemplate.scala 124:23]
  wire [8:0] readArb_io_in_0_bits_setIdx; // @[src/main/scala/utils/SRAMTemplate.scala 124:23]
  wire  readArb_io_out_ready; // @[src/main/scala/utils/SRAMTemplate.scala 124:23]
  wire  readArb_io_out_valid; // @[src/main/scala/utils/SRAMTemplate.scala 124:23]
  wire [8:0] readArb_io_out_bits_setIdx; // @[src/main/scala/utils/SRAMTemplate.scala 124:23]
  reg  REG; // @[src/main/scala/utils/SRAMTemplate.scala 130:58]
  reg [16:0] r_0_tag; // @[src/main/scala/utils/Hold.scala 23:65]
  reg  r_0_valid; // @[src/main/scala/utils/Hold.scala 23:65]
  reg  r_0_dirty; // @[src/main/scala/utils/Hold.scala 23:65]
  reg [16:0] r_1_tag; // @[src/main/scala/utils/Hold.scala 23:65]
  reg  r_1_valid; // @[src/main/scala/utils/Hold.scala 23:65]
  reg  r_1_dirty; // @[src/main/scala/utils/Hold.scala 23:65]
  reg [16:0] r_2_tag; // @[src/main/scala/utils/Hold.scala 23:65]
  reg  r_2_valid; // @[src/main/scala/utils/Hold.scala 23:65]
  reg  r_2_dirty; // @[src/main/scala/utils/Hold.scala 23:65]
  reg [16:0] r_3_tag; // @[src/main/scala/utils/Hold.scala 23:65]
  reg  r_3_valid; // @[src/main/scala/utils/Hold.scala 23:65]
  reg  r_3_dirty; // @[src/main/scala/utils/Hold.scala 23:65]
  SRAMTemplate_5 ram ( // @[src/main/scala/utils/SRAMTemplate.scala 121:19]
    .clock(ram_clock),
    .reset(ram_reset),
    .io_r_req_ready(ram_io_r_req_ready),
    .io_r_req_valid(ram_io_r_req_valid),
    .io_r_req_bits_setIdx(ram_io_r_req_bits_setIdx),
    .io_r_resp_data_0_tag(ram_io_r_resp_data_0_tag),
    .io_r_resp_data_0_valid(ram_io_r_resp_data_0_valid),
    .io_r_resp_data_0_dirty(ram_io_r_resp_data_0_dirty),
    .io_r_resp_data_1_tag(ram_io_r_resp_data_1_tag),
    .io_r_resp_data_1_valid(ram_io_r_resp_data_1_valid),
    .io_r_resp_data_1_dirty(ram_io_r_resp_data_1_dirty),
    .io_r_resp_data_2_tag(ram_io_r_resp_data_2_tag),
    .io_r_resp_data_2_valid(ram_io_r_resp_data_2_valid),
    .io_r_resp_data_2_dirty(ram_io_r_resp_data_2_dirty),
    .io_r_resp_data_3_tag(ram_io_r_resp_data_3_tag),
    .io_r_resp_data_3_valid(ram_io_r_resp_data_3_valid),
    .io_r_resp_data_3_dirty(ram_io_r_resp_data_3_dirty),
    .io_w_req_valid(ram_io_w_req_valid),
    .io_w_req_bits_setIdx(ram_io_w_req_bits_setIdx),
    .io_w_req_bits_data_tag(ram_io_w_req_bits_data_tag),
    .io_w_req_bits_data_dirty(ram_io_w_req_bits_data_dirty),
    .io_w_req_bits_waymask(ram_io_w_req_bits_waymask)
  );
  Arbiter_12 readArb ( // @[src/main/scala/utils/SRAMTemplate.scala 124:23]
    .io_in_0_ready(readArb_io_in_0_ready),
    .io_in_0_valid(readArb_io_in_0_valid),
    .io_in_0_bits_setIdx(readArb_io_in_0_bits_setIdx),
    .io_out_ready(readArb_io_out_ready),
    .io_out_valid(readArb_io_out_valid),
    .io_out_bits_setIdx(readArb_io_out_bits_setIdx)
  );
  assign io_r_0_req_ready = readArb_io_in_0_ready; // @[src/main/scala/utils/SRAMTemplate.scala 125:17]
  assign io_r_0_resp_data_0_tag = REG ? ram_io_r_resp_data_0_tag : r_0_tag; // @[src/main/scala/utils/Hold.scala 23:48]
  assign io_r_0_resp_data_0_valid = REG ? ram_io_r_resp_data_0_valid : r_0_valid; // @[src/main/scala/utils/Hold.scala 23:48]
  assign io_r_0_resp_data_0_dirty = REG ? ram_io_r_resp_data_0_dirty : r_0_dirty; // @[src/main/scala/utils/Hold.scala 23:48]
  assign io_r_0_resp_data_1_tag = REG ? ram_io_r_resp_data_1_tag : r_1_tag; // @[src/main/scala/utils/Hold.scala 23:48]
  assign io_r_0_resp_data_1_valid = REG ? ram_io_r_resp_data_1_valid : r_1_valid; // @[src/main/scala/utils/Hold.scala 23:48]
  assign io_r_0_resp_data_1_dirty = REG ? ram_io_r_resp_data_1_dirty : r_1_dirty; // @[src/main/scala/utils/Hold.scala 23:48]
  assign io_r_0_resp_data_2_tag = REG ? ram_io_r_resp_data_2_tag : r_2_tag; // @[src/main/scala/utils/Hold.scala 23:48]
  assign io_r_0_resp_data_2_valid = REG ? ram_io_r_resp_data_2_valid : r_2_valid; // @[src/main/scala/utils/Hold.scala 23:48]
  assign io_r_0_resp_data_2_dirty = REG ? ram_io_r_resp_data_2_dirty : r_2_dirty; // @[src/main/scala/utils/Hold.scala 23:48]
  assign io_r_0_resp_data_3_tag = REG ? ram_io_r_resp_data_3_tag : r_3_tag; // @[src/main/scala/utils/Hold.scala 23:48]
  assign io_r_0_resp_data_3_valid = REG ? ram_io_r_resp_data_3_valid : r_3_valid; // @[src/main/scala/utils/Hold.scala 23:48]
  assign io_r_0_resp_data_3_dirty = REG ? ram_io_r_resp_data_3_dirty : r_3_dirty; // @[src/main/scala/utils/Hold.scala 23:48]
  assign ram_clock = clock;
  assign ram_reset = reset;
  assign ram_io_r_req_valid = readArb_io_out_valid; // @[src/main/scala/utils/SRAMTemplate.scala 126:16]
  assign ram_io_r_req_bits_setIdx = readArb_io_out_bits_setIdx; // @[src/main/scala/utils/SRAMTemplate.scala 126:16]
  assign ram_io_w_req_valid = io_w_req_valid; // @[src/main/scala/utils/SRAMTemplate.scala 122:12]
  assign ram_io_w_req_bits_setIdx = io_w_req_bits_setIdx; // @[src/main/scala/utils/SRAMTemplate.scala 122:12]
  assign ram_io_w_req_bits_data_tag = io_w_req_bits_data_tag; // @[src/main/scala/utils/SRAMTemplate.scala 122:12]
  assign ram_io_w_req_bits_data_dirty = io_w_req_bits_data_dirty; // @[src/main/scala/utils/SRAMTemplate.scala 122:12]
  assign ram_io_w_req_bits_waymask = io_w_req_bits_waymask; // @[src/main/scala/utils/SRAMTemplate.scala 122:12]
  assign readArb_io_in_0_valid = io_r_0_req_valid; // @[src/main/scala/utils/SRAMTemplate.scala 125:17]
  assign readArb_io_in_0_bits_setIdx = io_r_0_req_bits_setIdx; // @[src/main/scala/utils/SRAMTemplate.scala 125:17]
  assign readArb_io_out_ready = ram_io_r_req_ready; // @[src/main/scala/utils/SRAMTemplate.scala 126:16]
  always @(posedge clock) begin
    REG <= io_r_0_req_ready & io_r_0_req_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
    if (reset) begin // @[src/main/scala/utils/Hold.scala 23:65]
      r_0_tag <= 17'h0; // @[src/main/scala/utils/Hold.scala 23:65]
    end else if (REG) begin // @[src/main/scala/utils/Hold.scala 23:65]
      r_0_tag <= ram_io_r_resp_data_0_tag; // @[src/main/scala/utils/Hold.scala 23:65]
    end
    if (reset) begin // @[src/main/scala/utils/Hold.scala 23:65]
      r_0_valid <= 1'h0; // @[src/main/scala/utils/Hold.scala 23:65]
    end else if (REG) begin // @[src/main/scala/utils/Hold.scala 23:65]
      r_0_valid <= ram_io_r_resp_data_0_valid; // @[src/main/scala/utils/Hold.scala 23:65]
    end
    if (reset) begin // @[src/main/scala/utils/Hold.scala 23:65]
      r_0_dirty <= 1'h0; // @[src/main/scala/utils/Hold.scala 23:65]
    end else if (REG) begin // @[src/main/scala/utils/Hold.scala 23:65]
      r_0_dirty <= ram_io_r_resp_data_0_dirty; // @[src/main/scala/utils/Hold.scala 23:65]
    end
    if (reset) begin // @[src/main/scala/utils/Hold.scala 23:65]
      r_1_tag <= 17'h0; // @[src/main/scala/utils/Hold.scala 23:65]
    end else if (REG) begin // @[src/main/scala/utils/Hold.scala 23:65]
      r_1_tag <= ram_io_r_resp_data_1_tag; // @[src/main/scala/utils/Hold.scala 23:65]
    end
    if (reset) begin // @[src/main/scala/utils/Hold.scala 23:65]
      r_1_valid <= 1'h0; // @[src/main/scala/utils/Hold.scala 23:65]
    end else if (REG) begin // @[src/main/scala/utils/Hold.scala 23:65]
      r_1_valid <= ram_io_r_resp_data_1_valid; // @[src/main/scala/utils/Hold.scala 23:65]
    end
    if (reset) begin // @[src/main/scala/utils/Hold.scala 23:65]
      r_1_dirty <= 1'h0; // @[src/main/scala/utils/Hold.scala 23:65]
    end else if (REG) begin // @[src/main/scala/utils/Hold.scala 23:65]
      r_1_dirty <= ram_io_r_resp_data_1_dirty; // @[src/main/scala/utils/Hold.scala 23:65]
    end
    if (reset) begin // @[src/main/scala/utils/Hold.scala 23:65]
      r_2_tag <= 17'h0; // @[src/main/scala/utils/Hold.scala 23:65]
    end else if (REG) begin // @[src/main/scala/utils/Hold.scala 23:65]
      r_2_tag <= ram_io_r_resp_data_2_tag; // @[src/main/scala/utils/Hold.scala 23:65]
    end
    if (reset) begin // @[src/main/scala/utils/Hold.scala 23:65]
      r_2_valid <= 1'h0; // @[src/main/scala/utils/Hold.scala 23:65]
    end else if (REG) begin // @[src/main/scala/utils/Hold.scala 23:65]
      r_2_valid <= ram_io_r_resp_data_2_valid; // @[src/main/scala/utils/Hold.scala 23:65]
    end
    if (reset) begin // @[src/main/scala/utils/Hold.scala 23:65]
      r_2_dirty <= 1'h0; // @[src/main/scala/utils/Hold.scala 23:65]
    end else if (REG) begin // @[src/main/scala/utils/Hold.scala 23:65]
      r_2_dirty <= ram_io_r_resp_data_2_dirty; // @[src/main/scala/utils/Hold.scala 23:65]
    end
    if (reset) begin // @[src/main/scala/utils/Hold.scala 23:65]
      r_3_tag <= 17'h0; // @[src/main/scala/utils/Hold.scala 23:65]
    end else if (REG) begin // @[src/main/scala/utils/Hold.scala 23:65]
      r_3_tag <= ram_io_r_resp_data_3_tag; // @[src/main/scala/utils/Hold.scala 23:65]
    end
    if (reset) begin // @[src/main/scala/utils/Hold.scala 23:65]
      r_3_valid <= 1'h0; // @[src/main/scala/utils/Hold.scala 23:65]
    end else if (REG) begin // @[src/main/scala/utils/Hold.scala 23:65]
      r_3_valid <= ram_io_r_resp_data_3_valid; // @[src/main/scala/utils/Hold.scala 23:65]
    end
    if (reset) begin // @[src/main/scala/utils/Hold.scala 23:65]
      r_3_dirty <= 1'h0; // @[src/main/scala/utils/Hold.scala 23:65]
    end else if (REG) begin // @[src/main/scala/utils/Hold.scala 23:65]
      r_3_dirty <= ram_io_r_resp_data_3_dirty; // @[src/main/scala/utils/Hold.scala 23:65]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  REG = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  r_0_tag = _RAND_1[16:0];
  _RAND_2 = {1{`RANDOM}};
  r_0_valid = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  r_0_dirty = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  r_1_tag = _RAND_4[16:0];
  _RAND_5 = {1{`RANDOM}};
  r_1_valid = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  r_1_dirty = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  r_2_tag = _RAND_7[16:0];
  _RAND_8 = {1{`RANDOM}};
  r_2_valid = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  r_2_dirty = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  r_3_tag = _RAND_10[16:0];
  _RAND_11 = {1{`RANDOM}};
  r_3_valid = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  r_3_dirty = _RAND_12[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module SRAMTemplate_6(
  input         clock,
  output        io_r_req_ready, // @[src/main/scala/utils/SRAMTemplate.scala 70:14]
  input         io_r_req_valid, // @[src/main/scala/utils/SRAMTemplate.scala 70:14]
  input  [11:0] io_r_req_bits_setIdx, // @[src/main/scala/utils/SRAMTemplate.scala 70:14]
  output [63:0] io_r_resp_data_0_data, // @[src/main/scala/utils/SRAMTemplate.scala 70:14]
  output [63:0] io_r_resp_data_1_data, // @[src/main/scala/utils/SRAMTemplate.scala 70:14]
  output [63:0] io_r_resp_data_2_data, // @[src/main/scala/utils/SRAMTemplate.scala 70:14]
  output [63:0] io_r_resp_data_3_data, // @[src/main/scala/utils/SRAMTemplate.scala 70:14]
  input         io_w_req_valid, // @[src/main/scala/utils/SRAMTemplate.scala 70:14]
  input  [11:0] io_w_req_bits_setIdx, // @[src/main/scala/utils/SRAMTemplate.scala 70:14]
  input  [63:0] io_w_req_bits_data_data, // @[src/main/scala/utils/SRAMTemplate.scala 70:14]
  input  [3:0]  io_w_req_bits_waymask // @[src/main/scala/utils/SRAMTemplate.scala 70:14]
);
`ifdef RANDOMIZE_MEM_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_9;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
`endif // RANDOMIZE_REG_INIT
  reg [63:0] array_0 [0:4095]; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
  wire  array_0_rdata_MPORT_en; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
  wire [11:0] array_0_rdata_MPORT_addr; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
  wire [63:0] array_0_rdata_MPORT_data; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
  wire [63:0] array_0_MPORT_data; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
  wire [11:0] array_0_MPORT_addr; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
  wire  array_0_MPORT_mask; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
  wire  array_0_MPORT_en; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
  reg  array_0_rdata_MPORT_en_pipe_0;
  reg [11:0] array_0_rdata_MPORT_addr_pipe_0;
  reg [63:0] array_1 [0:4095]; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
  wire  array_1_rdata_MPORT_en; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
  wire [11:0] array_1_rdata_MPORT_addr; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
  wire [63:0] array_1_rdata_MPORT_data; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
  wire [63:0] array_1_MPORT_data; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
  wire [11:0] array_1_MPORT_addr; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
  wire  array_1_MPORT_mask; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
  wire  array_1_MPORT_en; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
  reg  array_1_rdata_MPORT_en_pipe_0;
  reg [11:0] array_1_rdata_MPORT_addr_pipe_0;
  reg [63:0] array_2 [0:4095]; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
  wire  array_2_rdata_MPORT_en; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
  wire [11:0] array_2_rdata_MPORT_addr; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
  wire [63:0] array_2_rdata_MPORT_data; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
  wire [63:0] array_2_MPORT_data; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
  wire [11:0] array_2_MPORT_addr; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
  wire  array_2_MPORT_mask; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
  wire  array_2_MPORT_en; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
  reg  array_2_rdata_MPORT_en_pipe_0;
  reg [11:0] array_2_rdata_MPORT_addr_pipe_0;
  reg [63:0] array_3 [0:4095]; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
  wire  array_3_rdata_MPORT_en; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
  wire [11:0] array_3_rdata_MPORT_addr; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
  wire [63:0] array_3_rdata_MPORT_data; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
  wire [63:0] array_3_MPORT_data; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
  wire [11:0] array_3_MPORT_addr; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
  wire  array_3_MPORT_mask; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
  wire  array_3_MPORT_en; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
  reg  array_3_rdata_MPORT_en_pipe_0;
  reg [11:0] array_3_rdata_MPORT_addr_pipe_0;
  wire  _realRen_T = ~io_w_req_valid; // @[src/main/scala/utils/SRAMTemplate.scala 89:41]
  assign array_0_rdata_MPORT_en = array_0_rdata_MPORT_en_pipe_0;
  assign array_0_rdata_MPORT_addr = array_0_rdata_MPORT_addr_pipe_0;
  assign array_0_rdata_MPORT_data = array_0[array_0_rdata_MPORT_addr]; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
  assign array_0_MPORT_data = io_w_req_bits_data_data;
  assign array_0_MPORT_addr = io_w_req_bits_setIdx;
  assign array_0_MPORT_mask = io_w_req_bits_waymask[0];
  assign array_0_MPORT_en = io_w_req_valid;
  assign array_1_rdata_MPORT_en = array_1_rdata_MPORT_en_pipe_0;
  assign array_1_rdata_MPORT_addr = array_1_rdata_MPORT_addr_pipe_0;
  assign array_1_rdata_MPORT_data = array_1[array_1_rdata_MPORT_addr]; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
  assign array_1_MPORT_data = io_w_req_bits_data_data;
  assign array_1_MPORT_addr = io_w_req_bits_setIdx;
  assign array_1_MPORT_mask = io_w_req_bits_waymask[1];
  assign array_1_MPORT_en = io_w_req_valid;
  assign array_2_rdata_MPORT_en = array_2_rdata_MPORT_en_pipe_0;
  assign array_2_rdata_MPORT_addr = array_2_rdata_MPORT_addr_pipe_0;
  assign array_2_rdata_MPORT_data = array_2[array_2_rdata_MPORT_addr]; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
  assign array_2_MPORT_data = io_w_req_bits_data_data;
  assign array_2_MPORT_addr = io_w_req_bits_setIdx;
  assign array_2_MPORT_mask = io_w_req_bits_waymask[2];
  assign array_2_MPORT_en = io_w_req_valid;
  assign array_3_rdata_MPORT_en = array_3_rdata_MPORT_en_pipe_0;
  assign array_3_rdata_MPORT_addr = array_3_rdata_MPORT_addr_pipe_0;
  assign array_3_rdata_MPORT_data = array_3[array_3_rdata_MPORT_addr]; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
  assign array_3_MPORT_data = io_w_req_bits_data_data;
  assign array_3_MPORT_addr = io_w_req_bits_setIdx;
  assign array_3_MPORT_mask = io_w_req_bits_waymask[3];
  assign array_3_MPORT_en = io_w_req_valid;
  assign io_r_req_ready = ~io_w_req_valid; // @[src/main/scala/utils/SRAMTemplate.scala 101:53]
  assign io_r_resp_data_0_data = array_0_rdata_MPORT_data; // @[src/main/scala/utils/SRAMTemplate.scala 98:{78,78}]
  assign io_r_resp_data_1_data = array_1_rdata_MPORT_data; // @[src/main/scala/utils/SRAMTemplate.scala 98:{78,78}]
  assign io_r_resp_data_2_data = array_2_rdata_MPORT_data; // @[src/main/scala/utils/SRAMTemplate.scala 98:{78,78}]
  assign io_r_resp_data_3_data = array_3_rdata_MPORT_data; // @[src/main/scala/utils/SRAMTemplate.scala 98:{78,78}]
  always @(posedge clock) begin
    if (array_0_MPORT_en & array_0_MPORT_mask) begin
      array_0[array_0_MPORT_addr] <= array_0_MPORT_data; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
    end
    array_0_rdata_MPORT_en_pipe_0 <= io_r_req_valid & _realRen_T;
    if (io_r_req_valid & _realRen_T) begin
      array_0_rdata_MPORT_addr_pipe_0 <= io_r_req_bits_setIdx;
    end
    if (array_1_MPORT_en & array_1_MPORT_mask) begin
      array_1[array_1_MPORT_addr] <= array_1_MPORT_data; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
    end
    array_1_rdata_MPORT_en_pipe_0 <= io_r_req_valid & _realRen_T;
    if (io_r_req_valid & _realRen_T) begin
      array_1_rdata_MPORT_addr_pipe_0 <= io_r_req_bits_setIdx;
    end
    if (array_2_MPORT_en & array_2_MPORT_mask) begin
      array_2[array_2_MPORT_addr] <= array_2_MPORT_data; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
    end
    array_2_rdata_MPORT_en_pipe_0 <= io_r_req_valid & _realRen_T;
    if (io_r_req_valid & _realRen_T) begin
      array_2_rdata_MPORT_addr_pipe_0 <= io_r_req_bits_setIdx;
    end
    if (array_3_MPORT_en & array_3_MPORT_mask) begin
      array_3[array_3_MPORT_addr] <= array_3_MPORT_data; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
    end
    array_3_rdata_MPORT_en_pipe_0 <= io_r_req_valid & _realRen_T;
    if (io_r_req_valid & _realRen_T) begin
      array_3_rdata_MPORT_addr_pipe_0 <= io_r_req_bits_setIdx;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {2{`RANDOM}};
  for (initvar = 0; initvar < 4096; initvar = initvar+1)
    array_0[initvar] = _RAND_0[63:0];
  _RAND_3 = {2{`RANDOM}};
  for (initvar = 0; initvar < 4096; initvar = initvar+1)
    array_1[initvar] = _RAND_3[63:0];
  _RAND_6 = {2{`RANDOM}};
  for (initvar = 0; initvar < 4096; initvar = initvar+1)
    array_2[initvar] = _RAND_6[63:0];
  _RAND_9 = {2{`RANDOM}};
  for (initvar = 0; initvar < 4096; initvar = initvar+1)
    array_3[initvar] = _RAND_9[63:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  array_0_rdata_MPORT_en_pipe_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  array_0_rdata_MPORT_addr_pipe_0 = _RAND_2[11:0];
  _RAND_4 = {1{`RANDOM}};
  array_1_rdata_MPORT_en_pipe_0 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  array_1_rdata_MPORT_addr_pipe_0 = _RAND_5[11:0];
  _RAND_7 = {1{`RANDOM}};
  array_2_rdata_MPORT_en_pipe_0 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  array_2_rdata_MPORT_addr_pipe_0 = _RAND_8[11:0];
  _RAND_10 = {1{`RANDOM}};
  array_3_rdata_MPORT_en_pipe_0 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  array_3_rdata_MPORT_addr_pipe_0 = _RAND_11[11:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Arbiter_13(
  output        io_in_0_ready, // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
  input         io_in_0_valid, // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
  input  [11:0] io_in_0_bits_setIdx, // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
  output        io_in_1_ready, // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
  input         io_in_1_valid, // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
  input  [11:0] io_in_1_bits_setIdx, // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
  input         io_out_ready, // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
  output        io_out_valid, // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
  output [11:0] io_out_bits_setIdx // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
);
  wire  grant_1 = ~io_in_0_valid; // @[src/main/scala/chisel3/util/Arbiter.scala 45:78]
  assign io_in_0_ready = io_out_ready; // @[src/main/scala/chisel3/util/Arbiter.scala 147:19]
  assign io_in_1_ready = grant_1 & io_out_ready; // @[src/main/scala/chisel3/util/Arbiter.scala 147:19]
  assign io_out_valid = ~grant_1 | io_in_1_valid; // @[src/main/scala/chisel3/util/Arbiter.scala 148:31]
  assign io_out_bits_setIdx = io_in_0_valid ? io_in_0_bits_setIdx : io_in_1_bits_setIdx; // @[src/main/scala/chisel3/util/Arbiter.scala 137:15 139:26 141:19]
endmodule
module SRAMTemplateWithArbiter_5(
  input         clock,
  input         reset,
  output        io_r_0_req_ready, // @[src/main/scala/utils/SRAMTemplate.scala 116:14]
  input         io_r_0_req_valid, // @[src/main/scala/utils/SRAMTemplate.scala 116:14]
  input  [11:0] io_r_0_req_bits_setIdx, // @[src/main/scala/utils/SRAMTemplate.scala 116:14]
  output [63:0] io_r_0_resp_data_0_data, // @[src/main/scala/utils/SRAMTemplate.scala 116:14]
  output [63:0] io_r_0_resp_data_1_data, // @[src/main/scala/utils/SRAMTemplate.scala 116:14]
  output [63:0] io_r_0_resp_data_2_data, // @[src/main/scala/utils/SRAMTemplate.scala 116:14]
  output [63:0] io_r_0_resp_data_3_data, // @[src/main/scala/utils/SRAMTemplate.scala 116:14]
  output        io_r_1_req_ready, // @[src/main/scala/utils/SRAMTemplate.scala 116:14]
  input         io_r_1_req_valid, // @[src/main/scala/utils/SRAMTemplate.scala 116:14]
  input  [11:0] io_r_1_req_bits_setIdx, // @[src/main/scala/utils/SRAMTemplate.scala 116:14]
  output [63:0] io_r_1_resp_data_0_data, // @[src/main/scala/utils/SRAMTemplate.scala 116:14]
  output [63:0] io_r_1_resp_data_1_data, // @[src/main/scala/utils/SRAMTemplate.scala 116:14]
  output [63:0] io_r_1_resp_data_2_data, // @[src/main/scala/utils/SRAMTemplate.scala 116:14]
  output [63:0] io_r_1_resp_data_3_data, // @[src/main/scala/utils/SRAMTemplate.scala 116:14]
  input         io_w_req_valid, // @[src/main/scala/utils/SRAMTemplate.scala 116:14]
  input  [11:0] io_w_req_bits_setIdx, // @[src/main/scala/utils/SRAMTemplate.scala 116:14]
  input  [63:0] io_w_req_bits_data_data, // @[src/main/scala/utils/SRAMTemplate.scala 116:14]
  input  [3:0]  io_w_req_bits_waymask // @[src/main/scala/utils/SRAMTemplate.scala 116:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [63:0] _RAND_9;
`endif // RANDOMIZE_REG_INIT
  wire  ram_clock; // @[src/main/scala/utils/SRAMTemplate.scala 121:19]
  wire  ram_io_r_req_ready; // @[src/main/scala/utils/SRAMTemplate.scala 121:19]
  wire  ram_io_r_req_valid; // @[src/main/scala/utils/SRAMTemplate.scala 121:19]
  wire [11:0] ram_io_r_req_bits_setIdx; // @[src/main/scala/utils/SRAMTemplate.scala 121:19]
  wire [63:0] ram_io_r_resp_data_0_data; // @[src/main/scala/utils/SRAMTemplate.scala 121:19]
  wire [63:0] ram_io_r_resp_data_1_data; // @[src/main/scala/utils/SRAMTemplate.scala 121:19]
  wire [63:0] ram_io_r_resp_data_2_data; // @[src/main/scala/utils/SRAMTemplate.scala 121:19]
  wire [63:0] ram_io_r_resp_data_3_data; // @[src/main/scala/utils/SRAMTemplate.scala 121:19]
  wire  ram_io_w_req_valid; // @[src/main/scala/utils/SRAMTemplate.scala 121:19]
  wire [11:0] ram_io_w_req_bits_setIdx; // @[src/main/scala/utils/SRAMTemplate.scala 121:19]
  wire [63:0] ram_io_w_req_bits_data_data; // @[src/main/scala/utils/SRAMTemplate.scala 121:19]
  wire [3:0] ram_io_w_req_bits_waymask; // @[src/main/scala/utils/SRAMTemplate.scala 121:19]
  wire  readArb_io_in_0_ready; // @[src/main/scala/utils/SRAMTemplate.scala 124:23]
  wire  readArb_io_in_0_valid; // @[src/main/scala/utils/SRAMTemplate.scala 124:23]
  wire [11:0] readArb_io_in_0_bits_setIdx; // @[src/main/scala/utils/SRAMTemplate.scala 124:23]
  wire  readArb_io_in_1_ready; // @[src/main/scala/utils/SRAMTemplate.scala 124:23]
  wire  readArb_io_in_1_valid; // @[src/main/scala/utils/SRAMTemplate.scala 124:23]
  wire [11:0] readArb_io_in_1_bits_setIdx; // @[src/main/scala/utils/SRAMTemplate.scala 124:23]
  wire  readArb_io_out_ready; // @[src/main/scala/utils/SRAMTemplate.scala 124:23]
  wire  readArb_io_out_valid; // @[src/main/scala/utils/SRAMTemplate.scala 124:23]
  wire [11:0] readArb_io_out_bits_setIdx; // @[src/main/scala/utils/SRAMTemplate.scala 124:23]
  reg  REG; // @[src/main/scala/utils/SRAMTemplate.scala 130:58]
  reg [63:0] r__0_data; // @[src/main/scala/utils/Hold.scala 23:65]
  reg [63:0] r__1_data; // @[src/main/scala/utils/Hold.scala 23:65]
  reg [63:0] r__2_data; // @[src/main/scala/utils/Hold.scala 23:65]
  reg [63:0] r__3_data; // @[src/main/scala/utils/Hold.scala 23:65]
  reg  REG_1; // @[src/main/scala/utils/SRAMTemplate.scala 130:58]
  reg [63:0] r_1_0_data; // @[src/main/scala/utils/Hold.scala 23:65]
  reg [63:0] r_1_1_data; // @[src/main/scala/utils/Hold.scala 23:65]
  reg [63:0] r_1_2_data; // @[src/main/scala/utils/Hold.scala 23:65]
  reg [63:0] r_1_3_data; // @[src/main/scala/utils/Hold.scala 23:65]
  SRAMTemplate_6 ram ( // @[src/main/scala/utils/SRAMTemplate.scala 121:19]
    .clock(ram_clock),
    .io_r_req_ready(ram_io_r_req_ready),
    .io_r_req_valid(ram_io_r_req_valid),
    .io_r_req_bits_setIdx(ram_io_r_req_bits_setIdx),
    .io_r_resp_data_0_data(ram_io_r_resp_data_0_data),
    .io_r_resp_data_1_data(ram_io_r_resp_data_1_data),
    .io_r_resp_data_2_data(ram_io_r_resp_data_2_data),
    .io_r_resp_data_3_data(ram_io_r_resp_data_3_data),
    .io_w_req_valid(ram_io_w_req_valid),
    .io_w_req_bits_setIdx(ram_io_w_req_bits_setIdx),
    .io_w_req_bits_data_data(ram_io_w_req_bits_data_data),
    .io_w_req_bits_waymask(ram_io_w_req_bits_waymask)
  );
  Arbiter_13 readArb ( // @[src/main/scala/utils/SRAMTemplate.scala 124:23]
    .io_in_0_ready(readArb_io_in_0_ready),
    .io_in_0_valid(readArb_io_in_0_valid),
    .io_in_0_bits_setIdx(readArb_io_in_0_bits_setIdx),
    .io_in_1_ready(readArb_io_in_1_ready),
    .io_in_1_valid(readArb_io_in_1_valid),
    .io_in_1_bits_setIdx(readArb_io_in_1_bits_setIdx),
    .io_out_ready(readArb_io_out_ready),
    .io_out_valid(readArb_io_out_valid),
    .io_out_bits_setIdx(readArb_io_out_bits_setIdx)
  );
  assign io_r_0_req_ready = readArb_io_in_0_ready; // @[src/main/scala/utils/SRAMTemplate.scala 125:17]
  assign io_r_0_resp_data_0_data = REG ? ram_io_r_resp_data_0_data : r__0_data; // @[src/main/scala/utils/Hold.scala 23:48]
  assign io_r_0_resp_data_1_data = REG ? ram_io_r_resp_data_1_data : r__1_data; // @[src/main/scala/utils/Hold.scala 23:48]
  assign io_r_0_resp_data_2_data = REG ? ram_io_r_resp_data_2_data : r__2_data; // @[src/main/scala/utils/Hold.scala 23:48]
  assign io_r_0_resp_data_3_data = REG ? ram_io_r_resp_data_3_data : r__3_data; // @[src/main/scala/utils/Hold.scala 23:48]
  assign io_r_1_req_ready = readArb_io_in_1_ready; // @[src/main/scala/utils/SRAMTemplate.scala 125:17]
  assign io_r_1_resp_data_0_data = REG_1 ? ram_io_r_resp_data_0_data : r_1_0_data; // @[src/main/scala/utils/Hold.scala 23:48]
  assign io_r_1_resp_data_1_data = REG_1 ? ram_io_r_resp_data_1_data : r_1_1_data; // @[src/main/scala/utils/Hold.scala 23:48]
  assign io_r_1_resp_data_2_data = REG_1 ? ram_io_r_resp_data_2_data : r_1_2_data; // @[src/main/scala/utils/Hold.scala 23:48]
  assign io_r_1_resp_data_3_data = REG_1 ? ram_io_r_resp_data_3_data : r_1_3_data; // @[src/main/scala/utils/Hold.scala 23:48]
  assign ram_clock = clock;
  assign ram_io_r_req_valid = readArb_io_out_valid; // @[src/main/scala/utils/SRAMTemplate.scala 126:16]
  assign ram_io_r_req_bits_setIdx = readArb_io_out_bits_setIdx; // @[src/main/scala/utils/SRAMTemplate.scala 126:16]
  assign ram_io_w_req_valid = io_w_req_valid; // @[src/main/scala/utils/SRAMTemplate.scala 122:12]
  assign ram_io_w_req_bits_setIdx = io_w_req_bits_setIdx; // @[src/main/scala/utils/SRAMTemplate.scala 122:12]
  assign ram_io_w_req_bits_data_data = io_w_req_bits_data_data; // @[src/main/scala/utils/SRAMTemplate.scala 122:12]
  assign ram_io_w_req_bits_waymask = io_w_req_bits_waymask; // @[src/main/scala/utils/SRAMTemplate.scala 122:12]
  assign readArb_io_in_0_valid = io_r_0_req_valid; // @[src/main/scala/utils/SRAMTemplate.scala 125:17]
  assign readArb_io_in_0_bits_setIdx = io_r_0_req_bits_setIdx; // @[src/main/scala/utils/SRAMTemplate.scala 125:17]
  assign readArb_io_in_1_valid = io_r_1_req_valid; // @[src/main/scala/utils/SRAMTemplate.scala 125:17]
  assign readArb_io_in_1_bits_setIdx = io_r_1_req_bits_setIdx; // @[src/main/scala/utils/SRAMTemplate.scala 125:17]
  assign readArb_io_out_ready = ram_io_r_req_ready; // @[src/main/scala/utils/SRAMTemplate.scala 126:16]
  always @(posedge clock) begin
    REG <= io_r_0_req_ready & io_r_0_req_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
    if (reset) begin // @[src/main/scala/utils/Hold.scala 23:65]
      r__0_data <= 64'h0; // @[src/main/scala/utils/Hold.scala 23:65]
    end else if (REG) begin // @[src/main/scala/utils/Hold.scala 23:65]
      r__0_data <= ram_io_r_resp_data_0_data; // @[src/main/scala/utils/Hold.scala 23:65]
    end
    if (reset) begin // @[src/main/scala/utils/Hold.scala 23:65]
      r__1_data <= 64'h0; // @[src/main/scala/utils/Hold.scala 23:65]
    end else if (REG) begin // @[src/main/scala/utils/Hold.scala 23:65]
      r__1_data <= ram_io_r_resp_data_1_data; // @[src/main/scala/utils/Hold.scala 23:65]
    end
    if (reset) begin // @[src/main/scala/utils/Hold.scala 23:65]
      r__2_data <= 64'h0; // @[src/main/scala/utils/Hold.scala 23:65]
    end else if (REG) begin // @[src/main/scala/utils/Hold.scala 23:65]
      r__2_data <= ram_io_r_resp_data_2_data; // @[src/main/scala/utils/Hold.scala 23:65]
    end
    if (reset) begin // @[src/main/scala/utils/Hold.scala 23:65]
      r__3_data <= 64'h0; // @[src/main/scala/utils/Hold.scala 23:65]
    end else if (REG) begin // @[src/main/scala/utils/Hold.scala 23:65]
      r__3_data <= ram_io_r_resp_data_3_data; // @[src/main/scala/utils/Hold.scala 23:65]
    end
    REG_1 <= io_r_1_req_ready & io_r_1_req_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
    if (reset) begin // @[src/main/scala/utils/Hold.scala 23:65]
      r_1_0_data <= 64'h0; // @[src/main/scala/utils/Hold.scala 23:65]
    end else if (REG_1) begin // @[src/main/scala/utils/Hold.scala 23:65]
      r_1_0_data <= ram_io_r_resp_data_0_data; // @[src/main/scala/utils/Hold.scala 23:65]
    end
    if (reset) begin // @[src/main/scala/utils/Hold.scala 23:65]
      r_1_1_data <= 64'h0; // @[src/main/scala/utils/Hold.scala 23:65]
    end else if (REG_1) begin // @[src/main/scala/utils/Hold.scala 23:65]
      r_1_1_data <= ram_io_r_resp_data_1_data; // @[src/main/scala/utils/Hold.scala 23:65]
    end
    if (reset) begin // @[src/main/scala/utils/Hold.scala 23:65]
      r_1_2_data <= 64'h0; // @[src/main/scala/utils/Hold.scala 23:65]
    end else if (REG_1) begin // @[src/main/scala/utils/Hold.scala 23:65]
      r_1_2_data <= ram_io_r_resp_data_2_data; // @[src/main/scala/utils/Hold.scala 23:65]
    end
    if (reset) begin // @[src/main/scala/utils/Hold.scala 23:65]
      r_1_3_data <= 64'h0; // @[src/main/scala/utils/Hold.scala 23:65]
    end else if (REG_1) begin // @[src/main/scala/utils/Hold.scala 23:65]
      r_1_3_data <= ram_io_r_resp_data_3_data; // @[src/main/scala/utils/Hold.scala 23:65]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  REG = _RAND_0[0:0];
  _RAND_1 = {2{`RANDOM}};
  r__0_data = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  r__1_data = _RAND_2[63:0];
  _RAND_3 = {2{`RANDOM}};
  r__2_data = _RAND_3[63:0];
  _RAND_4 = {2{`RANDOM}};
  r__3_data = _RAND_4[63:0];
  _RAND_5 = {1{`RANDOM}};
  REG_1 = _RAND_5[0:0];
  _RAND_6 = {2{`RANDOM}};
  r_1_0_data = _RAND_6[63:0];
  _RAND_7 = {2{`RANDOM}};
  r_1_1_data = _RAND_7[63:0];
  _RAND_8 = {2{`RANDOM}};
  r_1_2_data = _RAND_8[63:0];
  _RAND_9 = {2{`RANDOM}};
  r_1_3_data = _RAND_9[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Cache_2(
  input         clock,
  input         reset,
  output        io_in_req_ready, // @[src/main/scala/nutcore/mem/Cache.scala 122:14]
  input         io_in_req_valid, // @[src/main/scala/nutcore/mem/Cache.scala 122:14]
  input  [31:0] io_in_req_bits_addr, // @[src/main/scala/nutcore/mem/Cache.scala 122:14]
  input  [2:0]  io_in_req_bits_size, // @[src/main/scala/nutcore/mem/Cache.scala 122:14]
  input  [3:0]  io_in_req_bits_cmd, // @[src/main/scala/nutcore/mem/Cache.scala 122:14]
  input  [7:0]  io_in_req_bits_wmask, // @[src/main/scala/nutcore/mem/Cache.scala 122:14]
  input  [63:0] io_in_req_bits_wdata, // @[src/main/scala/nutcore/mem/Cache.scala 122:14]
  output        io_in_resp_valid, // @[src/main/scala/nutcore/mem/Cache.scala 122:14]
  output [3:0]  io_in_resp_bits_cmd, // @[src/main/scala/nutcore/mem/Cache.scala 122:14]
  output [63:0] io_in_resp_bits_rdata, // @[src/main/scala/nutcore/mem/Cache.scala 122:14]
  input         io_out_mem_req_ready, // @[src/main/scala/nutcore/mem/Cache.scala 122:14]
  output        io_out_mem_req_valid, // @[src/main/scala/nutcore/mem/Cache.scala 122:14]
  output [31:0] io_out_mem_req_bits_addr, // @[src/main/scala/nutcore/mem/Cache.scala 122:14]
  output [3:0]  io_out_mem_req_bits_cmd, // @[src/main/scala/nutcore/mem/Cache.scala 122:14]
  output [63:0] io_out_mem_req_bits_wdata, // @[src/main/scala/nutcore/mem/Cache.scala 122:14]
  input         io_out_mem_resp_valid, // @[src/main/scala/nutcore/mem/Cache.scala 122:14]
  input  [3:0]  io_out_mem_resp_bits_cmd, // @[src/main/scala/nutcore/mem/Cache.scala 122:14]
  input  [63:0] io_out_mem_resp_bits_rdata, // @[src/main/scala/nutcore/mem/Cache.scala 122:14]
  input         DISPLAY_ENABLE
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [63:0] _RAND_24;
  reg [63:0] _RAND_25;
  reg [63:0] _RAND_26;
  reg [63:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [63:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [63:0] _RAND_34;
  reg [63:0] _RAND_35;
  reg [63:0] _RAND_36;
  reg [63:0] _RAND_37;
  reg [63:0] _RAND_38;
`endif // RANDOMIZE_REG_INIT
  wire  s1_clock; // @[src/main/scala/nutcore/mem/Cache.scala 480:18]
  wire  s1_reset; // @[src/main/scala/nutcore/mem/Cache.scala 480:18]
  wire  s1_io_in_ready; // @[src/main/scala/nutcore/mem/Cache.scala 480:18]
  wire  s1_io_in_valid; // @[src/main/scala/nutcore/mem/Cache.scala 480:18]
  wire [31:0] s1_io_in_bits_addr; // @[src/main/scala/nutcore/mem/Cache.scala 480:18]
  wire [2:0] s1_io_in_bits_size; // @[src/main/scala/nutcore/mem/Cache.scala 480:18]
  wire [3:0] s1_io_in_bits_cmd; // @[src/main/scala/nutcore/mem/Cache.scala 480:18]
  wire [7:0] s1_io_in_bits_wmask; // @[src/main/scala/nutcore/mem/Cache.scala 480:18]
  wire [63:0] s1_io_in_bits_wdata; // @[src/main/scala/nutcore/mem/Cache.scala 480:18]
  wire  s1_io_out_ready; // @[src/main/scala/nutcore/mem/Cache.scala 480:18]
  wire  s1_io_out_valid; // @[src/main/scala/nutcore/mem/Cache.scala 480:18]
  wire [31:0] s1_io_out_bits_req_addr; // @[src/main/scala/nutcore/mem/Cache.scala 480:18]
  wire [2:0] s1_io_out_bits_req_size; // @[src/main/scala/nutcore/mem/Cache.scala 480:18]
  wire [3:0] s1_io_out_bits_req_cmd; // @[src/main/scala/nutcore/mem/Cache.scala 480:18]
  wire [7:0] s1_io_out_bits_req_wmask; // @[src/main/scala/nutcore/mem/Cache.scala 480:18]
  wire [63:0] s1_io_out_bits_req_wdata; // @[src/main/scala/nutcore/mem/Cache.scala 480:18]
  wire  s1_io_metaReadBus_req_ready; // @[src/main/scala/nutcore/mem/Cache.scala 480:18]
  wire  s1_io_metaReadBus_req_valid; // @[src/main/scala/nutcore/mem/Cache.scala 480:18]
  wire [8:0] s1_io_metaReadBus_req_bits_setIdx; // @[src/main/scala/nutcore/mem/Cache.scala 480:18]
  wire [16:0] s1_io_metaReadBus_resp_data_0_tag; // @[src/main/scala/nutcore/mem/Cache.scala 480:18]
  wire  s1_io_metaReadBus_resp_data_0_valid; // @[src/main/scala/nutcore/mem/Cache.scala 480:18]
  wire  s1_io_metaReadBus_resp_data_0_dirty; // @[src/main/scala/nutcore/mem/Cache.scala 480:18]
  wire [16:0] s1_io_metaReadBus_resp_data_1_tag; // @[src/main/scala/nutcore/mem/Cache.scala 480:18]
  wire  s1_io_metaReadBus_resp_data_1_valid; // @[src/main/scala/nutcore/mem/Cache.scala 480:18]
  wire  s1_io_metaReadBus_resp_data_1_dirty; // @[src/main/scala/nutcore/mem/Cache.scala 480:18]
  wire [16:0] s1_io_metaReadBus_resp_data_2_tag; // @[src/main/scala/nutcore/mem/Cache.scala 480:18]
  wire  s1_io_metaReadBus_resp_data_2_valid; // @[src/main/scala/nutcore/mem/Cache.scala 480:18]
  wire  s1_io_metaReadBus_resp_data_2_dirty; // @[src/main/scala/nutcore/mem/Cache.scala 480:18]
  wire [16:0] s1_io_metaReadBus_resp_data_3_tag; // @[src/main/scala/nutcore/mem/Cache.scala 480:18]
  wire  s1_io_metaReadBus_resp_data_3_valid; // @[src/main/scala/nutcore/mem/Cache.scala 480:18]
  wire  s1_io_metaReadBus_resp_data_3_dirty; // @[src/main/scala/nutcore/mem/Cache.scala 480:18]
  wire  s1_io_dataReadBus_req_ready; // @[src/main/scala/nutcore/mem/Cache.scala 480:18]
  wire  s1_io_dataReadBus_req_valid; // @[src/main/scala/nutcore/mem/Cache.scala 480:18]
  wire [11:0] s1_io_dataReadBus_req_bits_setIdx; // @[src/main/scala/nutcore/mem/Cache.scala 480:18]
  wire [63:0] s1_io_dataReadBus_resp_data_0_data; // @[src/main/scala/nutcore/mem/Cache.scala 480:18]
  wire [63:0] s1_io_dataReadBus_resp_data_1_data; // @[src/main/scala/nutcore/mem/Cache.scala 480:18]
  wire [63:0] s1_io_dataReadBus_resp_data_2_data; // @[src/main/scala/nutcore/mem/Cache.scala 480:18]
  wire [63:0] s1_io_dataReadBus_resp_data_3_data; // @[src/main/scala/nutcore/mem/Cache.scala 480:18]
  wire  s1_DISPLAY_ENABLE; // @[src/main/scala/nutcore/mem/Cache.scala 480:18]
  wire  s2_clock; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire  s2_reset; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire  s2_io_in_ready; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire  s2_io_in_valid; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire [31:0] s2_io_in_bits_req_addr; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire [2:0] s2_io_in_bits_req_size; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire [3:0] s2_io_in_bits_req_cmd; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire [7:0] s2_io_in_bits_req_wmask; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire [63:0] s2_io_in_bits_req_wdata; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire  s2_io_out_ready; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire  s2_io_out_valid; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire [31:0] s2_io_out_bits_req_addr; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire [2:0] s2_io_out_bits_req_size; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire [3:0] s2_io_out_bits_req_cmd; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire [7:0] s2_io_out_bits_req_wmask; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire [63:0] s2_io_out_bits_req_wdata; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire [16:0] s2_io_out_bits_metas_0_tag; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire  s2_io_out_bits_metas_0_valid; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire  s2_io_out_bits_metas_0_dirty; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire [16:0] s2_io_out_bits_metas_1_tag; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire  s2_io_out_bits_metas_1_valid; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire  s2_io_out_bits_metas_1_dirty; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire [16:0] s2_io_out_bits_metas_2_tag; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire  s2_io_out_bits_metas_2_valid; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire  s2_io_out_bits_metas_2_dirty; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire [16:0] s2_io_out_bits_metas_3_tag; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire  s2_io_out_bits_metas_3_valid; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire  s2_io_out_bits_metas_3_dirty; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire [63:0] s2_io_out_bits_datas_0_data; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire [63:0] s2_io_out_bits_datas_1_data; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire [63:0] s2_io_out_bits_datas_2_data; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire [63:0] s2_io_out_bits_datas_3_data; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire  s2_io_out_bits_hit; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire [3:0] s2_io_out_bits_waymask; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire  s2_io_out_bits_mmio; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire  s2_io_out_bits_isForwardData; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire [63:0] s2_io_out_bits_forwardData_data_data; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire [3:0] s2_io_out_bits_forwardData_waymask; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire [16:0] s2_io_metaReadResp_0_tag; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire  s2_io_metaReadResp_0_valid; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire  s2_io_metaReadResp_0_dirty; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire [16:0] s2_io_metaReadResp_1_tag; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire  s2_io_metaReadResp_1_valid; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire  s2_io_metaReadResp_1_dirty; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire [16:0] s2_io_metaReadResp_2_tag; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire  s2_io_metaReadResp_2_valid; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire  s2_io_metaReadResp_2_dirty; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire [16:0] s2_io_metaReadResp_3_tag; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire  s2_io_metaReadResp_3_valid; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire  s2_io_metaReadResp_3_dirty; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire [63:0] s2_io_dataReadResp_0_data; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire [63:0] s2_io_dataReadResp_1_data; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire [63:0] s2_io_dataReadResp_2_data; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire [63:0] s2_io_dataReadResp_3_data; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire  s2_io_metaWriteBus_req_valid; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire [8:0] s2_io_metaWriteBus_req_bits_setIdx; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire [16:0] s2_io_metaWriteBus_req_bits_data_tag; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire  s2_io_metaWriteBus_req_bits_data_dirty; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire [3:0] s2_io_metaWriteBus_req_bits_waymask; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire  s2_io_dataWriteBus_req_valid; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire [11:0] s2_io_dataWriteBus_req_bits_setIdx; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire [63:0] s2_io_dataWriteBus_req_bits_data_data; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire [3:0] s2_io_dataWriteBus_req_bits_waymask; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire  s2_DISPLAY_ENABLE; // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
  wire  s3_clock; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire  s3_reset; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire  s3_io_in_ready; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire  s3_io_in_valid; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire [31:0] s3_io_in_bits_req_addr; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire [2:0] s3_io_in_bits_req_size; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire [3:0] s3_io_in_bits_req_cmd; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire [7:0] s3_io_in_bits_req_wmask; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire [63:0] s3_io_in_bits_req_wdata; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire [16:0] s3_io_in_bits_metas_0_tag; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire  s3_io_in_bits_metas_0_valid; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire  s3_io_in_bits_metas_0_dirty; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire [16:0] s3_io_in_bits_metas_1_tag; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire  s3_io_in_bits_metas_1_valid; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire  s3_io_in_bits_metas_1_dirty; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire [16:0] s3_io_in_bits_metas_2_tag; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire  s3_io_in_bits_metas_2_valid; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire  s3_io_in_bits_metas_2_dirty; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire [16:0] s3_io_in_bits_metas_3_tag; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire  s3_io_in_bits_metas_3_valid; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire  s3_io_in_bits_metas_3_dirty; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire [63:0] s3_io_in_bits_datas_0_data; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire [63:0] s3_io_in_bits_datas_1_data; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire [63:0] s3_io_in_bits_datas_2_data; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire [63:0] s3_io_in_bits_datas_3_data; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire  s3_io_in_bits_hit; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire [3:0] s3_io_in_bits_waymask; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire  s3_io_in_bits_mmio; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire  s3_io_in_bits_isForwardData; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire [63:0] s3_io_in_bits_forwardData_data_data; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire [3:0] s3_io_in_bits_forwardData_waymask; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire  s3_io_out_ready; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire  s3_io_out_valid; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire [3:0] s3_io_out_bits_cmd; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire [63:0] s3_io_out_bits_rdata; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire  s3_io_isFinish; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire  s3_io_dataReadBus_req_ready; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire  s3_io_dataReadBus_req_valid; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire [11:0] s3_io_dataReadBus_req_bits_setIdx; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire [63:0] s3_io_dataReadBus_resp_data_0_data; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire [63:0] s3_io_dataReadBus_resp_data_1_data; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire [63:0] s3_io_dataReadBus_resp_data_2_data; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire [63:0] s3_io_dataReadBus_resp_data_3_data; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire  s3_io_dataWriteBus_req_valid; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire [11:0] s3_io_dataWriteBus_req_bits_setIdx; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire [63:0] s3_io_dataWriteBus_req_bits_data_data; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire [3:0] s3_io_dataWriteBus_req_bits_waymask; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire  s3_io_metaWriteBus_req_valid; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire [8:0] s3_io_metaWriteBus_req_bits_setIdx; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire [16:0] s3_io_metaWriteBus_req_bits_data_tag; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire  s3_io_metaWriteBus_req_bits_data_valid; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire  s3_io_metaWriteBus_req_bits_data_dirty; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire [3:0] s3_io_metaWriteBus_req_bits_waymask; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire  s3_io_mem_req_ready; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire  s3_io_mem_req_valid; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire [31:0] s3_io_mem_req_bits_addr; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire [2:0] s3_io_mem_req_bits_size; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire [3:0] s3_io_mem_req_bits_cmd; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire [7:0] s3_io_mem_req_bits_wmask; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire [63:0] s3_io_mem_req_bits_wdata; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire  s3_io_mem_resp_ready; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire  s3_io_mem_resp_valid; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire [3:0] s3_io_mem_resp_bits_cmd; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire [63:0] s3_io_mem_resp_bits_rdata; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire  s3_io_cohResp_valid; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire  s3_io_dataReadRespToL1; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire  s3_DISPLAY_ENABLE; // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
  wire  metaArray_clock; // @[src/main/scala/nutcore/mem/Cache.scala 483:25]
  wire  metaArray_reset; // @[src/main/scala/nutcore/mem/Cache.scala 483:25]
  wire  metaArray_io_r_0_req_ready; // @[src/main/scala/nutcore/mem/Cache.scala 483:25]
  wire  metaArray_io_r_0_req_valid; // @[src/main/scala/nutcore/mem/Cache.scala 483:25]
  wire [8:0] metaArray_io_r_0_req_bits_setIdx; // @[src/main/scala/nutcore/mem/Cache.scala 483:25]
  wire [16:0] metaArray_io_r_0_resp_data_0_tag; // @[src/main/scala/nutcore/mem/Cache.scala 483:25]
  wire  metaArray_io_r_0_resp_data_0_valid; // @[src/main/scala/nutcore/mem/Cache.scala 483:25]
  wire  metaArray_io_r_0_resp_data_0_dirty; // @[src/main/scala/nutcore/mem/Cache.scala 483:25]
  wire [16:0] metaArray_io_r_0_resp_data_1_tag; // @[src/main/scala/nutcore/mem/Cache.scala 483:25]
  wire  metaArray_io_r_0_resp_data_1_valid; // @[src/main/scala/nutcore/mem/Cache.scala 483:25]
  wire  metaArray_io_r_0_resp_data_1_dirty; // @[src/main/scala/nutcore/mem/Cache.scala 483:25]
  wire [16:0] metaArray_io_r_0_resp_data_2_tag; // @[src/main/scala/nutcore/mem/Cache.scala 483:25]
  wire  metaArray_io_r_0_resp_data_2_valid; // @[src/main/scala/nutcore/mem/Cache.scala 483:25]
  wire  metaArray_io_r_0_resp_data_2_dirty; // @[src/main/scala/nutcore/mem/Cache.scala 483:25]
  wire [16:0] metaArray_io_r_0_resp_data_3_tag; // @[src/main/scala/nutcore/mem/Cache.scala 483:25]
  wire  metaArray_io_r_0_resp_data_3_valid; // @[src/main/scala/nutcore/mem/Cache.scala 483:25]
  wire  metaArray_io_r_0_resp_data_3_dirty; // @[src/main/scala/nutcore/mem/Cache.scala 483:25]
  wire  metaArray_io_w_req_valid; // @[src/main/scala/nutcore/mem/Cache.scala 483:25]
  wire [8:0] metaArray_io_w_req_bits_setIdx; // @[src/main/scala/nutcore/mem/Cache.scala 483:25]
  wire [16:0] metaArray_io_w_req_bits_data_tag; // @[src/main/scala/nutcore/mem/Cache.scala 483:25]
  wire  metaArray_io_w_req_bits_data_dirty; // @[src/main/scala/nutcore/mem/Cache.scala 483:25]
  wire [3:0] metaArray_io_w_req_bits_waymask; // @[src/main/scala/nutcore/mem/Cache.scala 483:25]
  wire  dataArray_clock; // @[src/main/scala/nutcore/mem/Cache.scala 484:25]
  wire  dataArray_reset; // @[src/main/scala/nutcore/mem/Cache.scala 484:25]
  wire  dataArray_io_r_0_req_ready; // @[src/main/scala/nutcore/mem/Cache.scala 484:25]
  wire  dataArray_io_r_0_req_valid; // @[src/main/scala/nutcore/mem/Cache.scala 484:25]
  wire [11:0] dataArray_io_r_0_req_bits_setIdx; // @[src/main/scala/nutcore/mem/Cache.scala 484:25]
  wire [63:0] dataArray_io_r_0_resp_data_0_data; // @[src/main/scala/nutcore/mem/Cache.scala 484:25]
  wire [63:0] dataArray_io_r_0_resp_data_1_data; // @[src/main/scala/nutcore/mem/Cache.scala 484:25]
  wire [63:0] dataArray_io_r_0_resp_data_2_data; // @[src/main/scala/nutcore/mem/Cache.scala 484:25]
  wire [63:0] dataArray_io_r_0_resp_data_3_data; // @[src/main/scala/nutcore/mem/Cache.scala 484:25]
  wire  dataArray_io_r_1_req_ready; // @[src/main/scala/nutcore/mem/Cache.scala 484:25]
  wire  dataArray_io_r_1_req_valid; // @[src/main/scala/nutcore/mem/Cache.scala 484:25]
  wire [11:0] dataArray_io_r_1_req_bits_setIdx; // @[src/main/scala/nutcore/mem/Cache.scala 484:25]
  wire [63:0] dataArray_io_r_1_resp_data_0_data; // @[src/main/scala/nutcore/mem/Cache.scala 484:25]
  wire [63:0] dataArray_io_r_1_resp_data_1_data; // @[src/main/scala/nutcore/mem/Cache.scala 484:25]
  wire [63:0] dataArray_io_r_1_resp_data_2_data; // @[src/main/scala/nutcore/mem/Cache.scala 484:25]
  wire [63:0] dataArray_io_r_1_resp_data_3_data; // @[src/main/scala/nutcore/mem/Cache.scala 484:25]
  wire  dataArray_io_w_req_valid; // @[src/main/scala/nutcore/mem/Cache.scala 484:25]
  wire [11:0] dataArray_io_w_req_bits_setIdx; // @[src/main/scala/nutcore/mem/Cache.scala 484:25]
  wire [63:0] dataArray_io_w_req_bits_data_data; // @[src/main/scala/nutcore/mem/Cache.scala 484:25]
  wire [3:0] dataArray_io_w_req_bits_waymask; // @[src/main/scala/nutcore/mem/Cache.scala 484:25]
  wire  arb_io_in_0_ready; // @[src/main/scala/nutcore/mem/Cache.scala 493:19]
  wire  arb_io_in_0_valid; // @[src/main/scala/nutcore/mem/Cache.scala 493:19]
  wire [31:0] arb_io_in_0_bits_addr; // @[src/main/scala/nutcore/mem/Cache.scala 493:19]
  wire [2:0] arb_io_in_0_bits_size; // @[src/main/scala/nutcore/mem/Cache.scala 493:19]
  wire [3:0] arb_io_in_0_bits_cmd; // @[src/main/scala/nutcore/mem/Cache.scala 493:19]
  wire [7:0] arb_io_in_0_bits_wmask; // @[src/main/scala/nutcore/mem/Cache.scala 493:19]
  wire [63:0] arb_io_in_0_bits_wdata; // @[src/main/scala/nutcore/mem/Cache.scala 493:19]
  wire  arb_io_in_1_ready; // @[src/main/scala/nutcore/mem/Cache.scala 493:19]
  wire  arb_io_in_1_valid; // @[src/main/scala/nutcore/mem/Cache.scala 493:19]
  wire [31:0] arb_io_in_1_bits_addr; // @[src/main/scala/nutcore/mem/Cache.scala 493:19]
  wire [2:0] arb_io_in_1_bits_size; // @[src/main/scala/nutcore/mem/Cache.scala 493:19]
  wire [3:0] arb_io_in_1_bits_cmd; // @[src/main/scala/nutcore/mem/Cache.scala 493:19]
  wire [7:0] arb_io_in_1_bits_wmask; // @[src/main/scala/nutcore/mem/Cache.scala 493:19]
  wire [63:0] arb_io_in_1_bits_wdata; // @[src/main/scala/nutcore/mem/Cache.scala 493:19]
  wire  arb_io_out_ready; // @[src/main/scala/nutcore/mem/Cache.scala 493:19]
  wire  arb_io_out_valid; // @[src/main/scala/nutcore/mem/Cache.scala 493:19]
  wire [31:0] arb_io_out_bits_addr; // @[src/main/scala/nutcore/mem/Cache.scala 493:19]
  wire [2:0] arb_io_out_bits_size; // @[src/main/scala/nutcore/mem/Cache.scala 493:19]
  wire [3:0] arb_io_out_bits_cmd; // @[src/main/scala/nutcore/mem/Cache.scala 493:19]
  wire [7:0] arb_io_out_bits_wmask; // @[src/main/scala/nutcore/mem/Cache.scala 493:19]
  wire [63:0] arb_io_out_bits_wdata; // @[src/main/scala/nutcore/mem/Cache.scala 493:19]
  wire  _T = s2_io_out_ready & s2_io_out_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  reg  valid; // @[src/main/scala/utils/Pipeline.scala 24:24]
  wire  _GEN_0 = _T ? 1'h0 : valid; // @[src/main/scala/utils/Pipeline.scala 24:24 25:{25,33}]
  wire  _T_2 = s1_io_out_valid & s2_io_in_ready; // @[src/main/scala/utils/Pipeline.scala 26:22]
  wire  _GEN_1 = s1_io_out_valid & s2_io_in_ready | _GEN_0; // @[src/main/scala/utils/Pipeline.scala 26:{38,46}]
  reg [31:0] s2_io_in_bits_r_req_addr; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg [2:0] s2_io_in_bits_r_req_size; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg [3:0] s2_io_in_bits_r_req_cmd; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg [7:0] s2_io_in_bits_r_req_wmask; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg [63:0] s2_io_in_bits_r_req_wdata; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg  valid_1; // @[src/main/scala/utils/Pipeline.scala 24:24]
  wire  _GEN_8 = s3_io_isFinish ? 1'h0 : valid_1; // @[src/main/scala/utils/Pipeline.scala 24:24 25:{25,33}]
  wire  _T_4 = s2_io_out_valid & s3_io_in_ready; // @[src/main/scala/utils/Pipeline.scala 26:22]
  wire  _GEN_9 = s2_io_out_valid & s3_io_in_ready | _GEN_8; // @[src/main/scala/utils/Pipeline.scala 26:{38,46}]
  reg [31:0] s3_io_in_bits_r_req_addr; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg [2:0] s3_io_in_bits_r_req_size; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg [3:0] s3_io_in_bits_r_req_cmd; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg [7:0] s3_io_in_bits_r_req_wmask; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg [63:0] s3_io_in_bits_r_req_wdata; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg [16:0] s3_io_in_bits_r_metas_0_tag; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg  s3_io_in_bits_r_metas_0_valid; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg  s3_io_in_bits_r_metas_0_dirty; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg [16:0] s3_io_in_bits_r_metas_1_tag; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg  s3_io_in_bits_r_metas_1_valid; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg  s3_io_in_bits_r_metas_1_dirty; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg [16:0] s3_io_in_bits_r_metas_2_tag; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg  s3_io_in_bits_r_metas_2_valid; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg  s3_io_in_bits_r_metas_2_dirty; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg [16:0] s3_io_in_bits_r_metas_3_tag; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg  s3_io_in_bits_r_metas_3_valid; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg  s3_io_in_bits_r_metas_3_dirty; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg [63:0] s3_io_in_bits_r_datas_0_data; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg [63:0] s3_io_in_bits_r_datas_1_data; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg [63:0] s3_io_in_bits_r_datas_2_data; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg [63:0] s3_io_in_bits_r_datas_3_data; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg  s3_io_in_bits_r_hit; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg [3:0] s3_io_in_bits_r_waymask; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg  s3_io_in_bits_r_mmio; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg  s3_io_in_bits_r_isForwardData; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg [63:0] s3_io_in_bits_r_forwardData_data_data; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg [3:0] s3_io_in_bits_r_forwardData_waymask; // @[src/main/scala/utils/Pipeline.scala 30:28]
  wire  _io_in_resp_valid_T = s3_io_out_bits_cmd == 4'h4; // @[src/main/scala/bus/simplebus/SimpleBus.scala 95:24]
  reg [63:0] c; // @[src/main/scala/utils/GTimer.scala 24:20]
  wire [63:0] _c_T_1 = c + 64'h1; // @[src/main/scala/utils/GTimer.scala 25:12]
  wire  _T_7 = ~reset; // @[src/main/scala/utils/Debug.scala 56:24]
  reg [63:0] c_1; // @[src/main/scala/utils/GTimer.scala 24:20]
  wire [63:0] _c_T_3 = c_1 + 64'h1; // @[src/main/scala/utils/GTimer.scala 25:12]
  reg [63:0] c_2; // @[src/main/scala/utils/GTimer.scala 24:20]
  wire [63:0] _c_T_5 = c_2 + 64'h1; // @[src/main/scala/utils/GTimer.scala 25:12]
  reg [63:0] c_3; // @[src/main/scala/utils/GTimer.scala 24:20]
  wire [63:0] _c_T_7 = c_3 + 64'h1; // @[src/main/scala/utils/GTimer.scala 25:12]
  reg [63:0] c_4; // @[src/main/scala/utils/GTimer.scala 24:20]
  wire [63:0] _c_T_9 = c_4 + 64'h1; // @[src/main/scala/utils/GTimer.scala 25:12]
  wire  _GEN_39 = s1_io_in_valid & DISPLAY_ENABLE; // @[src/main/scala/utils/Debug.scala 56:24]
  wire  _GEN_41 = s2_io_in_valid & DISPLAY_ENABLE; // @[src/main/scala/utils/Debug.scala 56:24]
  wire  _GEN_43 = s3_io_in_valid & DISPLAY_ENABLE; // @[src/main/scala/utils/Debug.scala 56:24]
  CacheStage1_2 s1 ( // @[src/main/scala/nutcore/mem/Cache.scala 480:18]
    .clock(s1_clock),
    .reset(s1_reset),
    .io_in_ready(s1_io_in_ready),
    .io_in_valid(s1_io_in_valid),
    .io_in_bits_addr(s1_io_in_bits_addr),
    .io_in_bits_size(s1_io_in_bits_size),
    .io_in_bits_cmd(s1_io_in_bits_cmd),
    .io_in_bits_wmask(s1_io_in_bits_wmask),
    .io_in_bits_wdata(s1_io_in_bits_wdata),
    .io_out_ready(s1_io_out_ready),
    .io_out_valid(s1_io_out_valid),
    .io_out_bits_req_addr(s1_io_out_bits_req_addr),
    .io_out_bits_req_size(s1_io_out_bits_req_size),
    .io_out_bits_req_cmd(s1_io_out_bits_req_cmd),
    .io_out_bits_req_wmask(s1_io_out_bits_req_wmask),
    .io_out_bits_req_wdata(s1_io_out_bits_req_wdata),
    .io_metaReadBus_req_ready(s1_io_metaReadBus_req_ready),
    .io_metaReadBus_req_valid(s1_io_metaReadBus_req_valid),
    .io_metaReadBus_req_bits_setIdx(s1_io_metaReadBus_req_bits_setIdx),
    .io_metaReadBus_resp_data_0_tag(s1_io_metaReadBus_resp_data_0_tag),
    .io_metaReadBus_resp_data_0_valid(s1_io_metaReadBus_resp_data_0_valid),
    .io_metaReadBus_resp_data_0_dirty(s1_io_metaReadBus_resp_data_0_dirty),
    .io_metaReadBus_resp_data_1_tag(s1_io_metaReadBus_resp_data_1_tag),
    .io_metaReadBus_resp_data_1_valid(s1_io_metaReadBus_resp_data_1_valid),
    .io_metaReadBus_resp_data_1_dirty(s1_io_metaReadBus_resp_data_1_dirty),
    .io_metaReadBus_resp_data_2_tag(s1_io_metaReadBus_resp_data_2_tag),
    .io_metaReadBus_resp_data_2_valid(s1_io_metaReadBus_resp_data_2_valid),
    .io_metaReadBus_resp_data_2_dirty(s1_io_metaReadBus_resp_data_2_dirty),
    .io_metaReadBus_resp_data_3_tag(s1_io_metaReadBus_resp_data_3_tag),
    .io_metaReadBus_resp_data_3_valid(s1_io_metaReadBus_resp_data_3_valid),
    .io_metaReadBus_resp_data_3_dirty(s1_io_metaReadBus_resp_data_3_dirty),
    .io_dataReadBus_req_ready(s1_io_dataReadBus_req_ready),
    .io_dataReadBus_req_valid(s1_io_dataReadBus_req_valid),
    .io_dataReadBus_req_bits_setIdx(s1_io_dataReadBus_req_bits_setIdx),
    .io_dataReadBus_resp_data_0_data(s1_io_dataReadBus_resp_data_0_data),
    .io_dataReadBus_resp_data_1_data(s1_io_dataReadBus_resp_data_1_data),
    .io_dataReadBus_resp_data_2_data(s1_io_dataReadBus_resp_data_2_data),
    .io_dataReadBus_resp_data_3_data(s1_io_dataReadBus_resp_data_3_data),
    .DISPLAY_ENABLE(s1_DISPLAY_ENABLE)
  );
  CacheStage2_2 s2 ( // @[src/main/scala/nutcore/mem/Cache.scala 481:18]
    .clock(s2_clock),
    .reset(s2_reset),
    .io_in_ready(s2_io_in_ready),
    .io_in_valid(s2_io_in_valid),
    .io_in_bits_req_addr(s2_io_in_bits_req_addr),
    .io_in_bits_req_size(s2_io_in_bits_req_size),
    .io_in_bits_req_cmd(s2_io_in_bits_req_cmd),
    .io_in_bits_req_wmask(s2_io_in_bits_req_wmask),
    .io_in_bits_req_wdata(s2_io_in_bits_req_wdata),
    .io_out_ready(s2_io_out_ready),
    .io_out_valid(s2_io_out_valid),
    .io_out_bits_req_addr(s2_io_out_bits_req_addr),
    .io_out_bits_req_size(s2_io_out_bits_req_size),
    .io_out_bits_req_cmd(s2_io_out_bits_req_cmd),
    .io_out_bits_req_wmask(s2_io_out_bits_req_wmask),
    .io_out_bits_req_wdata(s2_io_out_bits_req_wdata),
    .io_out_bits_metas_0_tag(s2_io_out_bits_metas_0_tag),
    .io_out_bits_metas_0_valid(s2_io_out_bits_metas_0_valid),
    .io_out_bits_metas_0_dirty(s2_io_out_bits_metas_0_dirty),
    .io_out_bits_metas_1_tag(s2_io_out_bits_metas_1_tag),
    .io_out_bits_metas_1_valid(s2_io_out_bits_metas_1_valid),
    .io_out_bits_metas_1_dirty(s2_io_out_bits_metas_1_dirty),
    .io_out_bits_metas_2_tag(s2_io_out_bits_metas_2_tag),
    .io_out_bits_metas_2_valid(s2_io_out_bits_metas_2_valid),
    .io_out_bits_metas_2_dirty(s2_io_out_bits_metas_2_dirty),
    .io_out_bits_metas_3_tag(s2_io_out_bits_metas_3_tag),
    .io_out_bits_metas_3_valid(s2_io_out_bits_metas_3_valid),
    .io_out_bits_metas_3_dirty(s2_io_out_bits_metas_3_dirty),
    .io_out_bits_datas_0_data(s2_io_out_bits_datas_0_data),
    .io_out_bits_datas_1_data(s2_io_out_bits_datas_1_data),
    .io_out_bits_datas_2_data(s2_io_out_bits_datas_2_data),
    .io_out_bits_datas_3_data(s2_io_out_bits_datas_3_data),
    .io_out_bits_hit(s2_io_out_bits_hit),
    .io_out_bits_waymask(s2_io_out_bits_waymask),
    .io_out_bits_mmio(s2_io_out_bits_mmio),
    .io_out_bits_isForwardData(s2_io_out_bits_isForwardData),
    .io_out_bits_forwardData_data_data(s2_io_out_bits_forwardData_data_data),
    .io_out_bits_forwardData_waymask(s2_io_out_bits_forwardData_waymask),
    .io_metaReadResp_0_tag(s2_io_metaReadResp_0_tag),
    .io_metaReadResp_0_valid(s2_io_metaReadResp_0_valid),
    .io_metaReadResp_0_dirty(s2_io_metaReadResp_0_dirty),
    .io_metaReadResp_1_tag(s2_io_metaReadResp_1_tag),
    .io_metaReadResp_1_valid(s2_io_metaReadResp_1_valid),
    .io_metaReadResp_1_dirty(s2_io_metaReadResp_1_dirty),
    .io_metaReadResp_2_tag(s2_io_metaReadResp_2_tag),
    .io_metaReadResp_2_valid(s2_io_metaReadResp_2_valid),
    .io_metaReadResp_2_dirty(s2_io_metaReadResp_2_dirty),
    .io_metaReadResp_3_tag(s2_io_metaReadResp_3_tag),
    .io_metaReadResp_3_valid(s2_io_metaReadResp_3_valid),
    .io_metaReadResp_3_dirty(s2_io_metaReadResp_3_dirty),
    .io_dataReadResp_0_data(s2_io_dataReadResp_0_data),
    .io_dataReadResp_1_data(s2_io_dataReadResp_1_data),
    .io_dataReadResp_2_data(s2_io_dataReadResp_2_data),
    .io_dataReadResp_3_data(s2_io_dataReadResp_3_data),
    .io_metaWriteBus_req_valid(s2_io_metaWriteBus_req_valid),
    .io_metaWriteBus_req_bits_setIdx(s2_io_metaWriteBus_req_bits_setIdx),
    .io_metaWriteBus_req_bits_data_tag(s2_io_metaWriteBus_req_bits_data_tag),
    .io_metaWriteBus_req_bits_data_dirty(s2_io_metaWriteBus_req_bits_data_dirty),
    .io_metaWriteBus_req_bits_waymask(s2_io_metaWriteBus_req_bits_waymask),
    .io_dataWriteBus_req_valid(s2_io_dataWriteBus_req_valid),
    .io_dataWriteBus_req_bits_setIdx(s2_io_dataWriteBus_req_bits_setIdx),
    .io_dataWriteBus_req_bits_data_data(s2_io_dataWriteBus_req_bits_data_data),
    .io_dataWriteBus_req_bits_waymask(s2_io_dataWriteBus_req_bits_waymask),
    .DISPLAY_ENABLE(s2_DISPLAY_ENABLE)
  );
  CacheStage3_2 s3 ( // @[src/main/scala/nutcore/mem/Cache.scala 482:18]
    .clock(s3_clock),
    .reset(s3_reset),
    .io_in_ready(s3_io_in_ready),
    .io_in_valid(s3_io_in_valid),
    .io_in_bits_req_addr(s3_io_in_bits_req_addr),
    .io_in_bits_req_size(s3_io_in_bits_req_size),
    .io_in_bits_req_cmd(s3_io_in_bits_req_cmd),
    .io_in_bits_req_wmask(s3_io_in_bits_req_wmask),
    .io_in_bits_req_wdata(s3_io_in_bits_req_wdata),
    .io_in_bits_metas_0_tag(s3_io_in_bits_metas_0_tag),
    .io_in_bits_metas_0_valid(s3_io_in_bits_metas_0_valid),
    .io_in_bits_metas_0_dirty(s3_io_in_bits_metas_0_dirty),
    .io_in_bits_metas_1_tag(s3_io_in_bits_metas_1_tag),
    .io_in_bits_metas_1_valid(s3_io_in_bits_metas_1_valid),
    .io_in_bits_metas_1_dirty(s3_io_in_bits_metas_1_dirty),
    .io_in_bits_metas_2_tag(s3_io_in_bits_metas_2_tag),
    .io_in_bits_metas_2_valid(s3_io_in_bits_metas_2_valid),
    .io_in_bits_metas_2_dirty(s3_io_in_bits_metas_2_dirty),
    .io_in_bits_metas_3_tag(s3_io_in_bits_metas_3_tag),
    .io_in_bits_metas_3_valid(s3_io_in_bits_metas_3_valid),
    .io_in_bits_metas_3_dirty(s3_io_in_bits_metas_3_dirty),
    .io_in_bits_datas_0_data(s3_io_in_bits_datas_0_data),
    .io_in_bits_datas_1_data(s3_io_in_bits_datas_1_data),
    .io_in_bits_datas_2_data(s3_io_in_bits_datas_2_data),
    .io_in_bits_datas_3_data(s3_io_in_bits_datas_3_data),
    .io_in_bits_hit(s3_io_in_bits_hit),
    .io_in_bits_waymask(s3_io_in_bits_waymask),
    .io_in_bits_mmio(s3_io_in_bits_mmio),
    .io_in_bits_isForwardData(s3_io_in_bits_isForwardData),
    .io_in_bits_forwardData_data_data(s3_io_in_bits_forwardData_data_data),
    .io_in_bits_forwardData_waymask(s3_io_in_bits_forwardData_waymask),
    .io_out_ready(s3_io_out_ready),
    .io_out_valid(s3_io_out_valid),
    .io_out_bits_cmd(s3_io_out_bits_cmd),
    .io_out_bits_rdata(s3_io_out_bits_rdata),
    .io_isFinish(s3_io_isFinish),
    .io_dataReadBus_req_ready(s3_io_dataReadBus_req_ready),
    .io_dataReadBus_req_valid(s3_io_dataReadBus_req_valid),
    .io_dataReadBus_req_bits_setIdx(s3_io_dataReadBus_req_bits_setIdx),
    .io_dataReadBus_resp_data_0_data(s3_io_dataReadBus_resp_data_0_data),
    .io_dataReadBus_resp_data_1_data(s3_io_dataReadBus_resp_data_1_data),
    .io_dataReadBus_resp_data_2_data(s3_io_dataReadBus_resp_data_2_data),
    .io_dataReadBus_resp_data_3_data(s3_io_dataReadBus_resp_data_3_data),
    .io_dataWriteBus_req_valid(s3_io_dataWriteBus_req_valid),
    .io_dataWriteBus_req_bits_setIdx(s3_io_dataWriteBus_req_bits_setIdx),
    .io_dataWriteBus_req_bits_data_data(s3_io_dataWriteBus_req_bits_data_data),
    .io_dataWriteBus_req_bits_waymask(s3_io_dataWriteBus_req_bits_waymask),
    .io_metaWriteBus_req_valid(s3_io_metaWriteBus_req_valid),
    .io_metaWriteBus_req_bits_setIdx(s3_io_metaWriteBus_req_bits_setIdx),
    .io_metaWriteBus_req_bits_data_tag(s3_io_metaWriteBus_req_bits_data_tag),
    .io_metaWriteBus_req_bits_data_valid(s3_io_metaWriteBus_req_bits_data_valid),
    .io_metaWriteBus_req_bits_data_dirty(s3_io_metaWriteBus_req_bits_data_dirty),
    .io_metaWriteBus_req_bits_waymask(s3_io_metaWriteBus_req_bits_waymask),
    .io_mem_req_ready(s3_io_mem_req_ready),
    .io_mem_req_valid(s3_io_mem_req_valid),
    .io_mem_req_bits_addr(s3_io_mem_req_bits_addr),
    .io_mem_req_bits_size(s3_io_mem_req_bits_size),
    .io_mem_req_bits_cmd(s3_io_mem_req_bits_cmd),
    .io_mem_req_bits_wmask(s3_io_mem_req_bits_wmask),
    .io_mem_req_bits_wdata(s3_io_mem_req_bits_wdata),
    .io_mem_resp_ready(s3_io_mem_resp_ready),
    .io_mem_resp_valid(s3_io_mem_resp_valid),
    .io_mem_resp_bits_cmd(s3_io_mem_resp_bits_cmd),
    .io_mem_resp_bits_rdata(s3_io_mem_resp_bits_rdata),
    .io_cohResp_valid(s3_io_cohResp_valid),
    .io_dataReadRespToL1(s3_io_dataReadRespToL1),
    .DISPLAY_ENABLE(s3_DISPLAY_ENABLE)
  );
  SRAMTemplateWithArbiter_4 metaArray ( // @[src/main/scala/nutcore/mem/Cache.scala 483:25]
    .clock(metaArray_clock),
    .reset(metaArray_reset),
    .io_r_0_req_ready(metaArray_io_r_0_req_ready),
    .io_r_0_req_valid(metaArray_io_r_0_req_valid),
    .io_r_0_req_bits_setIdx(metaArray_io_r_0_req_bits_setIdx),
    .io_r_0_resp_data_0_tag(metaArray_io_r_0_resp_data_0_tag),
    .io_r_0_resp_data_0_valid(metaArray_io_r_0_resp_data_0_valid),
    .io_r_0_resp_data_0_dirty(metaArray_io_r_0_resp_data_0_dirty),
    .io_r_0_resp_data_1_tag(metaArray_io_r_0_resp_data_1_tag),
    .io_r_0_resp_data_1_valid(metaArray_io_r_0_resp_data_1_valid),
    .io_r_0_resp_data_1_dirty(metaArray_io_r_0_resp_data_1_dirty),
    .io_r_0_resp_data_2_tag(metaArray_io_r_0_resp_data_2_tag),
    .io_r_0_resp_data_2_valid(metaArray_io_r_0_resp_data_2_valid),
    .io_r_0_resp_data_2_dirty(metaArray_io_r_0_resp_data_2_dirty),
    .io_r_0_resp_data_3_tag(metaArray_io_r_0_resp_data_3_tag),
    .io_r_0_resp_data_3_valid(metaArray_io_r_0_resp_data_3_valid),
    .io_r_0_resp_data_3_dirty(metaArray_io_r_0_resp_data_3_dirty),
    .io_w_req_valid(metaArray_io_w_req_valid),
    .io_w_req_bits_setIdx(metaArray_io_w_req_bits_setIdx),
    .io_w_req_bits_data_tag(metaArray_io_w_req_bits_data_tag),
    .io_w_req_bits_data_dirty(metaArray_io_w_req_bits_data_dirty),
    .io_w_req_bits_waymask(metaArray_io_w_req_bits_waymask)
  );
  SRAMTemplateWithArbiter_5 dataArray ( // @[src/main/scala/nutcore/mem/Cache.scala 484:25]
    .clock(dataArray_clock),
    .reset(dataArray_reset),
    .io_r_0_req_ready(dataArray_io_r_0_req_ready),
    .io_r_0_req_valid(dataArray_io_r_0_req_valid),
    .io_r_0_req_bits_setIdx(dataArray_io_r_0_req_bits_setIdx),
    .io_r_0_resp_data_0_data(dataArray_io_r_0_resp_data_0_data),
    .io_r_0_resp_data_1_data(dataArray_io_r_0_resp_data_1_data),
    .io_r_0_resp_data_2_data(dataArray_io_r_0_resp_data_2_data),
    .io_r_0_resp_data_3_data(dataArray_io_r_0_resp_data_3_data),
    .io_r_1_req_ready(dataArray_io_r_1_req_ready),
    .io_r_1_req_valid(dataArray_io_r_1_req_valid),
    .io_r_1_req_bits_setIdx(dataArray_io_r_1_req_bits_setIdx),
    .io_r_1_resp_data_0_data(dataArray_io_r_1_resp_data_0_data),
    .io_r_1_resp_data_1_data(dataArray_io_r_1_resp_data_1_data),
    .io_r_1_resp_data_2_data(dataArray_io_r_1_resp_data_2_data),
    .io_r_1_resp_data_3_data(dataArray_io_r_1_resp_data_3_data),
    .io_w_req_valid(dataArray_io_w_req_valid),
    .io_w_req_bits_setIdx(dataArray_io_w_req_bits_setIdx),
    .io_w_req_bits_data_data(dataArray_io_w_req_bits_data_data),
    .io_w_req_bits_waymask(dataArray_io_w_req_bits_waymask)
  );
  Arbiter_9 arb ( // @[src/main/scala/nutcore/mem/Cache.scala 493:19]
    .io_in_0_ready(arb_io_in_0_ready),
    .io_in_0_valid(arb_io_in_0_valid),
    .io_in_0_bits_addr(arb_io_in_0_bits_addr),
    .io_in_0_bits_size(arb_io_in_0_bits_size),
    .io_in_0_bits_cmd(arb_io_in_0_bits_cmd),
    .io_in_0_bits_wmask(arb_io_in_0_bits_wmask),
    .io_in_0_bits_wdata(arb_io_in_0_bits_wdata),
    .io_in_1_ready(arb_io_in_1_ready),
    .io_in_1_valid(arb_io_in_1_valid),
    .io_in_1_bits_addr(arb_io_in_1_bits_addr),
    .io_in_1_bits_size(arb_io_in_1_bits_size),
    .io_in_1_bits_cmd(arb_io_in_1_bits_cmd),
    .io_in_1_bits_wmask(arb_io_in_1_bits_wmask),
    .io_in_1_bits_wdata(arb_io_in_1_bits_wdata),
    .io_out_ready(arb_io_out_ready),
    .io_out_valid(arb_io_out_valid),
    .io_out_bits_addr(arb_io_out_bits_addr),
    .io_out_bits_size(arb_io_out_bits_size),
    .io_out_bits_cmd(arb_io_out_bits_cmd),
    .io_out_bits_wmask(arb_io_out_bits_wmask),
    .io_out_bits_wdata(arb_io_out_bits_wdata)
  );
  assign io_in_req_ready = arb_io_in_1_ready; // @[src/main/scala/nutcore/mem/Cache.scala 494:28]
  assign io_in_resp_valid = s3_io_out_valid & _io_in_resp_valid_T ? 1'h0 : s3_io_out_valid | s3_io_dataReadRespToL1; // @[src/main/scala/nutcore/mem/Cache.scala 510:26]
  assign io_in_resp_bits_cmd = s3_io_out_bits_cmd; // @[src/main/scala/nutcore/mem/Cache.scala 504:14]
  assign io_in_resp_bits_rdata = s3_io_out_bits_rdata; // @[src/main/scala/nutcore/mem/Cache.scala 504:14]
  assign io_out_mem_req_valid = s3_io_mem_req_valid; // @[src/main/scala/nutcore/mem/Cache.scala 506:14]
  assign io_out_mem_req_bits_addr = s3_io_mem_req_bits_addr; // @[src/main/scala/nutcore/mem/Cache.scala 506:14]
  assign io_out_mem_req_bits_cmd = s3_io_mem_req_bits_cmd; // @[src/main/scala/nutcore/mem/Cache.scala 506:14]
  assign io_out_mem_req_bits_wdata = s3_io_mem_req_bits_wdata; // @[src/main/scala/nutcore/mem/Cache.scala 506:14]
  assign s1_clock = clock;
  assign s1_reset = reset;
  assign s1_io_in_valid = arb_io_out_valid; // @[src/main/scala/nutcore/mem/Cache.scala 496:12]
  assign s1_io_in_bits_addr = arb_io_out_bits_addr; // @[src/main/scala/nutcore/mem/Cache.scala 496:12]
  assign s1_io_in_bits_size = arb_io_out_bits_size; // @[src/main/scala/nutcore/mem/Cache.scala 496:12]
  assign s1_io_in_bits_cmd = arb_io_out_bits_cmd; // @[src/main/scala/nutcore/mem/Cache.scala 496:12]
  assign s1_io_in_bits_wmask = arb_io_out_bits_wmask; // @[src/main/scala/nutcore/mem/Cache.scala 496:12]
  assign s1_io_in_bits_wdata = arb_io_out_bits_wdata; // @[src/main/scala/nutcore/mem/Cache.scala 496:12]
  assign s1_io_out_ready = s2_io_in_ready; // @[src/main/scala/utils/Pipeline.scala 29:16]
  assign s1_io_metaReadBus_req_ready = metaArray_io_r_0_req_ready; // @[src/main/scala/nutcore/mem/Cache.scala 528:21]
  assign s1_io_metaReadBus_resp_data_0_tag = metaArray_io_r_0_resp_data_0_tag; // @[src/main/scala/nutcore/mem/Cache.scala 528:21]
  assign s1_io_metaReadBus_resp_data_0_valid = metaArray_io_r_0_resp_data_0_valid; // @[src/main/scala/nutcore/mem/Cache.scala 528:21]
  assign s1_io_metaReadBus_resp_data_0_dirty = metaArray_io_r_0_resp_data_0_dirty; // @[src/main/scala/nutcore/mem/Cache.scala 528:21]
  assign s1_io_metaReadBus_resp_data_1_tag = metaArray_io_r_0_resp_data_1_tag; // @[src/main/scala/nutcore/mem/Cache.scala 528:21]
  assign s1_io_metaReadBus_resp_data_1_valid = metaArray_io_r_0_resp_data_1_valid; // @[src/main/scala/nutcore/mem/Cache.scala 528:21]
  assign s1_io_metaReadBus_resp_data_1_dirty = metaArray_io_r_0_resp_data_1_dirty; // @[src/main/scala/nutcore/mem/Cache.scala 528:21]
  assign s1_io_metaReadBus_resp_data_2_tag = metaArray_io_r_0_resp_data_2_tag; // @[src/main/scala/nutcore/mem/Cache.scala 528:21]
  assign s1_io_metaReadBus_resp_data_2_valid = metaArray_io_r_0_resp_data_2_valid; // @[src/main/scala/nutcore/mem/Cache.scala 528:21]
  assign s1_io_metaReadBus_resp_data_2_dirty = metaArray_io_r_0_resp_data_2_dirty; // @[src/main/scala/nutcore/mem/Cache.scala 528:21]
  assign s1_io_metaReadBus_resp_data_3_tag = metaArray_io_r_0_resp_data_3_tag; // @[src/main/scala/nutcore/mem/Cache.scala 528:21]
  assign s1_io_metaReadBus_resp_data_3_valid = metaArray_io_r_0_resp_data_3_valid; // @[src/main/scala/nutcore/mem/Cache.scala 528:21]
  assign s1_io_metaReadBus_resp_data_3_dirty = metaArray_io_r_0_resp_data_3_dirty; // @[src/main/scala/nutcore/mem/Cache.scala 528:21]
  assign s1_io_dataReadBus_req_ready = dataArray_io_r_0_req_ready; // @[src/main/scala/nutcore/mem/Cache.scala 529:21]
  assign s1_io_dataReadBus_resp_data_0_data = dataArray_io_r_0_resp_data_0_data; // @[src/main/scala/nutcore/mem/Cache.scala 529:21]
  assign s1_io_dataReadBus_resp_data_1_data = dataArray_io_r_0_resp_data_1_data; // @[src/main/scala/nutcore/mem/Cache.scala 529:21]
  assign s1_io_dataReadBus_resp_data_2_data = dataArray_io_r_0_resp_data_2_data; // @[src/main/scala/nutcore/mem/Cache.scala 529:21]
  assign s1_io_dataReadBus_resp_data_3_data = dataArray_io_r_0_resp_data_3_data; // @[src/main/scala/nutcore/mem/Cache.scala 529:21]
  assign s1_DISPLAY_ENABLE = DISPLAY_ENABLE;
  assign s2_clock = clock;
  assign s2_reset = reset;
  assign s2_io_in_valid = valid; // @[src/main/scala/utils/Pipeline.scala 31:17]
  assign s2_io_in_bits_req_addr = s2_io_in_bits_r_req_addr; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign s2_io_in_bits_req_size = s2_io_in_bits_r_req_size; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign s2_io_in_bits_req_cmd = s2_io_in_bits_r_req_cmd; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign s2_io_in_bits_req_wmask = s2_io_in_bits_r_req_wmask; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign s2_io_in_bits_req_wdata = s2_io_in_bits_r_req_wdata; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign s2_io_out_ready = s3_io_in_ready; // @[src/main/scala/utils/Pipeline.scala 29:16]
  assign s2_io_metaReadResp_0_tag = s1_io_metaReadBus_resp_data_0_tag; // @[src/main/scala/nutcore/mem/Cache.scala 535:22]
  assign s2_io_metaReadResp_0_valid = s1_io_metaReadBus_resp_data_0_valid; // @[src/main/scala/nutcore/mem/Cache.scala 535:22]
  assign s2_io_metaReadResp_0_dirty = s1_io_metaReadBus_resp_data_0_dirty; // @[src/main/scala/nutcore/mem/Cache.scala 535:22]
  assign s2_io_metaReadResp_1_tag = s1_io_metaReadBus_resp_data_1_tag; // @[src/main/scala/nutcore/mem/Cache.scala 535:22]
  assign s2_io_metaReadResp_1_valid = s1_io_metaReadBus_resp_data_1_valid; // @[src/main/scala/nutcore/mem/Cache.scala 535:22]
  assign s2_io_metaReadResp_1_dirty = s1_io_metaReadBus_resp_data_1_dirty; // @[src/main/scala/nutcore/mem/Cache.scala 535:22]
  assign s2_io_metaReadResp_2_tag = s1_io_metaReadBus_resp_data_2_tag; // @[src/main/scala/nutcore/mem/Cache.scala 535:22]
  assign s2_io_metaReadResp_2_valid = s1_io_metaReadBus_resp_data_2_valid; // @[src/main/scala/nutcore/mem/Cache.scala 535:22]
  assign s2_io_metaReadResp_2_dirty = s1_io_metaReadBus_resp_data_2_dirty; // @[src/main/scala/nutcore/mem/Cache.scala 535:22]
  assign s2_io_metaReadResp_3_tag = s1_io_metaReadBus_resp_data_3_tag; // @[src/main/scala/nutcore/mem/Cache.scala 535:22]
  assign s2_io_metaReadResp_3_valid = s1_io_metaReadBus_resp_data_3_valid; // @[src/main/scala/nutcore/mem/Cache.scala 535:22]
  assign s2_io_metaReadResp_3_dirty = s1_io_metaReadBus_resp_data_3_dirty; // @[src/main/scala/nutcore/mem/Cache.scala 535:22]
  assign s2_io_dataReadResp_0_data = s1_io_dataReadBus_resp_data_0_data; // @[src/main/scala/nutcore/mem/Cache.scala 536:22]
  assign s2_io_dataReadResp_1_data = s1_io_dataReadBus_resp_data_1_data; // @[src/main/scala/nutcore/mem/Cache.scala 536:22]
  assign s2_io_dataReadResp_2_data = s1_io_dataReadBus_resp_data_2_data; // @[src/main/scala/nutcore/mem/Cache.scala 536:22]
  assign s2_io_dataReadResp_3_data = s1_io_dataReadBus_resp_data_3_data; // @[src/main/scala/nutcore/mem/Cache.scala 536:22]
  assign s2_io_metaWriteBus_req_valid = s3_io_metaWriteBus_req_valid; // @[src/main/scala/nutcore/mem/Cache.scala 538:22]
  assign s2_io_metaWriteBus_req_bits_setIdx = s3_io_metaWriteBus_req_bits_setIdx; // @[src/main/scala/nutcore/mem/Cache.scala 538:22]
  assign s2_io_metaWriteBus_req_bits_data_tag = s3_io_metaWriteBus_req_bits_data_tag; // @[src/main/scala/nutcore/mem/Cache.scala 538:22]
  assign s2_io_metaWriteBus_req_bits_data_dirty = s3_io_metaWriteBus_req_bits_data_dirty; // @[src/main/scala/nutcore/mem/Cache.scala 538:22]
  assign s2_io_metaWriteBus_req_bits_waymask = s3_io_metaWriteBus_req_bits_waymask; // @[src/main/scala/nutcore/mem/Cache.scala 538:22]
  assign s2_io_dataWriteBus_req_valid = s3_io_dataWriteBus_req_valid; // @[src/main/scala/nutcore/mem/Cache.scala 537:22]
  assign s2_io_dataWriteBus_req_bits_setIdx = s3_io_dataWriteBus_req_bits_setIdx; // @[src/main/scala/nutcore/mem/Cache.scala 537:22]
  assign s2_io_dataWriteBus_req_bits_data_data = s3_io_dataWriteBus_req_bits_data_data; // @[src/main/scala/nutcore/mem/Cache.scala 537:22]
  assign s2_io_dataWriteBus_req_bits_waymask = s3_io_dataWriteBus_req_bits_waymask; // @[src/main/scala/nutcore/mem/Cache.scala 537:22]
  assign s2_DISPLAY_ENABLE = DISPLAY_ENABLE;
  assign s3_clock = clock;
  assign s3_reset = reset;
  assign s3_io_in_valid = valid_1; // @[src/main/scala/utils/Pipeline.scala 31:17]
  assign s3_io_in_bits_req_addr = s3_io_in_bits_r_req_addr; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign s3_io_in_bits_req_size = s3_io_in_bits_r_req_size; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign s3_io_in_bits_req_cmd = s3_io_in_bits_r_req_cmd; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign s3_io_in_bits_req_wmask = s3_io_in_bits_r_req_wmask; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign s3_io_in_bits_req_wdata = s3_io_in_bits_r_req_wdata; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign s3_io_in_bits_metas_0_tag = s3_io_in_bits_r_metas_0_tag; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign s3_io_in_bits_metas_0_valid = s3_io_in_bits_r_metas_0_valid; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign s3_io_in_bits_metas_0_dirty = s3_io_in_bits_r_metas_0_dirty; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign s3_io_in_bits_metas_1_tag = s3_io_in_bits_r_metas_1_tag; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign s3_io_in_bits_metas_1_valid = s3_io_in_bits_r_metas_1_valid; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign s3_io_in_bits_metas_1_dirty = s3_io_in_bits_r_metas_1_dirty; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign s3_io_in_bits_metas_2_tag = s3_io_in_bits_r_metas_2_tag; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign s3_io_in_bits_metas_2_valid = s3_io_in_bits_r_metas_2_valid; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign s3_io_in_bits_metas_2_dirty = s3_io_in_bits_r_metas_2_dirty; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign s3_io_in_bits_metas_3_tag = s3_io_in_bits_r_metas_3_tag; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign s3_io_in_bits_metas_3_valid = s3_io_in_bits_r_metas_3_valid; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign s3_io_in_bits_metas_3_dirty = s3_io_in_bits_r_metas_3_dirty; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign s3_io_in_bits_datas_0_data = s3_io_in_bits_r_datas_0_data; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign s3_io_in_bits_datas_1_data = s3_io_in_bits_r_datas_1_data; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign s3_io_in_bits_datas_2_data = s3_io_in_bits_r_datas_2_data; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign s3_io_in_bits_datas_3_data = s3_io_in_bits_r_datas_3_data; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign s3_io_in_bits_hit = s3_io_in_bits_r_hit; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign s3_io_in_bits_waymask = s3_io_in_bits_r_waymask; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign s3_io_in_bits_mmio = s3_io_in_bits_r_mmio; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign s3_io_in_bits_isForwardData = s3_io_in_bits_r_isForwardData; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign s3_io_in_bits_forwardData_data_data = s3_io_in_bits_r_forwardData_data_data; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign s3_io_in_bits_forwardData_waymask = s3_io_in_bits_r_forwardData_waymask; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign s3_io_out_ready = 1'h1; // @[src/main/scala/nutcore/mem/Cache.scala 504:14]
  assign s3_io_dataReadBus_req_ready = dataArray_io_r_1_req_ready; // @[src/main/scala/nutcore/mem/Cache.scala 530:21]
  assign s3_io_dataReadBus_resp_data_0_data = dataArray_io_r_1_resp_data_0_data; // @[src/main/scala/nutcore/mem/Cache.scala 530:21]
  assign s3_io_dataReadBus_resp_data_1_data = dataArray_io_r_1_resp_data_1_data; // @[src/main/scala/nutcore/mem/Cache.scala 530:21]
  assign s3_io_dataReadBus_resp_data_2_data = dataArray_io_r_1_resp_data_2_data; // @[src/main/scala/nutcore/mem/Cache.scala 530:21]
  assign s3_io_dataReadBus_resp_data_3_data = dataArray_io_r_1_resp_data_3_data; // @[src/main/scala/nutcore/mem/Cache.scala 530:21]
  assign s3_io_mem_req_ready = io_out_mem_req_ready; // @[src/main/scala/nutcore/mem/Cache.scala 506:14]
  assign s3_io_mem_resp_valid = io_out_mem_resp_valid; // @[src/main/scala/nutcore/mem/Cache.scala 506:14]
  assign s3_io_mem_resp_bits_cmd = io_out_mem_resp_bits_cmd; // @[src/main/scala/nutcore/mem/Cache.scala 506:14]
  assign s3_io_mem_resp_bits_rdata = io_out_mem_resp_bits_rdata; // @[src/main/scala/nutcore/mem/Cache.scala 506:14]
  assign s3_DISPLAY_ENABLE = DISPLAY_ENABLE;
  assign metaArray_clock = clock;
  assign metaArray_reset = reset;
  assign metaArray_io_r_0_req_valid = s1_io_metaReadBus_req_valid; // @[src/main/scala/nutcore/mem/Cache.scala 528:21]
  assign metaArray_io_r_0_req_bits_setIdx = s1_io_metaReadBus_req_bits_setIdx; // @[src/main/scala/nutcore/mem/Cache.scala 528:21]
  assign metaArray_io_w_req_valid = s3_io_metaWriteBus_req_valid; // @[src/main/scala/nutcore/mem/Cache.scala 532:18]
  assign metaArray_io_w_req_bits_setIdx = s3_io_metaWriteBus_req_bits_setIdx; // @[src/main/scala/nutcore/mem/Cache.scala 532:18]
  assign metaArray_io_w_req_bits_data_tag = s3_io_metaWriteBus_req_bits_data_tag; // @[src/main/scala/nutcore/mem/Cache.scala 532:18]
  assign metaArray_io_w_req_bits_data_dirty = s3_io_metaWriteBus_req_bits_data_dirty; // @[src/main/scala/nutcore/mem/Cache.scala 532:18]
  assign metaArray_io_w_req_bits_waymask = s3_io_metaWriteBus_req_bits_waymask; // @[src/main/scala/nutcore/mem/Cache.scala 532:18]
  assign dataArray_clock = clock;
  assign dataArray_reset = reset;
  assign dataArray_io_r_0_req_valid = s1_io_dataReadBus_req_valid; // @[src/main/scala/nutcore/mem/Cache.scala 529:21]
  assign dataArray_io_r_0_req_bits_setIdx = s1_io_dataReadBus_req_bits_setIdx; // @[src/main/scala/nutcore/mem/Cache.scala 529:21]
  assign dataArray_io_r_1_req_valid = s3_io_dataReadBus_req_valid; // @[src/main/scala/nutcore/mem/Cache.scala 530:21]
  assign dataArray_io_r_1_req_bits_setIdx = s3_io_dataReadBus_req_bits_setIdx; // @[src/main/scala/nutcore/mem/Cache.scala 530:21]
  assign dataArray_io_w_req_valid = s3_io_dataWriteBus_req_valid; // @[src/main/scala/nutcore/mem/Cache.scala 533:18]
  assign dataArray_io_w_req_bits_setIdx = s3_io_dataWriteBus_req_bits_setIdx; // @[src/main/scala/nutcore/mem/Cache.scala 533:18]
  assign dataArray_io_w_req_bits_data_data = s3_io_dataWriteBus_req_bits_data_data; // @[src/main/scala/nutcore/mem/Cache.scala 533:18]
  assign dataArray_io_w_req_bits_waymask = s3_io_dataWriteBus_req_bits_waymask; // @[src/main/scala/nutcore/mem/Cache.scala 533:18]
  assign arb_io_in_0_valid = 1'h0; // @[src/main/scala/nutcore/mem/Cache.scala 518:24]
  assign arb_io_in_0_bits_addr = 32'h0; // @[src/main/scala/nutcore/mem/Cache.scala 515:19 src/main/scala/bus/simplebus/SimpleBus.scala 64:15]
  assign arb_io_in_0_bits_size = 3'h0; // @[src/main/scala/nutcore/mem/Cache.scala 515:19 src/main/scala/bus/simplebus/SimpleBus.scala 66:15]
  assign arb_io_in_0_bits_cmd = 4'h0; // @[src/main/scala/nutcore/mem/Cache.scala 515:19 src/main/scala/bus/simplebus/SimpleBus.scala 65:14]
  assign arb_io_in_0_bits_wmask = 8'h0; // @[src/main/scala/nutcore/mem/Cache.scala 515:19 src/main/scala/bus/simplebus/SimpleBus.scala 68:16]
  assign arb_io_in_0_bits_wdata = 64'h0; // @[src/main/scala/nutcore/mem/Cache.scala 515:19 src/main/scala/bus/simplebus/SimpleBus.scala 67:16]
  assign arb_io_in_1_valid = io_in_req_valid; // @[src/main/scala/nutcore/mem/Cache.scala 494:28]
  assign arb_io_in_1_bits_addr = io_in_req_bits_addr; // @[src/main/scala/nutcore/mem/Cache.scala 494:28]
  assign arb_io_in_1_bits_size = io_in_req_bits_size; // @[src/main/scala/nutcore/mem/Cache.scala 494:28]
  assign arb_io_in_1_bits_cmd = io_in_req_bits_cmd; // @[src/main/scala/nutcore/mem/Cache.scala 494:28]
  assign arb_io_in_1_bits_wmask = io_in_req_bits_wmask; // @[src/main/scala/nutcore/mem/Cache.scala 494:28]
  assign arb_io_in_1_bits_wdata = io_in_req_bits_wdata; // @[src/main/scala/nutcore/mem/Cache.scala 494:28]
  assign arb_io_out_ready = s1_io_in_ready; // @[src/main/scala/nutcore/mem/Cache.scala 496:12]
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/utils/Pipeline.scala 24:24]
      valid <= 1'h0; // @[src/main/scala/utils/Pipeline.scala 24:24]
    end else begin
      valid <= _GEN_1;
    end
    if (_T_2) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      s2_io_in_bits_r_req_addr <= s1_io_out_bits_req_addr; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_2) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      s2_io_in_bits_r_req_size <= s1_io_out_bits_req_size; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_2) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      s2_io_in_bits_r_req_cmd <= s1_io_out_bits_req_cmd; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_2) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      s2_io_in_bits_r_req_wmask <= s1_io_out_bits_req_wmask; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_2) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      s2_io_in_bits_r_req_wdata <= s1_io_out_bits_req_wdata; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (reset) begin // @[src/main/scala/utils/Pipeline.scala 24:24]
      valid_1 <= 1'h0; // @[src/main/scala/utils/Pipeline.scala 24:24]
    end else begin
      valid_1 <= _GEN_9;
    end
    if (_T_4) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      s3_io_in_bits_r_req_addr <= s2_io_out_bits_req_addr; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_4) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      s3_io_in_bits_r_req_size <= s2_io_out_bits_req_size; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_4) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      s3_io_in_bits_r_req_cmd <= s2_io_out_bits_req_cmd; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_4) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      s3_io_in_bits_r_req_wmask <= s2_io_out_bits_req_wmask; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_4) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      s3_io_in_bits_r_req_wdata <= s2_io_out_bits_req_wdata; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_4) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      s3_io_in_bits_r_metas_0_tag <= s2_io_out_bits_metas_0_tag; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_4) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      s3_io_in_bits_r_metas_0_valid <= s2_io_out_bits_metas_0_valid; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_4) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      s3_io_in_bits_r_metas_0_dirty <= s2_io_out_bits_metas_0_dirty; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_4) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      s3_io_in_bits_r_metas_1_tag <= s2_io_out_bits_metas_1_tag; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_4) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      s3_io_in_bits_r_metas_1_valid <= s2_io_out_bits_metas_1_valid; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_4) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      s3_io_in_bits_r_metas_1_dirty <= s2_io_out_bits_metas_1_dirty; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_4) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      s3_io_in_bits_r_metas_2_tag <= s2_io_out_bits_metas_2_tag; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_4) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      s3_io_in_bits_r_metas_2_valid <= s2_io_out_bits_metas_2_valid; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_4) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      s3_io_in_bits_r_metas_2_dirty <= s2_io_out_bits_metas_2_dirty; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_4) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      s3_io_in_bits_r_metas_3_tag <= s2_io_out_bits_metas_3_tag; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_4) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      s3_io_in_bits_r_metas_3_valid <= s2_io_out_bits_metas_3_valid; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_4) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      s3_io_in_bits_r_metas_3_dirty <= s2_io_out_bits_metas_3_dirty; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_4) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      s3_io_in_bits_r_datas_0_data <= s2_io_out_bits_datas_0_data; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_4) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      s3_io_in_bits_r_datas_1_data <= s2_io_out_bits_datas_1_data; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_4) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      s3_io_in_bits_r_datas_2_data <= s2_io_out_bits_datas_2_data; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_4) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      s3_io_in_bits_r_datas_3_data <= s2_io_out_bits_datas_3_data; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_4) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      s3_io_in_bits_r_hit <= s2_io_out_bits_hit; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_4) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      s3_io_in_bits_r_waymask <= s2_io_out_bits_waymask; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_4) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      s3_io_in_bits_r_mmio <= s2_io_out_bits_mmio; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_4) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      s3_io_in_bits_r_isForwardData <= s2_io_out_bits_isForwardData; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_4) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      s3_io_in_bits_r_forwardData_data_data <= s2_io_out_bits_forwardData_data_data; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_4) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      s3_io_in_bits_r_forwardData_waymask <= s2_io_out_bits_forwardData_waymask; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (reset) begin // @[src/main/scala/utils/GTimer.scala 24:20]
      c <= 64'h0; // @[src/main/scala/utils/GTimer.scala 24:20]
    end else begin
      c <= _c_T_1; // @[src/main/scala/utils/GTimer.scala 25:7]
    end
    if (reset) begin // @[src/main/scala/utils/GTimer.scala 24:20]
      c_1 <= 64'h0; // @[src/main/scala/utils/GTimer.scala 24:20]
    end else begin
      c_1 <= _c_T_3; // @[src/main/scala/utils/GTimer.scala 25:7]
    end
    if (reset) begin // @[src/main/scala/utils/GTimer.scala 24:20]
      c_2 <= 64'h0; // @[src/main/scala/utils/GTimer.scala 24:20]
    end else begin
      c_2 <= _c_T_5; // @[src/main/scala/utils/GTimer.scala 25:7]
    end
    if (reset) begin // @[src/main/scala/utils/GTimer.scala 24:20]
      c_3 <= 64'h0; // @[src/main/scala/utils/GTimer.scala 24:20]
    end else begin
      c_3 <= _c_T_7; // @[src/main/scala/utils/GTimer.scala 25:7]
    end
    if (reset) begin // @[src/main/scala/utils/GTimer.scala 24:20]
      c_4 <= 64'h0; // @[src/main/scala/utils/GTimer.scala 24:20]
    end else begin
      c_4 <= _c_T_9; // @[src/main/scala/utils/GTimer.scala 25:7]
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & ~reset) begin
          $fwrite(32'h80000002,"[%d] Cache_2: ",c); // @[src/main/scala/utils/Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_7) begin
          $fwrite(32'h80000002,"InReq(%d, %d) InResp(%d, %d) \n",io_in_req_valid,io_in_req_ready,io_in_resp_valid,1'h1); // @[src/main/scala/utils/Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & ~reset) begin
          $fwrite(32'h80000002,"[%d] Cache_2: ",c_1); // @[src/main/scala/utils/Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_7) begin
          $fwrite(32'h80000002,"{IN s1:(%d,%d), s2:(%d,%d), s3:(%d,%d)} {OUT s1:(%d,%d), s2:(%d,%d), s3:(%d,%d)}\n",
            s1_io_in_valid,s1_io_in_ready,s2_io_in_valid,s2_io_in_ready,s3_io_in_valid,s3_io_in_ready,s1_io_out_valid,
            s1_io_out_ready,s2_io_out_valid,s2_io_out_ready,s3_io_out_valid,s3_io_out_ready); // @[src/main/scala/utils/Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (s1_io_in_valid & DISPLAY_ENABLE & ~reset) begin
          $fwrite(32'h80000002,"[%d] Cache_2: ",c_2); // @[src/main/scala/utils/Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_39 & _T_7) begin
          $fwrite(32'h80000002,"[l2cache.S1]: addr = 0x%x, cmd = %d, size = %d, wmask = 0x%x, wdata = 0x%x\n",
            s1_io_in_bits_addr,s1_io_in_bits_cmd,s1_io_in_bits_size,s1_io_in_bits_wmask,s1_io_in_bits_wdata); // @[src/main/scala/utils/Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (s2_io_in_valid & DISPLAY_ENABLE & ~reset) begin
          $fwrite(32'h80000002,"[%d] Cache_2: ",c_3); // @[src/main/scala/utils/Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_41 & _T_7) begin
          $fwrite(32'h80000002,"[l2cache.S2]: addr = 0x%x, cmd = %d, size = %d, wmask = 0x%x, wdata = 0x%x\n",
            s2_io_in_bits_req_addr,s2_io_in_bits_req_cmd,s2_io_in_bits_req_size,s2_io_in_bits_req_wmask,
            s2_io_in_bits_req_wdata); // @[src/main/scala/utils/Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (s3_io_in_valid & DISPLAY_ENABLE & ~reset) begin
          $fwrite(32'h80000002,"[%d] Cache_2: ",c_4); // @[src/main/scala/utils/Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_43 & _T_7) begin
          $fwrite(32'h80000002,"[l2cache.S3]: addr = 0x%x, cmd = %d, size = %d, wmask = 0x%x, wdata = 0x%x\n",
            s3_io_in_bits_req_addr,s3_io_in_bits_req_cmd,s3_io_in_bits_req_size,s3_io_in_bits_req_wmask,
            s3_io_in_bits_req_wdata); // @[src/main/scala/utils/Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  valid = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  s2_io_in_bits_r_req_addr = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  s2_io_in_bits_r_req_size = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  s2_io_in_bits_r_req_cmd = _RAND_3[3:0];
  _RAND_4 = {1{`RANDOM}};
  s2_io_in_bits_r_req_wmask = _RAND_4[7:0];
  _RAND_5 = {2{`RANDOM}};
  s2_io_in_bits_r_req_wdata = _RAND_5[63:0];
  _RAND_6 = {1{`RANDOM}};
  valid_1 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  s3_io_in_bits_r_req_addr = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  s3_io_in_bits_r_req_size = _RAND_8[2:0];
  _RAND_9 = {1{`RANDOM}};
  s3_io_in_bits_r_req_cmd = _RAND_9[3:0];
  _RAND_10 = {1{`RANDOM}};
  s3_io_in_bits_r_req_wmask = _RAND_10[7:0];
  _RAND_11 = {2{`RANDOM}};
  s3_io_in_bits_r_req_wdata = _RAND_11[63:0];
  _RAND_12 = {1{`RANDOM}};
  s3_io_in_bits_r_metas_0_tag = _RAND_12[16:0];
  _RAND_13 = {1{`RANDOM}};
  s3_io_in_bits_r_metas_0_valid = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  s3_io_in_bits_r_metas_0_dirty = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  s3_io_in_bits_r_metas_1_tag = _RAND_15[16:0];
  _RAND_16 = {1{`RANDOM}};
  s3_io_in_bits_r_metas_1_valid = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  s3_io_in_bits_r_metas_1_dirty = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  s3_io_in_bits_r_metas_2_tag = _RAND_18[16:0];
  _RAND_19 = {1{`RANDOM}};
  s3_io_in_bits_r_metas_2_valid = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  s3_io_in_bits_r_metas_2_dirty = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  s3_io_in_bits_r_metas_3_tag = _RAND_21[16:0];
  _RAND_22 = {1{`RANDOM}};
  s3_io_in_bits_r_metas_3_valid = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  s3_io_in_bits_r_metas_3_dirty = _RAND_23[0:0];
  _RAND_24 = {2{`RANDOM}};
  s3_io_in_bits_r_datas_0_data = _RAND_24[63:0];
  _RAND_25 = {2{`RANDOM}};
  s3_io_in_bits_r_datas_1_data = _RAND_25[63:0];
  _RAND_26 = {2{`RANDOM}};
  s3_io_in_bits_r_datas_2_data = _RAND_26[63:0];
  _RAND_27 = {2{`RANDOM}};
  s3_io_in_bits_r_datas_3_data = _RAND_27[63:0];
  _RAND_28 = {1{`RANDOM}};
  s3_io_in_bits_r_hit = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  s3_io_in_bits_r_waymask = _RAND_29[3:0];
  _RAND_30 = {1{`RANDOM}};
  s3_io_in_bits_r_mmio = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  s3_io_in_bits_r_isForwardData = _RAND_31[0:0];
  _RAND_32 = {2{`RANDOM}};
  s3_io_in_bits_r_forwardData_data_data = _RAND_32[63:0];
  _RAND_33 = {1{`RANDOM}};
  s3_io_in_bits_r_forwardData_waymask = _RAND_33[3:0];
  _RAND_34 = {2{`RANDOM}};
  c = _RAND_34[63:0];
  _RAND_35 = {2{`RANDOM}};
  c_1 = _RAND_35[63:0];
  _RAND_36 = {2{`RANDOM}};
  c_2 = _RAND_36[63:0];
  _RAND_37 = {2{`RANDOM}};
  c_3 = _RAND_37[63:0];
  _RAND_38 = {2{`RANDOM}};
  c_4 = _RAND_38[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module SimpleBusAddressMapper(
  output        io_in_req_ready, // @[src/main/scala/bus/simplebus/AddressMapper.scala 26:14]
  input         io_in_req_valid, // @[src/main/scala/bus/simplebus/AddressMapper.scala 26:14]
  input  [31:0] io_in_req_bits_addr, // @[src/main/scala/bus/simplebus/AddressMapper.scala 26:14]
  input  [3:0]  io_in_req_bits_cmd, // @[src/main/scala/bus/simplebus/AddressMapper.scala 26:14]
  input  [63:0] io_in_req_bits_wdata, // @[src/main/scala/bus/simplebus/AddressMapper.scala 26:14]
  output        io_in_resp_valid, // @[src/main/scala/bus/simplebus/AddressMapper.scala 26:14]
  output [3:0]  io_in_resp_bits_cmd, // @[src/main/scala/bus/simplebus/AddressMapper.scala 26:14]
  output [63:0] io_in_resp_bits_rdata, // @[src/main/scala/bus/simplebus/AddressMapper.scala 26:14]
  input         io_out_req_ready, // @[src/main/scala/bus/simplebus/AddressMapper.scala 26:14]
  output        io_out_req_valid, // @[src/main/scala/bus/simplebus/AddressMapper.scala 26:14]
  output [31:0] io_out_req_bits_addr, // @[src/main/scala/bus/simplebus/AddressMapper.scala 26:14]
  output [3:0]  io_out_req_bits_cmd, // @[src/main/scala/bus/simplebus/AddressMapper.scala 26:14]
  output [63:0] io_out_req_bits_wdata, // @[src/main/scala/bus/simplebus/AddressMapper.scala 26:14]
  input         io_out_resp_valid, // @[src/main/scala/bus/simplebus/AddressMapper.scala 26:14]
  input  [3:0]  io_out_resp_bits_cmd, // @[src/main/scala/bus/simplebus/AddressMapper.scala 26:14]
  input  [63:0] io_out_resp_bits_rdata // @[src/main/scala/bus/simplebus/AddressMapper.scala 26:14]
);
  assign io_in_req_ready = io_out_req_ready; // @[src/main/scala/bus/simplebus/AddressMapper.scala 31:10]
  assign io_in_resp_valid = io_out_resp_valid; // @[src/main/scala/bus/simplebus/AddressMapper.scala 31:10]
  assign io_in_resp_bits_cmd = io_out_resp_bits_cmd; // @[src/main/scala/bus/simplebus/AddressMapper.scala 31:10]
  assign io_in_resp_bits_rdata = io_out_resp_bits_rdata; // @[src/main/scala/bus/simplebus/AddressMapper.scala 31:10]
  assign io_out_req_valid = io_in_req_valid; // @[src/main/scala/bus/simplebus/AddressMapper.scala 31:10]
  assign io_out_req_bits_addr = io_in_req_bits_addr; // @[src/main/scala/bus/simplebus/AddressMapper.scala 31:10]
  assign io_out_req_bits_cmd = io_in_req_bits_cmd; // @[src/main/scala/bus/simplebus/AddressMapper.scala 31:10]
  assign io_out_req_bits_wdata = io_in_req_bits_wdata; // @[src/main/scala/bus/simplebus/AddressMapper.scala 31:10]
endmodule
module SimpleBus2AXI4Converter(
  input         clock,
  input         reset,
  output        io_in_req_ready, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input         io_in_req_valid, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input  [31:0] io_in_req_bits_addr, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input  [3:0]  io_in_req_bits_cmd, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input  [63:0] io_in_req_bits_wdata, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output        io_in_resp_valid, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output [3:0]  io_in_resp_bits_cmd, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output [63:0] io_in_resp_bits_rdata, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input         io_out_aw_ready, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output        io_out_aw_valid, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output [31:0] io_out_aw_bits_addr, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output [7:0]  io_out_aw_bits_len, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output [2:0]  io_out_aw_bits_size, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output [1:0]  io_out_aw_bits_burst, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input         io_out_w_ready, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output        io_out_w_valid, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output [63:0] io_out_w_bits_data, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output        io_out_w_bits_last, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input         io_out_b_valid, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input         io_out_ar_ready, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output        io_out_ar_valid, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output [31:0] io_out_ar_bits_addr, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output [7:0]  io_out_ar_bits_len, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output [2:0]  io_out_ar_bits_size, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output [1:0]  io_out_ar_bits_burst, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input         io_out_r_valid, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input  [63:0] io_out_r_bits_data, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input         io_out_r_bits_last // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  wire [2:0] _io_out_ar_bits_len_T_1 = io_in_req_bits_cmd[1] ? 3'h7 : 3'h0; // @[src/main/scala/bus/simplebus/ToAXI4.scala 169:30]
  wire  _io_out_w_bits_last_T = io_in_req_bits_cmd == 4'h7; // @[src/main/scala/bus/simplebus/SimpleBus.scala 78:27]
  wire  _io_out_w_bits_last_T_1 = io_in_req_bits_cmd == 4'h1; // @[src/main/scala/bus/simplebus/SimpleBus.scala 77:29]
  wire [2:0] _io_in_resp_bits_cmd_T = io_out_r_bits_last ? 3'h6 : 3'h0; // @[src/main/scala/bus/simplebus/ToAXI4.scala 184:28]
  wire  _awAck_T = io_out_aw_ready & io_out_aw_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  reg  awAck; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  _GEN_0 = _awAck_T | awAck; // @[src/main/scala/utils/StopWatch.scala 24:20 30:{20,24}]
  wire  _wSend_T_1 = io_out_w_ready & io_out_w_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  reg  wAck; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  wSend = _awAck_T & _wSend_T_1 & io_out_w_bits_last | awAck & wAck; // @[src/main/scala/bus/simplebus/ToAXI4.scala 189:49]
  wire  _wAck_T_1 = _wSend_T_1 & io_out_w_bits_last; // @[src/main/scala/bus/simplebus/ToAXI4.scala 188:39]
  wire  _GEN_2 = _wAck_T_1 | wAck; // @[src/main/scala/utils/StopWatch.scala 24:20 30:{20,24}]
  wire  _wen_T_1 = io_in_req_ready & io_in_req_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  reg  wen; // @[src/main/scala/bus/simplebus/ToAXI4.scala 190:22]
  wire  _io_out_ar_valid_T_4 = ~io_in_req_bits_cmd[0] & ~io_in_req_bits_cmd[3]; // @[src/main/scala/bus/simplebus/SimpleBus.scala 73:26]
  wire  _io_out_aw_valid_T_1 = io_in_req_valid & io_in_req_bits_cmd[0]; // @[src/main/scala/bus/simplebus/SimpleBus.scala 103:27]
  wire  _io_out_w_valid_T_2 = ~wAck; // @[src/main/scala/bus/simplebus/ToAXI4.scala 194:34]
  assign io_in_req_ready = io_in_req_bits_cmd[0] ? _io_out_w_valid_T_2 & io_out_w_ready : io_out_ar_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 195:24]
  assign io_in_resp_valid = wen ? io_out_b_valid : io_out_r_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 199:25]
  assign io_in_resp_bits_cmd = {{1'd0}, _io_in_resp_bits_cmd_T}; // @[src/main/scala/bus/simplebus/ToAXI4.scala 184:22]
  assign io_in_resp_bits_rdata = io_out_r_bits_data; // @[src/main/scala/bus/simplebus/ToAXI4.scala 183:23]
  assign io_out_aw_valid = _io_out_aw_valid_T_1 & ~awAck; // @[src/main/scala/bus/simplebus/ToAXI4.scala 193:31]
  assign io_out_aw_bits_addr = io_out_ar_bits_addr; // @[src/main/scala/bus/simplebus/ToAXI4.scala 182:6]
  assign io_out_aw_bits_len = io_out_ar_bits_len; // @[src/main/scala/bus/simplebus/ToAXI4.scala 182:6]
  assign io_out_aw_bits_size = io_out_ar_bits_size; // @[src/main/scala/bus/simplebus/ToAXI4.scala 182:6]
  assign io_out_aw_bits_burst = io_out_ar_bits_burst; // @[src/main/scala/bus/simplebus/ToAXI4.scala 182:6]
  assign io_out_w_valid = _io_out_aw_valid_T_1 & ~wAck; // @[src/main/scala/bus/simplebus/ToAXI4.scala 194:31]
  assign io_out_w_bits_data = io_in_req_bits_wdata; // @[src/main/scala/bus/simplebus/ToAXI4.scala 160:10]
  assign io_out_w_bits_last = _io_out_w_bits_last_T | _io_out_w_bits_last_T_1; // @[src/main/scala/bus/simplebus/ToAXI4.scala 177:54]
  assign io_out_ar_valid = io_in_req_valid & _io_out_ar_valid_T_4; // @[src/main/scala/bus/simplebus/SimpleBus.scala 104:27]
  assign io_out_ar_bits_addr = io_in_req_bits_addr; // @[src/main/scala/bus/simplebus/ToAXI4.scala 158:12]
  assign io_out_ar_bits_len = {{5'd0}, _io_out_ar_bits_len_T_1}; // @[src/main/scala/bus/simplebus/ToAXI4.scala 169:24]
  assign io_out_ar_bits_size = 3'h3; // @[src/main/scala/bus/simplebus/ToAXI4.scala 170:24]
  assign io_out_ar_bits_burst = 2'h2; // @[src/main/scala/bus/simplebus/ToAXI4.scala 171:24]
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      awAck <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else if (wSend) begin // @[src/main/scala/utils/StopWatch.scala 31:19]
      awAck <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 31:23]
    end else begin
      awAck <= _GEN_0;
    end
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      wAck <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else if (wSend) begin // @[src/main/scala/utils/StopWatch.scala 31:19]
      wAck <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 31:23]
    end else begin
      wAck <= _GEN_2;
    end
    if (_wen_T_1) begin // @[src/main/scala/bus/simplebus/ToAXI4.scala 190:22]
      wen <= io_in_req_bits_cmd[0]; // @[src/main/scala/bus/simplebus/ToAXI4.scala 190:22]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  awAck = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  wAck = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  wen = _RAND_2[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module SimpleBusCrossbar1toN(
  input         clock,
  input         reset,
  output        io_in_req_ready, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  input         io_in_req_valid, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  input  [31:0] io_in_req_bits_addr, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  input  [2:0]  io_in_req_bits_size, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  input  [3:0]  io_in_req_bits_cmd, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  input  [7:0]  io_in_req_bits_wmask, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  input  [63:0] io_in_req_bits_wdata, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output        io_in_resp_valid, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output [3:0]  io_in_resp_bits_cmd, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output [63:0] io_in_resp_bits_rdata, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  input         io_out_0_req_ready, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output        io_out_0_req_valid, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output [31:0] io_out_0_req_bits_addr, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output [3:0]  io_out_0_req_bits_cmd, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output [7:0]  io_out_0_req_bits_wmask, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output [63:0] io_out_0_req_bits_wdata, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output        io_out_0_resp_ready, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  input         io_out_0_resp_valid, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  input  [63:0] io_out_0_resp_bits_rdata, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  input         io_out_1_req_ready, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output        io_out_1_req_valid, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output [31:0] io_out_1_req_bits_addr, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output [3:0]  io_out_1_req_bits_cmd, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output [7:0]  io_out_1_req_bits_wmask, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output [63:0] io_out_1_req_bits_wdata, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output        io_out_1_resp_ready, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  input         io_out_1_resp_valid, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  input  [63:0] io_out_1_resp_bits_rdata, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  input         io_out_2_req_ready, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output        io_out_2_req_valid, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output [31:0] io_out_2_req_bits_addr, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output [2:0]  io_out_2_req_bits_size, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output [3:0]  io_out_2_req_bits_cmd, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output [7:0]  io_out_2_req_bits_wmask, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output [63:0] io_out_2_req_bits_wdata, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output        io_out_2_resp_ready, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  input         io_out_2_resp_valid, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  input  [3:0]  io_out_2_resp_bits_cmd, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  input  [63:0] io_out_2_resp_bits_rdata, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  input         DISPLAY_ENABLE
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
`endif // RANDOMIZE_REG_INIT
  reg [1:0] state; // @[src/main/scala/bus/simplebus/Crossbar.scala 32:22]
  wire  outMatchVec_0 = io_in_req_bits_addr >= 32'h38000000 & io_in_req_bits_addr < 32'h38010000; // @[src/main/scala/bus/simplebus/Crossbar.scala 37:34]
  wire  outMatchVec_1 = io_in_req_bits_addr >= 32'h3c000000 & io_in_req_bits_addr < 32'h40000000; // @[src/main/scala/bus/simplebus/Crossbar.scala 37:34]
  wire  outMatchVec_2 = io_in_req_bits_addr >= 32'h40000000 & io_in_req_bits_addr < 32'h80000000; // @[src/main/scala/bus/simplebus/Crossbar.scala 37:34]
  wire [2:0] _outSelVec_enc_T = outMatchVec_2 ? 3'h4 : 3'h0; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [2:0] _outSelVec_enc_T_1 = outMatchVec_1 ? 3'h2 : _outSelVec_enc_T; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [2:0] outSelVec_enc = outMatchVec_0 ? 3'h1 : _outSelVec_enc_T_1; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire  outSelVec_0 = outSelVec_enc[0]; // @[src/main/scala/chisel3/util/OneHot.scala 83:30]
  wire  outSelVec_1 = outSelVec_enc[1]; // @[src/main/scala/chisel3/util/OneHot.scala 83:30]
  wire  outSelVec_2 = outSelVec_enc[2]; // @[src/main/scala/chisel3/util/OneHot.scala 83:30]
  wire  _outSelRespVec_T = io_in_req_ready & io_in_req_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  wire  _outSelRespVec_T_1 = state == 2'h0; // @[src/main/scala/bus/simplebus/Crossbar.scala 41:57]
  wire  _outSelRespVec_T_2 = _outSelRespVec_T & state == 2'h0; // @[src/main/scala/bus/simplebus/Crossbar.scala 41:48]
  reg  outSelRespVec_0; // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
  reg  outSelRespVec_1; // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
  reg  outSelRespVec_2; // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
  wire [2:0] _reqInvalidAddr_T = {outSelVec_2,outSelVec_1,outSelVec_0}; // @[src/main/scala/bus/simplebus/Crossbar.scala 42:54]
  wire  reqInvalidAddr = io_in_req_valid & ~(|_reqInvalidAddr_T); // @[src/main/scala/bus/simplebus/Crossbar.scala 42:40]
  reg [63:0] c; // @[src/main/scala/utils/GTimer.scala 24:20]
  wire [63:0] _c_T_1 = c + 64'h1; // @[src/main/scala/utils/GTimer.scala 25:12]
  wire  _T_2 = ~reset; // @[src/main/scala/bus/simplebus/Crossbar.scala 46:13]
  wire [1:0] _GEN_5 = io_in_resp_valid ? 2'h0 : state; // @[src/main/scala/bus/simplebus/Crossbar.scala 32:22 56:{42,50}]
  wire  _io_in_req_ready_T_4 = outSelVec_0 & io_out_0_req_ready | outSelVec_1 & io_out_1_req_ready | outSelVec_2 &
    io_out_2_req_ready; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _io_in_resp_valid_T_4 = outSelRespVec_0 & io_out_0_resp_valid | outSelRespVec_1 & io_out_1_resp_valid |
    outSelRespVec_2 & io_out_2_resp_valid; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_in_resp_bits_T = outSelRespVec_0 ? io_out_0_resp_bits_rdata : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_in_resp_bits_T_1 = outSelRespVec_1 ? io_out_1_resp_bits_rdata : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_in_resp_bits_T_2 = outSelRespVec_2 ? io_out_2_resp_bits_rdata : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_in_resp_bits_T_3 = _io_in_resp_bits_T | _io_in_resp_bits_T_1; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [3:0] _io_in_resp_bits_T_5 = outSelRespVec_0 ? 4'h6 : 4'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [3:0] _io_in_resp_bits_T_6 = outSelRespVec_1 ? 4'h6 : 4'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [3:0] _io_in_resp_bits_T_7 = outSelRespVec_2 ? io_out_2_resp_bits_cmd : 4'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [3:0] _io_in_resp_bits_T_8 = _io_in_resp_bits_T_5 | _io_in_resp_bits_T_6; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  reg [63:0] c_1; // @[src/main/scala/utils/GTimer.scala 24:20]
  wire [63:0] _c_T_3 = c_1 + 64'h1; // @[src/main/scala/utils/GTimer.scala 25:12]
  reg [63:0] c_2; // @[src/main/scala/utils/GTimer.scala 24:20]
  wire [63:0] _c_T_5 = c_2 + 64'h1; // @[src/main/scala/utils/GTimer.scala 25:12]
  assign io_in_req_ready = _io_in_req_ready_T_4 | reqInvalidAddr; // @[src/main/scala/bus/simplebus/Crossbar.scala 61:64]
  assign io_in_resp_valid = _io_in_resp_valid_T_4 | state == 2'h2; // @[src/main/scala/bus/simplebus/Crossbar.scala 71:70]
  assign io_in_resp_bits_cmd = _io_in_resp_bits_T_8 | _io_in_resp_bits_T_7; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign io_in_resp_bits_rdata = _io_in_resp_bits_T_3 | _io_in_resp_bits_T_2; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign io_out_0_req_valid = outSelVec_0 & io_in_req_valid & _outSelRespVec_T_1; // @[src/main/scala/bus/simplebus/Crossbar.scala 63:60]
  assign io_out_0_req_bits_addr = io_in_req_bits_addr; // @[src/main/scala/bus/simplebus/Crossbar.scala 64:24]
  assign io_out_0_req_bits_cmd = io_in_req_bits_cmd; // @[src/main/scala/bus/simplebus/Crossbar.scala 64:24]
  assign io_out_0_req_bits_wmask = io_in_req_bits_wmask; // @[src/main/scala/bus/simplebus/Crossbar.scala 64:24]
  assign io_out_0_req_bits_wdata = io_in_req_bits_wdata; // @[src/main/scala/bus/simplebus/Crossbar.scala 64:24]
  assign io_out_0_resp_ready = outSelRespVec_0 & state == 2'h1; // @[src/main/scala/bus/simplebus/Crossbar.scala 69:66]
  assign io_out_1_req_valid = outSelVec_1 & io_in_req_valid & _outSelRespVec_T_1; // @[src/main/scala/bus/simplebus/Crossbar.scala 63:60]
  assign io_out_1_req_bits_addr = io_in_req_bits_addr; // @[src/main/scala/bus/simplebus/Crossbar.scala 64:24]
  assign io_out_1_req_bits_cmd = io_in_req_bits_cmd; // @[src/main/scala/bus/simplebus/Crossbar.scala 64:24]
  assign io_out_1_req_bits_wmask = io_in_req_bits_wmask; // @[src/main/scala/bus/simplebus/Crossbar.scala 64:24]
  assign io_out_1_req_bits_wdata = io_in_req_bits_wdata; // @[src/main/scala/bus/simplebus/Crossbar.scala 64:24]
  assign io_out_1_resp_ready = outSelRespVec_1 & state == 2'h1; // @[src/main/scala/bus/simplebus/Crossbar.scala 69:66]
  assign io_out_2_req_valid = outSelVec_2 & io_in_req_valid & _outSelRespVec_T_1; // @[src/main/scala/bus/simplebus/Crossbar.scala 63:60]
  assign io_out_2_req_bits_addr = io_in_req_bits_addr; // @[src/main/scala/bus/simplebus/Crossbar.scala 64:24]
  assign io_out_2_req_bits_size = io_in_req_bits_size; // @[src/main/scala/bus/simplebus/Crossbar.scala 64:24]
  assign io_out_2_req_bits_cmd = io_in_req_bits_cmd; // @[src/main/scala/bus/simplebus/Crossbar.scala 64:24]
  assign io_out_2_req_bits_wmask = io_in_req_bits_wmask; // @[src/main/scala/bus/simplebus/Crossbar.scala 64:24]
  assign io_out_2_req_bits_wdata = io_in_req_bits_wdata; // @[src/main/scala/bus/simplebus/Crossbar.scala 64:24]
  assign io_out_2_resp_ready = outSelRespVec_2 & state == 2'h1; // @[src/main/scala/bus/simplebus/Crossbar.scala 69:66]
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 32:22]
      state <= 2'h0; // @[src/main/scala/bus/simplebus/Crossbar.scala 32:22]
    end else if (2'h0 == state) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 51:18]
      if (reqInvalidAddr) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 54:29]
        state <= 2'h2; // @[src/main/scala/bus/simplebus/Crossbar.scala 54:37]
      end else if (_outSelRespVec_T) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 53:29]
        state <= 2'h1; // @[src/main/scala/bus/simplebus/Crossbar.scala 53:37]
      end
    end else if (2'h1 == state) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 51:18]
      state <= _GEN_5;
    end else if (2'h2 == state) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 51:18]
      state <= _GEN_5;
    end
    if (reset) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
      outSelRespVec_0 <= 1'h0; // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
    end else if (_outSelRespVec_T_2) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
      outSelRespVec_0 <= outSelVec_0; // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
    end
    if (reset) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
      outSelRespVec_1 <= 1'h0; // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
    end else if (_outSelRespVec_T_2) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
      outSelRespVec_1 <= outSelVec_1; // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
    end
    if (reset) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
      outSelRespVec_2 <= 1'h0; // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
    end else if (_outSelRespVec_T_2) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
      outSelRespVec_2 <= outSelVec_2; // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
    end
    if (reset) begin // @[src/main/scala/utils/GTimer.scala 24:20]
      c <= 64'h0; // @[src/main/scala/utils/GTimer.scala 24:20]
    end else begin
      c <= _c_T_1; // @[src/main/scala/utils/GTimer.scala 25:7]
    end
    if (reset) begin // @[src/main/scala/utils/GTimer.scala 24:20]
      c_1 <= 64'h0; // @[src/main/scala/utils/GTimer.scala 24:20]
    end else begin
      c_1 <= _c_T_3; // @[src/main/scala/utils/GTimer.scala 25:7]
    end
    if (reset) begin // @[src/main/scala/utils/GTimer.scala 24:20]
      c_2 <= 64'h0; // @[src/main/scala/utils/GTimer.scala 24:20]
    end else begin
      c_2 <= _c_T_5; // @[src/main/scala/utils/GTimer.scala 25:7]
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (reqInvalidAddr & DISPLAY_ENABLE & ~reset) begin
          $fwrite(32'h80000002,"crossbar access bad addr %x, time %d\n",io_in_req_bits_addr,c); // @[src/main/scala/bus/simplebus/Crossbar.scala 46:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2 & ~(~reqInvalidAddr)) begin
          $fwrite(32'h80000002,
            "Assertion failed: address decode error, bad addr = 0x%x\n\n    at Crossbar.scala:49 assert(!reqInvalidAddr, \"address decode error, bad addr = 0x%%%%x\\n\", addr)\n"
            ,io_in_req_bits_addr); // @[src/main/scala/bus/simplebus/Crossbar.scala 49:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~reqInvalidAddr) & _T_2) begin
          $fatal; // @[src/main/scala/bus/simplebus/Crossbar.scala 49:9]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _outSelRespVec_T & _T_2) begin
          $fwrite(32'h80000002,
            "%d: xbar: outSelVec = Vec(%d, %d, %d), outSel.req: addr = 0x%x, cmd = %d, size = %d, wmask = 0x%x, wdata = 0x%x\n"
            ,c_1,outSelVec_0,outSelVec_1,outSelVec_2,io_in_req_bits_addr,io_in_req_bits_cmd,io_in_req_bits_size,
            io_in_req_bits_wmask,io_in_req_bits_wdata); // @[src/main/scala/bus/simplebus/Crossbar.scala 77:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & io_in_resp_valid & _T_2) begin
          $fwrite(32'h80000002,"%d: xbar: outSelVec = Vec(%d, %d, %d), outSel.resp: rdata = %x, cmd = %d\n",c_2,
            outSelVec_0,outSelVec_1,outSelVec_2,io_in_resp_bits_rdata,io_in_resp_bits_cmd); // @[src/main/scala/bus/simplebus/Crossbar.scala 80:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  outSelRespVec_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  outSelRespVec_1 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  outSelRespVec_2 = _RAND_3[0:0];
  _RAND_4 = {2{`RANDOM}};
  c = _RAND_4[63:0];
  _RAND_5 = {2{`RANDOM}};
  c_1 = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  c_2 = _RAND_6[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module AXI4CLINT(
  input         clock,
  input         reset,
  output        io__in_aw_ready, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input         io__in_aw_valid, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input  [31:0] io__in_aw_bits_addr, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output        io__in_w_ready, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input         io__in_w_valid, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input  [63:0] io__in_w_bits_data, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input  [7:0]  io__in_w_bits_strb, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input         io__in_b_ready, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output        io__in_b_valid, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output        io__in_ar_ready, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input         io__in_ar_valid, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input  [31:0] io__in_ar_bits_addr, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input         io__in_r_ready, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output        io__in_r_valid, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output [63:0] io__in_r_bits_data, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output        io__extra_mtip, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output        io__extra_msip, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input         isWFI_0,
  output        io_extra_mtip,
  output        io_extra_msip
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
`endif // RANDOMIZE_REG_INIT
  wire [7:0] _fullMask_T_9 = io__in_w_bits_strb[0] ? 8'hff : 8'h0; // @[src/main/scala/utils/BitUtils.scala 27:45]
  wire [7:0] _fullMask_T_11 = io__in_w_bits_strb[1] ? 8'hff : 8'h0; // @[src/main/scala/utils/BitUtils.scala 27:45]
  wire [7:0] _fullMask_T_13 = io__in_w_bits_strb[2] ? 8'hff : 8'h0; // @[src/main/scala/utils/BitUtils.scala 27:45]
  wire [7:0] _fullMask_T_15 = io__in_w_bits_strb[3] ? 8'hff : 8'h0; // @[src/main/scala/utils/BitUtils.scala 27:45]
  wire [7:0] _fullMask_T_17 = io__in_w_bits_strb[4] ? 8'hff : 8'h0; // @[src/main/scala/utils/BitUtils.scala 27:45]
  wire [7:0] _fullMask_T_19 = io__in_w_bits_strb[5] ? 8'hff : 8'h0; // @[src/main/scala/utils/BitUtils.scala 27:45]
  wire [7:0] _fullMask_T_21 = io__in_w_bits_strb[6] ? 8'hff : 8'h0; // @[src/main/scala/utils/BitUtils.scala 27:45]
  wire [7:0] _fullMask_T_23 = io__in_w_bits_strb[7] ? 8'hff : 8'h0; // @[src/main/scala/utils/BitUtils.scala 27:45]
  wire [63:0] fullMask = {_fullMask_T_23,_fullMask_T_21,_fullMask_T_19,_fullMask_T_17,_fullMask_T_15,_fullMask_T_13,
    _fullMask_T_11,_fullMask_T_9}; // @[src/main/scala/utils/BitUtils.scala 27:26]
  wire  _r_busy_T = io__in_ar_ready & io__in_ar_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  wire  _r_busy_T_1 = io__in_r_ready & io__in_r_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  reg  r_busy; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  _GEN_0 = _r_busy_T_1 ? 1'h0 : r_busy; // @[src/main/scala/utils/StopWatch.scala 26:19 24:20 26:23]
  wire  _GEN_1 = _r_busy_T | _GEN_0; // @[src/main/scala/utils/StopWatch.scala 27:{20,24}]
  reg  ren_REG; // @[src/main/scala/device/AXI4Slave.scala 73:17]
  wire  _io_in_r_valid_T_2 = ren_REG & (_r_busy_T | r_busy); // @[src/main/scala/device/AXI4Slave.scala 74:35]
  reg  io_in_r_valid_r; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  _GEN_2 = _r_busy_T_1 ? 1'h0 : io_in_r_valid_r; // @[src/main/scala/utils/StopWatch.scala 26:19 24:20 26:23]
  wire  _GEN_3 = _io_in_r_valid_T_2 | _GEN_2; // @[src/main/scala/utils/StopWatch.scala 27:{20,24}]
  wire  _w_busy_T = io__in_aw_ready & io__in_aw_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  wire  _w_busy_T_1 = io__in_b_ready & io__in_b_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  reg  w_busy; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  _GEN_4 = _w_busy_T_1 ? 1'h0 : w_busy; // @[src/main/scala/utils/StopWatch.scala 26:19 24:20 26:23]
  wire  _GEN_5 = _w_busy_T | _GEN_4; // @[src/main/scala/utils/StopWatch.scala 27:{20,24}]
  wire  _io_in_b_valid_T = io__in_w_ready & io__in_w_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  reg  io_in_b_valid_r; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  _GEN_6 = _w_busy_T_1 ? 1'h0 : io_in_b_valid_r; // @[src/main/scala/utils/StopWatch.scala 26:19 24:20 26:23]
  wire  _GEN_7 = _io_in_b_valid_T | _GEN_6; // @[src/main/scala/utils/StopWatch.scala 27:{20,24}]
  reg [63:0] mtime; // @[src/main/scala/device/AXI4CLINT.scala 32:22]
  reg [63:0] mtimecmp; // @[src/main/scala/device/AXI4CLINT.scala 33:25]
  reg [63:0] msip; // @[src/main/scala/device/AXI4CLINT.scala 34:21]
  reg [63:0] freq_reg; // @[src/main/scala/device/AXI4CLINT.scala 37:25]
  wire [15:0] freq = freq_reg[15:0]; // @[src/main/scala/device/AXI4CLINT.scala 38:22]
  reg [63:0] inc_reg; // @[src/main/scala/device/AXI4CLINT.scala 39:24]
  wire [15:0] inc = inc_reg[15:0]; // @[src/main/scala/device/AXI4CLINT.scala 40:20]
  reg [15:0] cnt; // @[src/main/scala/device/AXI4CLINT.scala 42:20]
  wire [15:0] nextCnt = cnt + 16'h1; // @[src/main/scala/device/AXI4CLINT.scala 43:21]
  wire  tick = nextCnt == freq; // @[src/main/scala/device/AXI4CLINT.scala 45:23]
  wire [63:0] _GEN_15 = {{48'd0}, inc}; // @[src/main/scala/device/AXI4CLINT.scala 46:32]
  wire [63:0] _mtime_T_1 = mtime + _GEN_15; // @[src/main/scala/device/AXI4CLINT.scala 46:32]
  wire [63:0] _mtime_T_3 = mtime + 64'h186a0; // @[src/main/scala/device/AXI4CLINT.scala 51:35]
  wire  _io_in_r_bits_data_T = 16'h0 == io__in_ar_bits_addr[15:0]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _io_in_r_bits_data_T_1 = 16'h8000 == io__in_ar_bits_addr[15:0]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _io_in_r_bits_data_T_2 = 16'hbff8 == io__in_ar_bits_addr[15:0]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _io_in_r_bits_data_T_3 = 16'h8008 == io__in_ar_bits_addr[15:0]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _io_in_r_bits_data_T_4 = 16'h4000 == io__in_ar_bits_addr[15:0]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _io_in_r_bits_data_T_5 = _io_in_r_bits_data_T ? msip : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_in_r_bits_data_T_6 = _io_in_r_bits_data_T_1 ? freq_reg : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_in_r_bits_data_T_7 = _io_in_r_bits_data_T_2 ? mtime : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_in_r_bits_data_T_8 = _io_in_r_bits_data_T_3 ? inc_reg : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_in_r_bits_data_T_9 = _io_in_r_bits_data_T_4 ? mtimecmp : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_in_r_bits_data_T_10 = _io_in_r_bits_data_T_5 | _io_in_r_bits_data_T_6; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_in_r_bits_data_T_11 = _io_in_r_bits_data_T_10 | _io_in_r_bits_data_T_7; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_in_r_bits_data_T_12 = _io_in_r_bits_data_T_11 | _io_in_r_bits_data_T_8; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _msip_T = io__in_w_bits_data & fullMask; // @[src/main/scala/utils/BitUtils.scala 34:14]
  wire [63:0] _msip_T_1 = ~fullMask; // @[src/main/scala/utils/BitUtils.scala 34:39]
  wire [63:0] _msip_T_2 = msip & _msip_T_1; // @[src/main/scala/utils/BitUtils.scala 34:37]
  wire [63:0] _msip_T_3 = _msip_T | _msip_T_2; // @[src/main/scala/utils/BitUtils.scala 34:26]
  wire [63:0] _freq_reg_T_2 = freq_reg & _msip_T_1; // @[src/main/scala/utils/BitUtils.scala 34:37]
  wire [63:0] _freq_reg_T_3 = _msip_T | _freq_reg_T_2; // @[src/main/scala/utils/BitUtils.scala 34:26]
  wire [63:0] _mtime_T_6 = mtime & _msip_T_1; // @[src/main/scala/utils/BitUtils.scala 34:37]
  wire [63:0] _mtime_T_7 = _msip_T | _mtime_T_6; // @[src/main/scala/utils/BitUtils.scala 34:26]
  wire [63:0] _inc_reg_T_2 = inc_reg & _msip_T_1; // @[src/main/scala/utils/BitUtils.scala 34:37]
  wire [63:0] _inc_reg_T_3 = _msip_T | _inc_reg_T_2; // @[src/main/scala/utils/BitUtils.scala 34:26]
  wire [63:0] _mtimecmp_T_2 = mtimecmp & _msip_T_1; // @[src/main/scala/utils/BitUtils.scala 34:37]
  wire [63:0] _mtimecmp_T_3 = _msip_T | _mtimecmp_T_2; // @[src/main/scala/utils/BitUtils.scala 34:26]
  reg  io_extra_mtip_REG; // @[src/main/scala/device/AXI4CLINT.scala 66:31]
  reg  io_extra_msip_REG; // @[src/main/scala/device/AXI4CLINT.scala 67:31]
  assign io__in_aw_ready = ~w_busy; // @[src/main/scala/device/AXI4Slave.scala 94:18]
  assign io__in_w_ready = io__in_aw_valid | w_busy; // @[src/main/scala/device/AXI4Slave.scala 95:30]
  assign io__in_b_valid = io_in_b_valid_r; // @[src/main/scala/device/AXI4Slave.scala 97:14]
  assign io__in_ar_ready = io__in_r_ready | ~r_busy; // @[src/main/scala/device/AXI4Slave.scala 71:29]
  assign io__in_r_valid = io_in_r_valid_r; // @[src/main/scala/device/AXI4Slave.scala 74:14]
  assign io__in_r_bits_data = _io_in_r_bits_data_T_12 | _io_in_r_bits_data_T_9; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign io__extra_mtip = io_extra_mtip_REG; // @[src/main/scala/device/AXI4CLINT.scala 66:21]
  assign io__extra_msip = io_extra_msip_REG; // @[src/main/scala/device/AXI4CLINT.scala 67:21]
  assign io_extra_mtip = io__extra_mtip;
  assign io_extra_msip = io__extra_msip;
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      r_busy <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else begin
      r_busy <= _GEN_1;
    end
    if (reset) begin // @[src/main/scala/device/AXI4Slave.scala 73:17]
      ren_REG <= 1'h0; // @[src/main/scala/device/AXI4Slave.scala 73:17]
    end else begin
      ren_REG <= _r_busy_T; // @[src/main/scala/device/AXI4Slave.scala 73:17]
    end
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      io_in_r_valid_r <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else begin
      io_in_r_valid_r <= _GEN_3;
    end
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      w_busy <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else begin
      w_busy <= _GEN_5;
    end
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      io_in_b_valid_r <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else begin
      io_in_b_valid_r <= _GEN_7;
    end
    if (reset) begin // @[src/main/scala/device/AXI4CLINT.scala 32:22]
      mtime <= 64'h0; // @[src/main/scala/device/AXI4CLINT.scala 32:22]
    end else if (_io_in_b_valid_T & io__in_aw_bits_addr[15:0] == 16'hbff8) begin // @[src/main/scala/utils/RegMap.scala 32:48]
      mtime <= _mtime_T_7; // @[src/main/scala/utils/RegMap.scala 32:52]
    end else if (isWFI_0) begin // @[src/main/scala/device/AXI4CLINT.scala 51:18]
      mtime <= _mtime_T_3; // @[src/main/scala/device/AXI4CLINT.scala 51:26]
    end else if (tick) begin // @[src/main/scala/device/AXI4CLINT.scala 46:15]
      mtime <= _mtime_T_1; // @[src/main/scala/device/AXI4CLINT.scala 46:23]
    end
    if (reset) begin // @[src/main/scala/device/AXI4CLINT.scala 33:25]
      mtimecmp <= 64'h0; // @[src/main/scala/device/AXI4CLINT.scala 33:25]
    end else if (_io_in_b_valid_T & io__in_aw_bits_addr[15:0] == 16'h4000) begin // @[src/main/scala/utils/RegMap.scala 32:48]
      mtimecmp <= _mtimecmp_T_3; // @[src/main/scala/utils/RegMap.scala 32:52]
    end
    if (reset) begin // @[src/main/scala/device/AXI4CLINT.scala 34:21]
      msip <= 64'h0; // @[src/main/scala/device/AXI4CLINT.scala 34:21]
    end else if (_io_in_b_valid_T & io__in_aw_bits_addr[15:0] == 16'h0) begin // @[src/main/scala/utils/RegMap.scala 32:48]
      msip <= _msip_T_3; // @[src/main/scala/utils/RegMap.scala 32:52]
    end
    if (reset) begin // @[src/main/scala/device/AXI4CLINT.scala 37:25]
      freq_reg <= 64'h2710; // @[src/main/scala/device/AXI4CLINT.scala 37:25]
    end else if (_io_in_b_valid_T & io__in_aw_bits_addr[15:0] == 16'h8000) begin // @[src/main/scala/utils/RegMap.scala 32:48]
      freq_reg <= _freq_reg_T_3; // @[src/main/scala/utils/RegMap.scala 32:52]
    end
    if (reset) begin // @[src/main/scala/device/AXI4CLINT.scala 39:24]
      inc_reg <= 64'h1; // @[src/main/scala/device/AXI4CLINT.scala 39:24]
    end else if (_io_in_b_valid_T & io__in_aw_bits_addr[15:0] == 16'h8008) begin // @[src/main/scala/utils/RegMap.scala 32:48]
      inc_reg <= _inc_reg_T_3; // @[src/main/scala/utils/RegMap.scala 32:52]
    end
    if (reset) begin // @[src/main/scala/device/AXI4CLINT.scala 42:20]
      cnt <= 16'h0; // @[src/main/scala/device/AXI4CLINT.scala 42:20]
    end else if (nextCnt < freq) begin // @[src/main/scala/device/AXI4CLINT.scala 44:13]
      cnt <= nextCnt;
    end else begin
      cnt <= 16'h0;
    end
    io_extra_mtip_REG <= mtime >= mtimecmp; // @[src/main/scala/device/AXI4CLINT.scala 66:38]
    io_extra_msip_REG <= msip != 64'h0; // @[src/main/scala/device/AXI4CLINT.scala 67:37]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  r_busy = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  ren_REG = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  io_in_r_valid_r = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  w_busy = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  io_in_b_valid_r = _RAND_4[0:0];
  _RAND_5 = {2{`RANDOM}};
  mtime = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  mtimecmp = _RAND_6[63:0];
  _RAND_7 = {2{`RANDOM}};
  msip = _RAND_7[63:0];
  _RAND_8 = {2{`RANDOM}};
  freq_reg = _RAND_8[63:0];
  _RAND_9 = {2{`RANDOM}};
  inc_reg = _RAND_9[63:0];
  _RAND_10 = {1{`RANDOM}};
  cnt = _RAND_10[15:0];
  _RAND_11 = {1{`RANDOM}};
  io_extra_mtip_REG = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  io_extra_msip_REG = _RAND_12[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module SimpleBus2AXI4Converter_1(
  input         clock,
  input         reset,
  output        io_in_req_ready, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input         io_in_req_valid, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input  [31:0] io_in_req_bits_addr, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input  [3:0]  io_in_req_bits_cmd, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input  [7:0]  io_in_req_bits_wmask, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input  [63:0] io_in_req_bits_wdata, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input         io_in_resp_ready, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output        io_in_resp_valid, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output [63:0] io_in_resp_bits_rdata, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input         io_out_aw_ready, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output        io_out_aw_valid, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output [31:0] io_out_aw_bits_addr, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input         io_out_w_ready, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output        io_out_w_valid, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output [63:0] io_out_w_bits_data, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output [7:0]  io_out_w_bits_strb, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output        io_out_b_ready, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input         io_out_b_valid, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input         io_out_ar_ready, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output        io_out_ar_valid, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output [31:0] io_out_ar_bits_addr, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output        io_out_r_ready, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input         io_out_r_valid, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input  [63:0] io_out_r_bits_data // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  wire  toAXI4Lite = ~(io_in_req_valid & io_in_req_bits_cmd[1]); // @[src/main/scala/bus/simplebus/ToAXI4.scala 151:20]
  wire  _awAck_T = io_out_aw_ready & io_out_aw_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  reg  awAck; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  _GEN_0 = _awAck_T | awAck; // @[src/main/scala/utils/StopWatch.scala 24:20 30:{20,24}]
  wire  _wSend_T_1 = io_out_w_ready & io_out_w_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  reg  wAck; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  wSend = _awAck_T & _wSend_T_1 | awAck & wAck; // @[src/main/scala/bus/simplebus/ToAXI4.scala 189:49]
  wire  _GEN_2 = _wSend_T_1 | wAck; // @[src/main/scala/utils/StopWatch.scala 24:20 30:{20,24}]
  wire  _wen_T_1 = io_in_req_ready & io_in_req_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  reg  wen; // @[src/main/scala/bus/simplebus/ToAXI4.scala 190:22]
  wire  _io_out_ar_valid_T_4 = ~io_in_req_bits_cmd[0] & ~io_in_req_bits_cmd[3]; // @[src/main/scala/bus/simplebus/SimpleBus.scala 73:26]
  wire  _io_out_aw_valid_T_1 = io_in_req_valid & io_in_req_bits_cmd[0]; // @[src/main/scala/bus/simplebus/SimpleBus.scala 103:27]
  wire  _io_out_w_valid_T_2 = ~wAck; // @[src/main/scala/bus/simplebus/ToAXI4.scala 194:34]
  assign io_in_req_ready = io_in_req_bits_cmd[0] ? _io_out_w_valid_T_2 & io_out_w_ready : io_out_ar_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 195:24]
  assign io_in_resp_valid = wen ? io_out_b_valid : io_out_r_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 199:25]
  assign io_in_resp_bits_rdata = io_out_r_bits_data; // @[src/main/scala/bus/simplebus/ToAXI4.scala 183:23]
  assign io_out_aw_valid = _io_out_aw_valid_T_1 & ~awAck; // @[src/main/scala/bus/simplebus/ToAXI4.scala 193:31]
  assign io_out_aw_bits_addr = io_out_ar_bits_addr; // @[src/main/scala/bus/simplebus/ToAXI4.scala 182:6]
  assign io_out_w_valid = _io_out_aw_valid_T_1 & ~wAck; // @[src/main/scala/bus/simplebus/ToAXI4.scala 194:31]
  assign io_out_w_bits_data = io_in_req_bits_wdata; // @[src/main/scala/bus/simplebus/ToAXI4.scala 160:10]
  assign io_out_w_bits_strb = io_in_req_bits_wmask; // @[src/main/scala/bus/simplebus/ToAXI4.scala 161:10]
  assign io_out_b_ready = io_in_resp_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 198:16]
  assign io_out_ar_valid = io_in_req_valid & _io_out_ar_valid_T_4; // @[src/main/scala/bus/simplebus/SimpleBus.scala 104:27]
  assign io_out_ar_bits_addr = io_in_req_bits_addr; // @[src/main/scala/bus/simplebus/ToAXI4.scala 158:12]
  assign io_out_r_ready = io_in_resp_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 197:16]
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      awAck <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else if (wSend) begin // @[src/main/scala/utils/StopWatch.scala 31:19]
      awAck <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 31:23]
    end else begin
      awAck <= _GEN_0;
    end
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      wAck <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else if (wSend) begin // @[src/main/scala/utils/StopWatch.scala 31:19]
      wAck <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 31:23]
    end else begin
      wAck <= _GEN_2;
    end
    if (_wen_T_1) begin // @[src/main/scala/bus/simplebus/ToAXI4.scala 190:22]
      wen <= io_in_req_bits_cmd[0]; // @[src/main/scala/bus/simplebus/ToAXI4.scala 190:22]
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~toAXI4Lite) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:153 assert(toAXI4Lite || toAXI4)\n"); // @[src/main/scala/bus/simplebus/ToAXI4.scala 153:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~toAXI4Lite & ~reset) begin
          $fatal; // @[src/main/scala/bus/simplebus/ToAXI4.scala 153:9]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  awAck = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  wAck = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  wen = _RAND_2[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module AXI4PLIC(
  input         clock,
  input         reset,
  output        io__in_aw_ready, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input         io__in_aw_valid, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input  [31:0] io__in_aw_bits_addr, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output        io__in_w_ready, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input         io__in_w_valid, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input  [63:0] io__in_w_bits_data, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input  [7:0]  io__in_w_bits_strb, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input         io__in_b_ready, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output        io__in_b_valid, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output        io__in_ar_ready, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input         io__in_ar_valid, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input  [31:0] io__in_ar_bits_addr, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input         io__in_r_ready, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output        io__in_r_valid, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output [63:0] io__in_r_bits_data, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input         io__extra_intrVec, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output        io__extra_meip_0, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output        io_extra_meip_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
`endif // RANDOMIZE_REG_INIT
  wire  _r_busy_T = io__in_ar_ready & io__in_ar_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  wire  _r_busy_T_1 = io__in_r_ready & io__in_r_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  reg  r_busy; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  _GEN_0 = _r_busy_T_1 ? 1'h0 : r_busy; // @[src/main/scala/utils/StopWatch.scala 26:19 24:20 26:23]
  wire  _GEN_1 = _r_busy_T | _GEN_0; // @[src/main/scala/utils/StopWatch.scala 27:{20,24}]
  reg  ren_REG; // @[src/main/scala/device/AXI4Slave.scala 73:17]
  wire  _io_in_r_valid_T_2 = ren_REG & (_r_busy_T | r_busy); // @[src/main/scala/device/AXI4Slave.scala 74:35]
  reg  io_in_r_valid_r; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  _GEN_2 = _r_busy_T_1 ? 1'h0 : io_in_r_valid_r; // @[src/main/scala/utils/StopWatch.scala 26:19 24:20 26:23]
  wire  _GEN_3 = _io_in_r_valid_T_2 | _GEN_2; // @[src/main/scala/utils/StopWatch.scala 27:{20,24}]
  wire  _w_busy_T = io__in_aw_ready & io__in_aw_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  wire  _w_busy_T_1 = io__in_b_ready & io__in_b_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  reg  w_busy; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  _GEN_4 = _w_busy_T_1 ? 1'h0 : w_busy; // @[src/main/scala/utils/StopWatch.scala 26:19 24:20 26:23]
  wire  _GEN_5 = _w_busy_T | _GEN_4; // @[src/main/scala/utils/StopWatch.scala 27:{20,24}]
  wire  _io_in_b_valid_T = io__in_w_ready & io__in_w_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  reg  io_in_b_valid_r; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  _GEN_6 = _w_busy_T_1 ? 1'h0 : io_in_b_valid_r; // @[src/main/scala/utils/StopWatch.scala 26:19 24:20 26:23]
  wire  _GEN_7 = _io_in_b_valid_T | _GEN_6; // @[src/main/scala/utils/StopWatch.scala 27:{20,24}]
  reg [31:0] priority_0; // @[src/main/scala/device/AXI4PLIC.scala 37:39]
  reg  pending_0_1; // @[src/main/scala/device/AXI4PLIC.scala 43:46]
  wire [31:0] _T = {16'h0,8'h0,4'h0,2'h0,pending_0_1,1'h0}; // @[src/main/scala/device/AXI4PLIC.scala 45:38]
  reg [31:0] enable_0_0; // @[src/main/scala/device/AXI4PLIC.scala 48:64]
  reg [31:0] threshold_0; // @[src/main/scala/device/AXI4PLIC.scala 53:40]
  reg  inHandle_1; // @[src/main/scala/device/AXI4PLIC.scala 58:25]
  reg [31:0] claimCompletion_0; // @[src/main/scala/device/AXI4PLIC.scala 64:46]
  wire  _GEN_11 = _r_busy_T_1 & io__in_ar_bits_addr[25:0] == 26'h200004 ? claimCompletion_0[0] | inHandle_1 : inHandle_1
    ; // @[src/main/scala/device/AXI4PLIC.scala 58:25 68:57]
  wire  _GEN_12 = io__extra_intrVec | pending_0_1; // @[src/main/scala/device/AXI4PLIC.scala 75:{17,45} 43:46]
  wire [31:0] takenVec = _T & enable_0_0; // @[src/main/scala/device/AXI4PLIC.scala 81:31]
  wire [4:0] _claimCompletion_0_T_33 = takenVec[30] ? 5'h1e : 5'h1f; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [4:0] _claimCompletion_0_T_34 = takenVec[29] ? 5'h1d : _claimCompletion_0_T_33; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [4:0] _claimCompletion_0_T_35 = takenVec[28] ? 5'h1c : _claimCompletion_0_T_34; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [4:0] _claimCompletion_0_T_36 = takenVec[27] ? 5'h1b : _claimCompletion_0_T_35; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [4:0] _claimCompletion_0_T_37 = takenVec[26] ? 5'h1a : _claimCompletion_0_T_36; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [4:0] _claimCompletion_0_T_38 = takenVec[25] ? 5'h19 : _claimCompletion_0_T_37; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [4:0] _claimCompletion_0_T_39 = takenVec[24] ? 5'h18 : _claimCompletion_0_T_38; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [4:0] _claimCompletion_0_T_40 = takenVec[23] ? 5'h17 : _claimCompletion_0_T_39; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [4:0] _claimCompletion_0_T_41 = takenVec[22] ? 5'h16 : _claimCompletion_0_T_40; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [4:0] _claimCompletion_0_T_42 = takenVec[21] ? 5'h15 : _claimCompletion_0_T_41; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [4:0] _claimCompletion_0_T_43 = takenVec[20] ? 5'h14 : _claimCompletion_0_T_42; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [4:0] _claimCompletion_0_T_44 = takenVec[19] ? 5'h13 : _claimCompletion_0_T_43; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [4:0] _claimCompletion_0_T_45 = takenVec[18] ? 5'h12 : _claimCompletion_0_T_44; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [4:0] _claimCompletion_0_T_46 = takenVec[17] ? 5'h11 : _claimCompletion_0_T_45; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [4:0] _claimCompletion_0_T_47 = takenVec[16] ? 5'h10 : _claimCompletion_0_T_46; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [4:0] _claimCompletion_0_T_48 = takenVec[15] ? 5'hf : _claimCompletion_0_T_47; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [4:0] _claimCompletion_0_T_49 = takenVec[14] ? 5'he : _claimCompletion_0_T_48; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [4:0] _claimCompletion_0_T_50 = takenVec[13] ? 5'hd : _claimCompletion_0_T_49; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [4:0] _claimCompletion_0_T_51 = takenVec[12] ? 5'hc : _claimCompletion_0_T_50; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [4:0] _claimCompletion_0_T_52 = takenVec[11] ? 5'hb : _claimCompletion_0_T_51; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [4:0] _claimCompletion_0_T_53 = takenVec[10] ? 5'ha : _claimCompletion_0_T_52; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [4:0] _claimCompletion_0_T_54 = takenVec[9] ? 5'h9 : _claimCompletion_0_T_53; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [4:0] _claimCompletion_0_T_55 = takenVec[8] ? 5'h8 : _claimCompletion_0_T_54; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [4:0] _claimCompletion_0_T_56 = takenVec[7] ? 5'h7 : _claimCompletion_0_T_55; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [4:0] _claimCompletion_0_T_57 = takenVec[6] ? 5'h6 : _claimCompletion_0_T_56; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [4:0] _claimCompletion_0_T_58 = takenVec[5] ? 5'h5 : _claimCompletion_0_T_57; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [4:0] _claimCompletion_0_T_59 = takenVec[4] ? 5'h4 : _claimCompletion_0_T_58; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [4:0] _claimCompletion_0_T_60 = takenVec[3] ? 5'h3 : _claimCompletion_0_T_59; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [4:0] _claimCompletion_0_T_61 = takenVec[2] ? 5'h2 : _claimCompletion_0_T_60; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [4:0] _claimCompletion_0_T_62 = takenVec[1] ? 5'h1 : _claimCompletion_0_T_61; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [4:0] _claimCompletion_0_T_63 = takenVec[0] ? 5'h0 : _claimCompletion_0_T_62; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [4:0] _claimCompletion_0_T_64 = takenVec == 32'h0 ? 5'h0 : _claimCompletion_0_T_63; // @[src/main/scala/device/AXI4PLIC.scala 82:13]
  wire [7:0] _T_12 = io__in_w_bits_strb >> io__in_aw_bits_addr[2:0]; // @[src/main/scala/device/AXI4PLIC.scala 90:31]
  wire [7:0] _T_22 = _T_12[0] ? 8'hff : 8'h0; // @[src/main/scala/utils/BitUtils.scala 27:45]
  wire [7:0] _T_24 = _T_12[1] ? 8'hff : 8'h0; // @[src/main/scala/utils/BitUtils.scala 27:45]
  wire [7:0] _T_26 = _T_12[2] ? 8'hff : 8'h0; // @[src/main/scala/utils/BitUtils.scala 27:45]
  wire [7:0] _T_28 = _T_12[3] ? 8'hff : 8'h0; // @[src/main/scala/utils/BitUtils.scala 27:45]
  wire [7:0] _T_30 = _T_12[4] ? 8'hff : 8'h0; // @[src/main/scala/utils/BitUtils.scala 27:45]
  wire [7:0] _T_32 = _T_12[5] ? 8'hff : 8'h0; // @[src/main/scala/utils/BitUtils.scala 27:45]
  wire [7:0] _T_34 = _T_12[6] ? 8'hff : 8'h0; // @[src/main/scala/utils/BitUtils.scala 27:45]
  wire [7:0] _T_36 = _T_12[7] ? 8'hff : 8'h0; // @[src/main/scala/utils/BitUtils.scala 27:45]
  wire [63:0] _T_37 = {_T_36,_T_34,_T_32,_T_30,_T_28,_T_26,_T_24,_T_22}; // @[src/main/scala/utils/BitUtils.scala 27:26]
  wire  _rdata_T = 26'h1000 == io__in_ar_bits_addr[25:0]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _rdata_T_1 = 26'h2000 == io__in_ar_bits_addr[25:0]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _rdata_T_2 = 26'h200004 == io__in_ar_bits_addr[25:0]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _rdata_T_3 = 26'h4 == io__in_ar_bits_addr[25:0]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _rdata_T_4 = 26'h200000 == io__in_ar_bits_addr[25:0]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [31:0] _rdata_T_5 = _rdata_T ? _T : 32'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] _rdata_T_6 = _rdata_T_1 ? enable_0_0 : 32'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] _rdata_T_7 = _rdata_T_2 ? claimCompletion_0 : 32'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] _rdata_T_8 = _rdata_T_3 ? priority_0 : 32'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] _rdata_T_9 = _rdata_T_4 ? threshold_0 : 32'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] _rdata_T_10 = _rdata_T_5 | _rdata_T_6; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] _rdata_T_11 = _rdata_T_10 | _rdata_T_7; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] _rdata_T_12 = _rdata_T_11 | _rdata_T_8; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] rdata = _rdata_T_12 | _rdata_T_9; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] _enable_0_0_T = io__in_w_bits_data[31:0] & _T_37[31:0]; // @[src/main/scala/utils/BitUtils.scala 34:14]
  wire [31:0] _enable_0_0_T_1 = ~_T_37[31:0]; // @[src/main/scala/utils/BitUtils.scala 34:39]
  wire [31:0] _enable_0_0_T_2 = enable_0_0 & _enable_0_0_T_1; // @[src/main/scala/utils/BitUtils.scala 34:37]
  wire [31:0] _enable_0_0_T_3 = _enable_0_0_T | _enable_0_0_T_2; // @[src/main/scala/utils/BitUtils.scala 34:26]
  wire [31:0] _claimCompletion_0_T_67 = claimCompletion_0 & _enable_0_0_T_1; // @[src/main/scala/utils/BitUtils.scala 34:37]
  wire [31:0] _claimCompletion_0_T_68 = _enable_0_0_T | _claimCompletion_0_T_67; // @[src/main/scala/utils/BitUtils.scala 34:26]
  wire [4:0] _GEN_19 = _io_in_b_valid_T & io__in_aw_bits_addr[25:0] == 26'h200004 ? 5'h0 : _claimCompletion_0_T_64; // @[src/main/scala/utils/RegMap.scala 32:{48,52} src/main/scala/device/AXI4PLIC.scala 82:7]
  wire [31:0] _priority_0_T_2 = priority_0 & _enable_0_0_T_1; // @[src/main/scala/utils/BitUtils.scala 34:37]
  wire [31:0] _priority_0_T_3 = _enable_0_0_T | _priority_0_T_2; // @[src/main/scala/utils/BitUtils.scala 34:26]
  wire [31:0] _threshold_0_T_2 = threshold_0 & _enable_0_0_T_1; // @[src/main/scala/utils/BitUtils.scala 34:37]
  wire [31:0] _threshold_0_T_3 = _enable_0_0_T | _threshold_0_T_2; // @[src/main/scala/utils/BitUtils.scala 34:26]
  assign io__in_aw_ready = ~w_busy; // @[src/main/scala/device/AXI4Slave.scala 94:18]
  assign io__in_w_ready = io__in_aw_valid | w_busy; // @[src/main/scala/device/AXI4Slave.scala 95:30]
  assign io__in_b_valid = io_in_b_valid_r; // @[src/main/scala/device/AXI4Slave.scala 97:14]
  assign io__in_ar_ready = io__in_r_ready | ~r_busy; // @[src/main/scala/device/AXI4Slave.scala 71:29]
  assign io__in_r_valid = io_in_r_valid_r; // @[src/main/scala/device/AXI4Slave.scala 74:14]
  assign io__in_r_bits_data = {rdata,rdata}; // @[src/main/scala/device/AXI4PLIC.scala 93:25]
  assign io__extra_meip_0 = claimCompletion_0 != 32'h0; // @[src/main/scala/device/AXI4PLIC.scala 95:87]
  assign io_extra_meip_0 = io__extra_meip_0;
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      r_busy <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else begin
      r_busy <= _GEN_1;
    end
    if (reset) begin // @[src/main/scala/device/AXI4Slave.scala 73:17]
      ren_REG <= 1'h0; // @[src/main/scala/device/AXI4Slave.scala 73:17]
    end else begin
      ren_REG <= _r_busy_T; // @[src/main/scala/device/AXI4Slave.scala 73:17]
    end
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      io_in_r_valid_r <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else begin
      io_in_r_valid_r <= _GEN_3;
    end
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      w_busy <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else begin
      w_busy <= _GEN_5;
    end
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      io_in_b_valid_r <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else begin
      io_in_b_valid_r <= _GEN_7;
    end
    if (_io_in_b_valid_T & io__in_aw_bits_addr[25:0] == 26'h4) begin // @[src/main/scala/utils/RegMap.scala 32:48]
      priority_0 <= _priority_0_T_3; // @[src/main/scala/utils/RegMap.scala 32:52]
    end
    if (reset) begin // @[src/main/scala/device/AXI4PLIC.scala 43:46]
      pending_0_1 <= 1'h0; // @[src/main/scala/device/AXI4PLIC.scala 43:46]
    end else if (inHandle_1) begin // @[src/main/scala/device/AXI4PLIC.scala 76:25]
      pending_0_1 <= 1'h0; // @[src/main/scala/device/AXI4PLIC.scala 76:53]
    end else begin
      pending_0_1 <= _GEN_12;
    end
    if (reset) begin // @[src/main/scala/device/AXI4PLIC.scala 48:64]
      enable_0_0 <= 32'h0; // @[src/main/scala/device/AXI4PLIC.scala 48:64]
    end else if (_io_in_b_valid_T & io__in_aw_bits_addr[25:0] == 26'h2000) begin // @[src/main/scala/utils/RegMap.scala 32:48]
      enable_0_0 <= _enable_0_0_T_3; // @[src/main/scala/utils/RegMap.scala 32:52]
    end
    if (_io_in_b_valid_T & io__in_aw_bits_addr[25:0] == 26'h200000) begin // @[src/main/scala/utils/RegMap.scala 32:48]
      threshold_0 <= _threshold_0_T_3; // @[src/main/scala/utils/RegMap.scala 32:52]
    end
    if (reset) begin // @[src/main/scala/device/AXI4PLIC.scala 58:25]
      inHandle_1 <= 1'h0; // @[src/main/scala/device/AXI4PLIC.scala 58:25]
    end else if (_io_in_b_valid_T & io__in_aw_bits_addr[25:0] == 26'h200004) begin // @[src/main/scala/utils/RegMap.scala 32:48]
      if (_claimCompletion_0_T_68[0]) begin // @[src/main/scala/device/AXI4PLIC.scala 60:27]
        inHandle_1 <= 1'h0; // @[src/main/scala/device/AXI4PLIC.scala 60:27]
      end else begin
        inHandle_1 <= _GEN_11;
      end
    end else begin
      inHandle_1 <= _GEN_11;
    end
    claimCompletion_0 <= {{27'd0}, _GEN_19};
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  r_busy = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  ren_REG = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  io_in_r_valid_r = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  w_busy = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  io_in_b_valid_r = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  priority_0 = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  pending_0_1 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  enable_0_0 = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  threshold_0 = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  inHandle_1 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  claimCompletion_0 = _RAND_10[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module NutShell(
  input         clock,
  input         reset,
  input         io_mem_aw_ready, // @[src/main/scala/system/NutShell.scala 45:14]
  output        io_mem_aw_valid, // @[src/main/scala/system/NutShell.scala 45:14]
  output [31:0] io_mem_aw_bits_addr, // @[src/main/scala/system/NutShell.scala 45:14]
  output [7:0]  io_mem_aw_bits_len, // @[src/main/scala/system/NutShell.scala 45:14]
  output [2:0]  io_mem_aw_bits_size, // @[src/main/scala/system/NutShell.scala 45:14]
  output [1:0]  io_mem_aw_bits_burst, // @[src/main/scala/system/NutShell.scala 45:14]
  input         io_mem_w_ready, // @[src/main/scala/system/NutShell.scala 45:14]
  output        io_mem_w_valid, // @[src/main/scala/system/NutShell.scala 45:14]
  output [63:0] io_mem_w_bits_data, // @[src/main/scala/system/NutShell.scala 45:14]
  output        io_mem_w_bits_last, // @[src/main/scala/system/NutShell.scala 45:14]
  input         io_mem_b_valid, // @[src/main/scala/system/NutShell.scala 45:14]
  input         io_mem_ar_ready, // @[src/main/scala/system/NutShell.scala 45:14]
  output        io_mem_ar_valid, // @[src/main/scala/system/NutShell.scala 45:14]
  output [31:0] io_mem_ar_bits_addr, // @[src/main/scala/system/NutShell.scala 45:14]
  output [7:0]  io_mem_ar_bits_len, // @[src/main/scala/system/NutShell.scala 45:14]
  input         io_mem_r_valid, // @[src/main/scala/system/NutShell.scala 45:14]
  input  [63:0] io_mem_r_bits_data, // @[src/main/scala/system/NutShell.scala 45:14]
  input         io_mem_r_bits_last, // @[src/main/scala/system/NutShell.scala 45:14]
  input         io_mmio_req_ready, // @[src/main/scala/system/NutShell.scala 45:14]
  output        io_mmio_req_valid, // @[src/main/scala/system/NutShell.scala 45:14]
  output [31:0] io_mmio_req_bits_addr, // @[src/main/scala/system/NutShell.scala 45:14]
  output [2:0]  io_mmio_req_bits_size, // @[src/main/scala/system/NutShell.scala 45:14]
  output [3:0]  io_mmio_req_bits_cmd, // @[src/main/scala/system/NutShell.scala 45:14]
  output [7:0]  io_mmio_req_bits_wmask, // @[src/main/scala/system/NutShell.scala 45:14]
  output [63:0] io_mmio_req_bits_wdata, // @[src/main/scala/system/NutShell.scala 45:14]
  output        io_mmio_resp_ready, // @[src/main/scala/system/NutShell.scala 45:14]
  input         io_mmio_resp_valid, // @[src/main/scala/system/NutShell.scala 45:14]
  input  [3:0]  io_mmio_resp_bits_cmd, // @[src/main/scala/system/NutShell.scala 45:14]
  input  [63:0] io_mmio_resp_bits_rdata, // @[src/main/scala/system/NutShell.scala 45:14]
  output        io_frontend_aw_ready, // @[src/main/scala/system/NutShell.scala 45:14]
  input         io_frontend_aw_valid, // @[src/main/scala/system/NutShell.scala 45:14]
  input  [31:0] io_frontend_aw_bits_addr, // @[src/main/scala/system/NutShell.scala 45:14]
  input  [7:0]  io_frontend_aw_bits_len, // @[src/main/scala/system/NutShell.scala 45:14]
  input  [2:0]  io_frontend_aw_bits_size, // @[src/main/scala/system/NutShell.scala 45:14]
  output        io_frontend_w_ready, // @[src/main/scala/system/NutShell.scala 45:14]
  input         io_frontend_w_valid, // @[src/main/scala/system/NutShell.scala 45:14]
  input  [63:0] io_frontend_w_bits_data, // @[src/main/scala/system/NutShell.scala 45:14]
  input  [7:0]  io_frontend_w_bits_strb, // @[src/main/scala/system/NutShell.scala 45:14]
  input         io_frontend_b_ready, // @[src/main/scala/system/NutShell.scala 45:14]
  output        io_frontend_b_valid, // @[src/main/scala/system/NutShell.scala 45:14]
  output        io_frontend_ar_ready, // @[src/main/scala/system/NutShell.scala 45:14]
  input         io_frontend_ar_valid, // @[src/main/scala/system/NutShell.scala 45:14]
  input  [31:0] io_frontend_ar_bits_addr, // @[src/main/scala/system/NutShell.scala 45:14]
  input         io_frontend_r_ready, // @[src/main/scala/system/NutShell.scala 45:14]
  output        io_frontend_r_valid, // @[src/main/scala/system/NutShell.scala 45:14]
  output [63:0] io_frontend_r_bits_data, // @[src/main/scala/system/NutShell.scala 45:14]
  input         io_meip, // @[src/main/scala/system/NutShell.scala 45:14]
  input         _WIRE_4
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  wire  nutcore_clock; // @[src/main/scala/system/NutShell.scala 53:23]
  wire  nutcore_reset; // @[src/main/scala/system/NutShell.scala 53:23]
  wire  nutcore_io_imem_mem_req_ready; // @[src/main/scala/system/NutShell.scala 53:23]
  wire  nutcore_io_imem_mem_req_valid; // @[src/main/scala/system/NutShell.scala 53:23]
  wire [31:0] nutcore_io_imem_mem_req_bits_addr; // @[src/main/scala/system/NutShell.scala 53:23]
  wire [3:0] nutcore_io_imem_mem_req_bits_cmd; // @[src/main/scala/system/NutShell.scala 53:23]
  wire [63:0] nutcore_io_imem_mem_req_bits_wdata; // @[src/main/scala/system/NutShell.scala 53:23]
  wire  nutcore_io_imem_mem_resp_valid; // @[src/main/scala/system/NutShell.scala 53:23]
  wire [3:0] nutcore_io_imem_mem_resp_bits_cmd; // @[src/main/scala/system/NutShell.scala 53:23]
  wire [63:0] nutcore_io_imem_mem_resp_bits_rdata; // @[src/main/scala/system/NutShell.scala 53:23]
  wire  nutcore_io_dmem_mem_req_ready; // @[src/main/scala/system/NutShell.scala 53:23]
  wire  nutcore_io_dmem_mem_req_valid; // @[src/main/scala/system/NutShell.scala 53:23]
  wire [31:0] nutcore_io_dmem_mem_req_bits_addr; // @[src/main/scala/system/NutShell.scala 53:23]
  wire [3:0] nutcore_io_dmem_mem_req_bits_cmd; // @[src/main/scala/system/NutShell.scala 53:23]
  wire [63:0] nutcore_io_dmem_mem_req_bits_wdata; // @[src/main/scala/system/NutShell.scala 53:23]
  wire  nutcore_io_dmem_mem_resp_valid; // @[src/main/scala/system/NutShell.scala 53:23]
  wire [3:0] nutcore_io_dmem_mem_resp_bits_cmd; // @[src/main/scala/system/NutShell.scala 53:23]
  wire [63:0] nutcore_io_dmem_mem_resp_bits_rdata; // @[src/main/scala/system/NutShell.scala 53:23]
  wire  nutcore_io_dmem_coh_req_ready; // @[src/main/scala/system/NutShell.scala 53:23]
  wire  nutcore_io_dmem_coh_req_valid; // @[src/main/scala/system/NutShell.scala 53:23]
  wire [31:0] nutcore_io_dmem_coh_req_bits_addr; // @[src/main/scala/system/NutShell.scala 53:23]
  wire [63:0] nutcore_io_dmem_coh_req_bits_wdata; // @[src/main/scala/system/NutShell.scala 53:23]
  wire  nutcore_io_dmem_coh_resp_valid; // @[src/main/scala/system/NutShell.scala 53:23]
  wire [3:0] nutcore_io_dmem_coh_resp_bits_cmd; // @[src/main/scala/system/NutShell.scala 53:23]
  wire [63:0] nutcore_io_dmem_coh_resp_bits_rdata; // @[src/main/scala/system/NutShell.scala 53:23]
  wire  nutcore_io_mmio_req_ready; // @[src/main/scala/system/NutShell.scala 53:23]
  wire  nutcore_io_mmio_req_valid; // @[src/main/scala/system/NutShell.scala 53:23]
  wire [31:0] nutcore_io_mmio_req_bits_addr; // @[src/main/scala/system/NutShell.scala 53:23]
  wire [2:0] nutcore_io_mmio_req_bits_size; // @[src/main/scala/system/NutShell.scala 53:23]
  wire [3:0] nutcore_io_mmio_req_bits_cmd; // @[src/main/scala/system/NutShell.scala 53:23]
  wire [7:0] nutcore_io_mmio_req_bits_wmask; // @[src/main/scala/system/NutShell.scala 53:23]
  wire [63:0] nutcore_io_mmio_req_bits_wdata; // @[src/main/scala/system/NutShell.scala 53:23]
  wire  nutcore_io_mmio_resp_valid; // @[src/main/scala/system/NutShell.scala 53:23]
  wire [3:0] nutcore_io_mmio_resp_bits_cmd; // @[src/main/scala/system/NutShell.scala 53:23]
  wire [63:0] nutcore_io_mmio_resp_bits_rdata; // @[src/main/scala/system/NutShell.scala 53:23]
  wire  nutcore_io_frontend_req_ready; // @[src/main/scala/system/NutShell.scala 53:23]
  wire  nutcore_io_frontend_req_valid; // @[src/main/scala/system/NutShell.scala 53:23]
  wire [31:0] nutcore_io_frontend_req_bits_addr; // @[src/main/scala/system/NutShell.scala 53:23]
  wire [2:0] nutcore_io_frontend_req_bits_size; // @[src/main/scala/system/NutShell.scala 53:23]
  wire [3:0] nutcore_io_frontend_req_bits_cmd; // @[src/main/scala/system/NutShell.scala 53:23]
  wire [7:0] nutcore_io_frontend_req_bits_wmask; // @[src/main/scala/system/NutShell.scala 53:23]
  wire [63:0] nutcore_io_frontend_req_bits_wdata; // @[src/main/scala/system/NutShell.scala 53:23]
  wire  nutcore_io_frontend_resp_ready; // @[src/main/scala/system/NutShell.scala 53:23]
  wire  nutcore_io_frontend_resp_valid; // @[src/main/scala/system/NutShell.scala 53:23]
  wire [3:0] nutcore_io_frontend_resp_bits_cmd; // @[src/main/scala/system/NutShell.scala 53:23]
  wire [63:0] nutcore_io_frontend_resp_bits_rdata; // @[src/main/scala/system/NutShell.scala 53:23]
  wire  nutcore_io_extra_meip_0; // @[src/main/scala/system/NutShell.scala 53:23]
  wire  nutcore__WIRE_0; // @[src/main/scala/system/NutShell.scala 53:23]
  wire  nutcore_DISPLAY_ENABLE; // @[src/main/scala/system/NutShell.scala 53:23]
  wire  nutcore_io_extra_mtip; // @[src/main/scala/system/NutShell.scala 53:23]
  wire  nutcore_io_extra_msip; // @[src/main/scala/system/NutShell.scala 53:23]
  wire  cohMg_clock; // @[src/main/scala/system/NutShell.scala 54:21]
  wire  cohMg_reset; // @[src/main/scala/system/NutShell.scala 54:21]
  wire  cohMg_io_in_req_ready; // @[src/main/scala/system/NutShell.scala 54:21]
  wire  cohMg_io_in_req_valid; // @[src/main/scala/system/NutShell.scala 54:21]
  wire [31:0] cohMg_io_in_req_bits_addr; // @[src/main/scala/system/NutShell.scala 54:21]
  wire [3:0] cohMg_io_in_req_bits_cmd; // @[src/main/scala/system/NutShell.scala 54:21]
  wire [63:0] cohMg_io_in_req_bits_wdata; // @[src/main/scala/system/NutShell.scala 54:21]
  wire  cohMg_io_in_resp_valid; // @[src/main/scala/system/NutShell.scala 54:21]
  wire [3:0] cohMg_io_in_resp_bits_cmd; // @[src/main/scala/system/NutShell.scala 54:21]
  wire [63:0] cohMg_io_in_resp_bits_rdata; // @[src/main/scala/system/NutShell.scala 54:21]
  wire  cohMg_io_out_mem_req_ready; // @[src/main/scala/system/NutShell.scala 54:21]
  wire  cohMg_io_out_mem_req_valid; // @[src/main/scala/system/NutShell.scala 54:21]
  wire [31:0] cohMg_io_out_mem_req_bits_addr; // @[src/main/scala/system/NutShell.scala 54:21]
  wire [3:0] cohMg_io_out_mem_req_bits_cmd; // @[src/main/scala/system/NutShell.scala 54:21]
  wire [63:0] cohMg_io_out_mem_req_bits_wdata; // @[src/main/scala/system/NutShell.scala 54:21]
  wire  cohMg_io_out_mem_resp_ready; // @[src/main/scala/system/NutShell.scala 54:21]
  wire  cohMg_io_out_mem_resp_valid; // @[src/main/scala/system/NutShell.scala 54:21]
  wire [3:0] cohMg_io_out_mem_resp_bits_cmd; // @[src/main/scala/system/NutShell.scala 54:21]
  wire [63:0] cohMg_io_out_mem_resp_bits_rdata; // @[src/main/scala/system/NutShell.scala 54:21]
  wire  cohMg_io_out_coh_req_ready; // @[src/main/scala/system/NutShell.scala 54:21]
  wire  cohMg_io_out_coh_req_valid; // @[src/main/scala/system/NutShell.scala 54:21]
  wire [31:0] cohMg_io_out_coh_req_bits_addr; // @[src/main/scala/system/NutShell.scala 54:21]
  wire [63:0] cohMg_io_out_coh_req_bits_wdata; // @[src/main/scala/system/NutShell.scala 54:21]
  wire  cohMg_io_out_coh_resp_ready; // @[src/main/scala/system/NutShell.scala 54:21]
  wire  cohMg_io_out_coh_resp_valid; // @[src/main/scala/system/NutShell.scala 54:21]
  wire [3:0] cohMg_io_out_coh_resp_bits_cmd; // @[src/main/scala/system/NutShell.scala 54:21]
  wire [63:0] cohMg_io_out_coh_resp_bits_rdata; // @[src/main/scala/system/NutShell.scala 54:21]
  wire  xbar_clock; // @[src/main/scala/system/NutShell.scala 55:20]
  wire  xbar_reset; // @[src/main/scala/system/NutShell.scala 55:20]
  wire  xbar_io_in_0_req_ready; // @[src/main/scala/system/NutShell.scala 55:20]
  wire  xbar_io_in_0_req_valid; // @[src/main/scala/system/NutShell.scala 55:20]
  wire [31:0] xbar_io_in_0_req_bits_addr; // @[src/main/scala/system/NutShell.scala 55:20]
  wire [3:0] xbar_io_in_0_req_bits_cmd; // @[src/main/scala/system/NutShell.scala 55:20]
  wire [7:0] xbar_io_in_0_req_bits_wmask; // @[src/main/scala/system/NutShell.scala 55:20]
  wire [63:0] xbar_io_in_0_req_bits_wdata; // @[src/main/scala/system/NutShell.scala 55:20]
  wire  xbar_io_in_0_resp_valid; // @[src/main/scala/system/NutShell.scala 55:20]
  wire [3:0] xbar_io_in_0_resp_bits_cmd; // @[src/main/scala/system/NutShell.scala 55:20]
  wire [63:0] xbar_io_in_0_resp_bits_rdata; // @[src/main/scala/system/NutShell.scala 55:20]
  wire  xbar_io_in_1_req_ready; // @[src/main/scala/system/NutShell.scala 55:20]
  wire  xbar_io_in_1_req_valid; // @[src/main/scala/system/NutShell.scala 55:20]
  wire [31:0] xbar_io_in_1_req_bits_addr; // @[src/main/scala/system/NutShell.scala 55:20]
  wire [2:0] xbar_io_in_1_req_bits_size; // @[src/main/scala/system/NutShell.scala 55:20]
  wire [3:0] xbar_io_in_1_req_bits_cmd; // @[src/main/scala/system/NutShell.scala 55:20]
  wire [7:0] xbar_io_in_1_req_bits_wmask; // @[src/main/scala/system/NutShell.scala 55:20]
  wire [63:0] xbar_io_in_1_req_bits_wdata; // @[src/main/scala/system/NutShell.scala 55:20]
  wire  xbar_io_in_1_resp_valid; // @[src/main/scala/system/NutShell.scala 55:20]
  wire [3:0] xbar_io_in_1_resp_bits_cmd; // @[src/main/scala/system/NutShell.scala 55:20]
  wire [63:0] xbar_io_in_1_resp_bits_rdata; // @[src/main/scala/system/NutShell.scala 55:20]
  wire  xbar_io_out_req_ready; // @[src/main/scala/system/NutShell.scala 55:20]
  wire  xbar_io_out_req_valid; // @[src/main/scala/system/NutShell.scala 55:20]
  wire [31:0] xbar_io_out_req_bits_addr; // @[src/main/scala/system/NutShell.scala 55:20]
  wire [2:0] xbar_io_out_req_bits_size; // @[src/main/scala/system/NutShell.scala 55:20]
  wire [3:0] xbar_io_out_req_bits_cmd; // @[src/main/scala/system/NutShell.scala 55:20]
  wire [7:0] xbar_io_out_req_bits_wmask; // @[src/main/scala/system/NutShell.scala 55:20]
  wire [63:0] xbar_io_out_req_bits_wdata; // @[src/main/scala/system/NutShell.scala 55:20]
  wire  xbar_io_out_resp_ready; // @[src/main/scala/system/NutShell.scala 55:20]
  wire  xbar_io_out_resp_valid; // @[src/main/scala/system/NutShell.scala 55:20]
  wire [3:0] xbar_io_out_resp_bits_cmd; // @[src/main/scala/system/NutShell.scala 55:20]
  wire [63:0] xbar_io_out_resp_bits_rdata; // @[src/main/scala/system/NutShell.scala 55:20]
  wire  axi2sb_clock; // @[src/main/scala/system/NutShell.scala 61:22]
  wire  axi2sb_reset; // @[src/main/scala/system/NutShell.scala 61:22]
  wire  axi2sb_io_in_aw_ready; // @[src/main/scala/system/NutShell.scala 61:22]
  wire  axi2sb_io_in_aw_valid; // @[src/main/scala/system/NutShell.scala 61:22]
  wire [31:0] axi2sb_io_in_aw_bits_addr; // @[src/main/scala/system/NutShell.scala 61:22]
  wire [7:0] axi2sb_io_in_aw_bits_len; // @[src/main/scala/system/NutShell.scala 61:22]
  wire [2:0] axi2sb_io_in_aw_bits_size; // @[src/main/scala/system/NutShell.scala 61:22]
  wire  axi2sb_io_in_w_ready; // @[src/main/scala/system/NutShell.scala 61:22]
  wire  axi2sb_io_in_w_valid; // @[src/main/scala/system/NutShell.scala 61:22]
  wire [63:0] axi2sb_io_in_w_bits_data; // @[src/main/scala/system/NutShell.scala 61:22]
  wire [7:0] axi2sb_io_in_w_bits_strb; // @[src/main/scala/system/NutShell.scala 61:22]
  wire  axi2sb_io_in_b_ready; // @[src/main/scala/system/NutShell.scala 61:22]
  wire  axi2sb_io_in_b_valid; // @[src/main/scala/system/NutShell.scala 61:22]
  wire  axi2sb_io_in_ar_ready; // @[src/main/scala/system/NutShell.scala 61:22]
  wire  axi2sb_io_in_ar_valid; // @[src/main/scala/system/NutShell.scala 61:22]
  wire [31:0] axi2sb_io_in_ar_bits_addr; // @[src/main/scala/system/NutShell.scala 61:22]
  wire  axi2sb_io_in_r_ready; // @[src/main/scala/system/NutShell.scala 61:22]
  wire  axi2sb_io_in_r_valid; // @[src/main/scala/system/NutShell.scala 61:22]
  wire [63:0] axi2sb_io_in_r_bits_data; // @[src/main/scala/system/NutShell.scala 61:22]
  wire  axi2sb_io_out_req_ready; // @[src/main/scala/system/NutShell.scala 61:22]
  wire  axi2sb_io_out_req_valid; // @[src/main/scala/system/NutShell.scala 61:22]
  wire [31:0] axi2sb_io_out_req_bits_addr; // @[src/main/scala/system/NutShell.scala 61:22]
  wire [2:0] axi2sb_io_out_req_bits_size; // @[src/main/scala/system/NutShell.scala 61:22]
  wire [3:0] axi2sb_io_out_req_bits_cmd; // @[src/main/scala/system/NutShell.scala 61:22]
  wire [7:0] axi2sb_io_out_req_bits_wmask; // @[src/main/scala/system/NutShell.scala 61:22]
  wire [63:0] axi2sb_io_out_req_bits_wdata; // @[src/main/scala/system/NutShell.scala 61:22]
  wire  axi2sb_io_out_resp_ready; // @[src/main/scala/system/NutShell.scala 61:22]
  wire  axi2sb_io_out_resp_valid; // @[src/main/scala/system/NutShell.scala 61:22]
  wire [3:0] axi2sb_io_out_resp_bits_cmd; // @[src/main/scala/system/NutShell.scala 61:22]
  wire [63:0] axi2sb_io_out_resp_bits_rdata; // @[src/main/scala/system/NutShell.scala 61:22]
  wire  mem_l2cacheIn_prefetcher_clock; // @[src/main/scala/system/NutShell.scala 73:30]
  wire  mem_l2cacheIn_prefetcher_reset; // @[src/main/scala/system/NutShell.scala 73:30]
  wire  mem_l2cacheIn_prefetcher_io_in_ready; // @[src/main/scala/system/NutShell.scala 73:30]
  wire  mem_l2cacheIn_prefetcher_io_in_valid; // @[src/main/scala/system/NutShell.scala 73:30]
  wire [31:0] mem_l2cacheIn_prefetcher_io_in_bits_addr; // @[src/main/scala/system/NutShell.scala 73:30]
  wire [2:0] mem_l2cacheIn_prefetcher_io_in_bits_size; // @[src/main/scala/system/NutShell.scala 73:30]
  wire [3:0] mem_l2cacheIn_prefetcher_io_in_bits_cmd; // @[src/main/scala/system/NutShell.scala 73:30]
  wire [7:0] mem_l2cacheIn_prefetcher_io_in_bits_wmask; // @[src/main/scala/system/NutShell.scala 73:30]
  wire [63:0] mem_l2cacheIn_prefetcher_io_in_bits_wdata; // @[src/main/scala/system/NutShell.scala 73:30]
  wire  mem_l2cacheIn_prefetcher_io_out_ready; // @[src/main/scala/system/NutShell.scala 73:30]
  wire  mem_l2cacheIn_prefetcher_io_out_valid; // @[src/main/scala/system/NutShell.scala 73:30]
  wire [31:0] mem_l2cacheIn_prefetcher_io_out_bits_addr; // @[src/main/scala/system/NutShell.scala 73:30]
  wire [2:0] mem_l2cacheIn_prefetcher_io_out_bits_size; // @[src/main/scala/system/NutShell.scala 73:30]
  wire [3:0] mem_l2cacheIn_prefetcher_io_out_bits_cmd; // @[src/main/scala/system/NutShell.scala 73:30]
  wire [7:0] mem_l2cacheIn_prefetcher_io_out_bits_wmask; // @[src/main/scala/system/NutShell.scala 73:30]
  wire [63:0] mem_l2cacheIn_prefetcher_io_out_bits_wdata; // @[src/main/scala/system/NutShell.scala 73:30]
  wire  mem_l2cacheIn_prefetcher_DISPLAY_ENABLE; // @[src/main/scala/system/NutShell.scala 73:30]
  wire  mem_l2cacheOut_cache_clock; // @[src/main/scala/nutcore/mem/Cache.scala 668:35]
  wire  mem_l2cacheOut_cache_reset; // @[src/main/scala/nutcore/mem/Cache.scala 668:35]
  wire  mem_l2cacheOut_cache_io_in_req_ready; // @[src/main/scala/nutcore/mem/Cache.scala 668:35]
  wire  mem_l2cacheOut_cache_io_in_req_valid; // @[src/main/scala/nutcore/mem/Cache.scala 668:35]
  wire [31:0] mem_l2cacheOut_cache_io_in_req_bits_addr; // @[src/main/scala/nutcore/mem/Cache.scala 668:35]
  wire [2:0] mem_l2cacheOut_cache_io_in_req_bits_size; // @[src/main/scala/nutcore/mem/Cache.scala 668:35]
  wire [3:0] mem_l2cacheOut_cache_io_in_req_bits_cmd; // @[src/main/scala/nutcore/mem/Cache.scala 668:35]
  wire [7:0] mem_l2cacheOut_cache_io_in_req_bits_wmask; // @[src/main/scala/nutcore/mem/Cache.scala 668:35]
  wire [63:0] mem_l2cacheOut_cache_io_in_req_bits_wdata; // @[src/main/scala/nutcore/mem/Cache.scala 668:35]
  wire  mem_l2cacheOut_cache_io_in_resp_valid; // @[src/main/scala/nutcore/mem/Cache.scala 668:35]
  wire [3:0] mem_l2cacheOut_cache_io_in_resp_bits_cmd; // @[src/main/scala/nutcore/mem/Cache.scala 668:35]
  wire [63:0] mem_l2cacheOut_cache_io_in_resp_bits_rdata; // @[src/main/scala/nutcore/mem/Cache.scala 668:35]
  wire  mem_l2cacheOut_cache_io_out_mem_req_ready; // @[src/main/scala/nutcore/mem/Cache.scala 668:35]
  wire  mem_l2cacheOut_cache_io_out_mem_req_valid; // @[src/main/scala/nutcore/mem/Cache.scala 668:35]
  wire [31:0] mem_l2cacheOut_cache_io_out_mem_req_bits_addr; // @[src/main/scala/nutcore/mem/Cache.scala 668:35]
  wire [3:0] mem_l2cacheOut_cache_io_out_mem_req_bits_cmd; // @[src/main/scala/nutcore/mem/Cache.scala 668:35]
  wire [63:0] mem_l2cacheOut_cache_io_out_mem_req_bits_wdata; // @[src/main/scala/nutcore/mem/Cache.scala 668:35]
  wire  mem_l2cacheOut_cache_io_out_mem_resp_valid; // @[src/main/scala/nutcore/mem/Cache.scala 668:35]
  wire [3:0] mem_l2cacheOut_cache_io_out_mem_resp_bits_cmd; // @[src/main/scala/nutcore/mem/Cache.scala 668:35]
  wire [63:0] mem_l2cacheOut_cache_io_out_mem_resp_bits_rdata; // @[src/main/scala/nutcore/mem/Cache.scala 668:35]
  wire  mem_l2cacheOut_cache_DISPLAY_ENABLE; // @[src/main/scala/nutcore/mem/Cache.scala 668:35]
  wire  memAddrMap_io_in_req_ready; // @[src/main/scala/system/NutShell.scala 93:26]
  wire  memAddrMap_io_in_req_valid; // @[src/main/scala/system/NutShell.scala 93:26]
  wire [31:0] memAddrMap_io_in_req_bits_addr; // @[src/main/scala/system/NutShell.scala 93:26]
  wire [3:0] memAddrMap_io_in_req_bits_cmd; // @[src/main/scala/system/NutShell.scala 93:26]
  wire [63:0] memAddrMap_io_in_req_bits_wdata; // @[src/main/scala/system/NutShell.scala 93:26]
  wire  memAddrMap_io_in_resp_valid; // @[src/main/scala/system/NutShell.scala 93:26]
  wire [3:0] memAddrMap_io_in_resp_bits_cmd; // @[src/main/scala/system/NutShell.scala 93:26]
  wire [63:0] memAddrMap_io_in_resp_bits_rdata; // @[src/main/scala/system/NutShell.scala 93:26]
  wire  memAddrMap_io_out_req_ready; // @[src/main/scala/system/NutShell.scala 93:26]
  wire  memAddrMap_io_out_req_valid; // @[src/main/scala/system/NutShell.scala 93:26]
  wire [31:0] memAddrMap_io_out_req_bits_addr; // @[src/main/scala/system/NutShell.scala 93:26]
  wire [3:0] memAddrMap_io_out_req_bits_cmd; // @[src/main/scala/system/NutShell.scala 93:26]
  wire [63:0] memAddrMap_io_out_req_bits_wdata; // @[src/main/scala/system/NutShell.scala 93:26]
  wire  memAddrMap_io_out_resp_valid; // @[src/main/scala/system/NutShell.scala 93:26]
  wire [3:0] memAddrMap_io_out_resp_bits_cmd; // @[src/main/scala/system/NutShell.scala 93:26]
  wire [63:0] memAddrMap_io_out_resp_bits_rdata; // @[src/main/scala/system/NutShell.scala 93:26]
  wire  io_mem_bridge_clock; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  io_mem_bridge_reset; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  io_mem_bridge_io_in_req_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  io_mem_bridge_io_in_req_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [31:0] io_mem_bridge_io_in_req_bits_addr; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [3:0] io_mem_bridge_io_in_req_bits_cmd; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [63:0] io_mem_bridge_io_in_req_bits_wdata; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  io_mem_bridge_io_in_resp_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [3:0] io_mem_bridge_io_in_resp_bits_cmd; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [63:0] io_mem_bridge_io_in_resp_bits_rdata; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  io_mem_bridge_io_out_aw_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  io_mem_bridge_io_out_aw_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [31:0] io_mem_bridge_io_out_aw_bits_addr; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [7:0] io_mem_bridge_io_out_aw_bits_len; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [2:0] io_mem_bridge_io_out_aw_bits_size; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [1:0] io_mem_bridge_io_out_aw_bits_burst; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  io_mem_bridge_io_out_w_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  io_mem_bridge_io_out_w_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [63:0] io_mem_bridge_io_out_w_bits_data; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  io_mem_bridge_io_out_w_bits_last; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  io_mem_bridge_io_out_b_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  io_mem_bridge_io_out_ar_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  io_mem_bridge_io_out_ar_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [31:0] io_mem_bridge_io_out_ar_bits_addr; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [7:0] io_mem_bridge_io_out_ar_bits_len; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [2:0] io_mem_bridge_io_out_ar_bits_size; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [1:0] io_mem_bridge_io_out_ar_bits_burst; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  io_mem_bridge_io_out_r_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [63:0] io_mem_bridge_io_out_r_bits_data; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  io_mem_bridge_io_out_r_bits_last; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  mmioXbar_clock; // @[src/main/scala/system/NutShell.scala 106:24]
  wire  mmioXbar_reset; // @[src/main/scala/system/NutShell.scala 106:24]
  wire  mmioXbar_io_in_req_ready; // @[src/main/scala/system/NutShell.scala 106:24]
  wire  mmioXbar_io_in_req_valid; // @[src/main/scala/system/NutShell.scala 106:24]
  wire [31:0] mmioXbar_io_in_req_bits_addr; // @[src/main/scala/system/NutShell.scala 106:24]
  wire [2:0] mmioXbar_io_in_req_bits_size; // @[src/main/scala/system/NutShell.scala 106:24]
  wire [3:0] mmioXbar_io_in_req_bits_cmd; // @[src/main/scala/system/NutShell.scala 106:24]
  wire [7:0] mmioXbar_io_in_req_bits_wmask; // @[src/main/scala/system/NutShell.scala 106:24]
  wire [63:0] mmioXbar_io_in_req_bits_wdata; // @[src/main/scala/system/NutShell.scala 106:24]
  wire  mmioXbar_io_in_resp_valid; // @[src/main/scala/system/NutShell.scala 106:24]
  wire [3:0] mmioXbar_io_in_resp_bits_cmd; // @[src/main/scala/system/NutShell.scala 106:24]
  wire [63:0] mmioXbar_io_in_resp_bits_rdata; // @[src/main/scala/system/NutShell.scala 106:24]
  wire  mmioXbar_io_out_0_req_ready; // @[src/main/scala/system/NutShell.scala 106:24]
  wire  mmioXbar_io_out_0_req_valid; // @[src/main/scala/system/NutShell.scala 106:24]
  wire [31:0] mmioXbar_io_out_0_req_bits_addr; // @[src/main/scala/system/NutShell.scala 106:24]
  wire [3:0] mmioXbar_io_out_0_req_bits_cmd; // @[src/main/scala/system/NutShell.scala 106:24]
  wire [7:0] mmioXbar_io_out_0_req_bits_wmask; // @[src/main/scala/system/NutShell.scala 106:24]
  wire [63:0] mmioXbar_io_out_0_req_bits_wdata; // @[src/main/scala/system/NutShell.scala 106:24]
  wire  mmioXbar_io_out_0_resp_ready; // @[src/main/scala/system/NutShell.scala 106:24]
  wire  mmioXbar_io_out_0_resp_valid; // @[src/main/scala/system/NutShell.scala 106:24]
  wire [63:0] mmioXbar_io_out_0_resp_bits_rdata; // @[src/main/scala/system/NutShell.scala 106:24]
  wire  mmioXbar_io_out_1_req_ready; // @[src/main/scala/system/NutShell.scala 106:24]
  wire  mmioXbar_io_out_1_req_valid; // @[src/main/scala/system/NutShell.scala 106:24]
  wire [31:0] mmioXbar_io_out_1_req_bits_addr; // @[src/main/scala/system/NutShell.scala 106:24]
  wire [3:0] mmioXbar_io_out_1_req_bits_cmd; // @[src/main/scala/system/NutShell.scala 106:24]
  wire [7:0] mmioXbar_io_out_1_req_bits_wmask; // @[src/main/scala/system/NutShell.scala 106:24]
  wire [63:0] mmioXbar_io_out_1_req_bits_wdata; // @[src/main/scala/system/NutShell.scala 106:24]
  wire  mmioXbar_io_out_1_resp_ready; // @[src/main/scala/system/NutShell.scala 106:24]
  wire  mmioXbar_io_out_1_resp_valid; // @[src/main/scala/system/NutShell.scala 106:24]
  wire [63:0] mmioXbar_io_out_1_resp_bits_rdata; // @[src/main/scala/system/NutShell.scala 106:24]
  wire  mmioXbar_io_out_2_req_ready; // @[src/main/scala/system/NutShell.scala 106:24]
  wire  mmioXbar_io_out_2_req_valid; // @[src/main/scala/system/NutShell.scala 106:24]
  wire [31:0] mmioXbar_io_out_2_req_bits_addr; // @[src/main/scala/system/NutShell.scala 106:24]
  wire [2:0] mmioXbar_io_out_2_req_bits_size; // @[src/main/scala/system/NutShell.scala 106:24]
  wire [3:0] mmioXbar_io_out_2_req_bits_cmd; // @[src/main/scala/system/NutShell.scala 106:24]
  wire [7:0] mmioXbar_io_out_2_req_bits_wmask; // @[src/main/scala/system/NutShell.scala 106:24]
  wire [63:0] mmioXbar_io_out_2_req_bits_wdata; // @[src/main/scala/system/NutShell.scala 106:24]
  wire  mmioXbar_io_out_2_resp_ready; // @[src/main/scala/system/NutShell.scala 106:24]
  wire  mmioXbar_io_out_2_resp_valid; // @[src/main/scala/system/NutShell.scala 106:24]
  wire [3:0] mmioXbar_io_out_2_resp_bits_cmd; // @[src/main/scala/system/NutShell.scala 106:24]
  wire [63:0] mmioXbar_io_out_2_resp_bits_rdata; // @[src/main/scala/system/NutShell.scala 106:24]
  wire  mmioXbar_DISPLAY_ENABLE; // @[src/main/scala/system/NutShell.scala 106:24]
  wire  clint_clock; // @[src/main/scala/system/NutShell.scala 113:21]
  wire  clint_reset; // @[src/main/scala/system/NutShell.scala 113:21]
  wire  clint_io__in_aw_ready; // @[src/main/scala/system/NutShell.scala 113:21]
  wire  clint_io__in_aw_valid; // @[src/main/scala/system/NutShell.scala 113:21]
  wire [31:0] clint_io__in_aw_bits_addr; // @[src/main/scala/system/NutShell.scala 113:21]
  wire  clint_io__in_w_ready; // @[src/main/scala/system/NutShell.scala 113:21]
  wire  clint_io__in_w_valid; // @[src/main/scala/system/NutShell.scala 113:21]
  wire [63:0] clint_io__in_w_bits_data; // @[src/main/scala/system/NutShell.scala 113:21]
  wire [7:0] clint_io__in_w_bits_strb; // @[src/main/scala/system/NutShell.scala 113:21]
  wire  clint_io__in_b_ready; // @[src/main/scala/system/NutShell.scala 113:21]
  wire  clint_io__in_b_valid; // @[src/main/scala/system/NutShell.scala 113:21]
  wire  clint_io__in_ar_ready; // @[src/main/scala/system/NutShell.scala 113:21]
  wire  clint_io__in_ar_valid; // @[src/main/scala/system/NutShell.scala 113:21]
  wire [31:0] clint_io__in_ar_bits_addr; // @[src/main/scala/system/NutShell.scala 113:21]
  wire  clint_io__in_r_ready; // @[src/main/scala/system/NutShell.scala 113:21]
  wire  clint_io__in_r_valid; // @[src/main/scala/system/NutShell.scala 113:21]
  wire [63:0] clint_io__in_r_bits_data; // @[src/main/scala/system/NutShell.scala 113:21]
  wire  clint_io__extra_mtip; // @[src/main/scala/system/NutShell.scala 113:21]
  wire  clint_io__extra_msip; // @[src/main/scala/system/NutShell.scala 113:21]
  wire  clint_isWFI_0; // @[src/main/scala/system/NutShell.scala 113:21]
  wire  clint_io_extra_mtip; // @[src/main/scala/system/NutShell.scala 113:21]
  wire  clint_io_extra_msip; // @[src/main/scala/system/NutShell.scala 113:21]
  wire  clint_io_in_bridge_clock; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  clint_io_in_bridge_reset; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  clint_io_in_bridge_io_in_req_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  clint_io_in_bridge_io_in_req_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [31:0] clint_io_in_bridge_io_in_req_bits_addr; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [3:0] clint_io_in_bridge_io_in_req_bits_cmd; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [7:0] clint_io_in_bridge_io_in_req_bits_wmask; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [63:0] clint_io_in_bridge_io_in_req_bits_wdata; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  clint_io_in_bridge_io_in_resp_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  clint_io_in_bridge_io_in_resp_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [63:0] clint_io_in_bridge_io_in_resp_bits_rdata; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  clint_io_in_bridge_io_out_aw_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  clint_io_in_bridge_io_out_aw_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [31:0] clint_io_in_bridge_io_out_aw_bits_addr; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  clint_io_in_bridge_io_out_w_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  clint_io_in_bridge_io_out_w_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [63:0] clint_io_in_bridge_io_out_w_bits_data; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [7:0] clint_io_in_bridge_io_out_w_bits_strb; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  clint_io_in_bridge_io_out_b_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  clint_io_in_bridge_io_out_b_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  clint_io_in_bridge_io_out_ar_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  clint_io_in_bridge_io_out_ar_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [31:0] clint_io_in_bridge_io_out_ar_bits_addr; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  clint_io_in_bridge_io_out_r_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  clint_io_in_bridge_io_out_r_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [63:0] clint_io_in_bridge_io_out_r_bits_data; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  plic_clock; // @[src/main/scala/system/NutShell.scala 120:20]
  wire  plic_reset; // @[src/main/scala/system/NutShell.scala 120:20]
  wire  plic_io__in_aw_ready; // @[src/main/scala/system/NutShell.scala 120:20]
  wire  plic_io__in_aw_valid; // @[src/main/scala/system/NutShell.scala 120:20]
  wire [31:0] plic_io__in_aw_bits_addr; // @[src/main/scala/system/NutShell.scala 120:20]
  wire  plic_io__in_w_ready; // @[src/main/scala/system/NutShell.scala 120:20]
  wire  plic_io__in_w_valid; // @[src/main/scala/system/NutShell.scala 120:20]
  wire [63:0] plic_io__in_w_bits_data; // @[src/main/scala/system/NutShell.scala 120:20]
  wire [7:0] plic_io__in_w_bits_strb; // @[src/main/scala/system/NutShell.scala 120:20]
  wire  plic_io__in_b_ready; // @[src/main/scala/system/NutShell.scala 120:20]
  wire  plic_io__in_b_valid; // @[src/main/scala/system/NutShell.scala 120:20]
  wire  plic_io__in_ar_ready; // @[src/main/scala/system/NutShell.scala 120:20]
  wire  plic_io__in_ar_valid; // @[src/main/scala/system/NutShell.scala 120:20]
  wire [31:0] plic_io__in_ar_bits_addr; // @[src/main/scala/system/NutShell.scala 120:20]
  wire  plic_io__in_r_ready; // @[src/main/scala/system/NutShell.scala 120:20]
  wire  plic_io__in_r_valid; // @[src/main/scala/system/NutShell.scala 120:20]
  wire [63:0] plic_io__in_r_bits_data; // @[src/main/scala/system/NutShell.scala 120:20]
  wire  plic_io__extra_intrVec; // @[src/main/scala/system/NutShell.scala 120:20]
  wire  plic_io__extra_meip_0; // @[src/main/scala/system/NutShell.scala 120:20]
  wire  plic_io_extra_meip_0; // @[src/main/scala/system/NutShell.scala 120:20]
  wire  plic_io_in_bridge_clock; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  plic_io_in_bridge_reset; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  plic_io_in_bridge_io_in_req_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  plic_io_in_bridge_io_in_req_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [31:0] plic_io_in_bridge_io_in_req_bits_addr; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [3:0] plic_io_in_bridge_io_in_req_bits_cmd; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [7:0] plic_io_in_bridge_io_in_req_bits_wmask; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [63:0] plic_io_in_bridge_io_in_req_bits_wdata; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  plic_io_in_bridge_io_in_resp_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  plic_io_in_bridge_io_in_resp_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [63:0] plic_io_in_bridge_io_in_resp_bits_rdata; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  plic_io_in_bridge_io_out_aw_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  plic_io_in_bridge_io_out_aw_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [31:0] plic_io_in_bridge_io_out_aw_bits_addr; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  plic_io_in_bridge_io_out_w_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  plic_io_in_bridge_io_out_w_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [63:0] plic_io_in_bridge_io_out_w_bits_data; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [7:0] plic_io_in_bridge_io_out_w_bits_strb; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  plic_io_in_bridge_io_out_b_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  plic_io_in_bridge_io_out_b_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  plic_io_in_bridge_io_out_ar_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  plic_io_in_bridge_io_out_ar_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [31:0] plic_io_in_bridge_io_out_ar_bits_addr; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  plic_io_in_bridge_io_out_r_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  plic_io_in_bridge_io_out_r_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [63:0] plic_io_in_bridge_io_out_r_bits_data; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  reg  plic_io_extra_intrVec_REG; // @[src/main/scala/system/NutShell.scala 122:47]
  reg  plic_io_extra_intrVec_REG_1; // @[src/main/scala/system/NutShell.scala 122:39]
  NutCore nutcore ( // @[src/main/scala/system/NutShell.scala 53:23]
    .clock(nutcore_clock),
    .reset(nutcore_reset),
    .io_imem_mem_req_ready(nutcore_io_imem_mem_req_ready),
    .io_imem_mem_req_valid(nutcore_io_imem_mem_req_valid),
    .io_imem_mem_req_bits_addr(nutcore_io_imem_mem_req_bits_addr),
    .io_imem_mem_req_bits_cmd(nutcore_io_imem_mem_req_bits_cmd),
    .io_imem_mem_req_bits_wdata(nutcore_io_imem_mem_req_bits_wdata),
    .io_imem_mem_resp_valid(nutcore_io_imem_mem_resp_valid),
    .io_imem_mem_resp_bits_cmd(nutcore_io_imem_mem_resp_bits_cmd),
    .io_imem_mem_resp_bits_rdata(nutcore_io_imem_mem_resp_bits_rdata),
    .io_dmem_mem_req_ready(nutcore_io_dmem_mem_req_ready),
    .io_dmem_mem_req_valid(nutcore_io_dmem_mem_req_valid),
    .io_dmem_mem_req_bits_addr(nutcore_io_dmem_mem_req_bits_addr),
    .io_dmem_mem_req_bits_cmd(nutcore_io_dmem_mem_req_bits_cmd),
    .io_dmem_mem_req_bits_wdata(nutcore_io_dmem_mem_req_bits_wdata),
    .io_dmem_mem_resp_valid(nutcore_io_dmem_mem_resp_valid),
    .io_dmem_mem_resp_bits_cmd(nutcore_io_dmem_mem_resp_bits_cmd),
    .io_dmem_mem_resp_bits_rdata(nutcore_io_dmem_mem_resp_bits_rdata),
    .io_dmem_coh_req_ready(nutcore_io_dmem_coh_req_ready),
    .io_dmem_coh_req_valid(nutcore_io_dmem_coh_req_valid),
    .io_dmem_coh_req_bits_addr(nutcore_io_dmem_coh_req_bits_addr),
    .io_dmem_coh_req_bits_wdata(nutcore_io_dmem_coh_req_bits_wdata),
    .io_dmem_coh_resp_valid(nutcore_io_dmem_coh_resp_valid),
    .io_dmem_coh_resp_bits_cmd(nutcore_io_dmem_coh_resp_bits_cmd),
    .io_dmem_coh_resp_bits_rdata(nutcore_io_dmem_coh_resp_bits_rdata),
    .io_mmio_req_ready(nutcore_io_mmio_req_ready),
    .io_mmio_req_valid(nutcore_io_mmio_req_valid),
    .io_mmio_req_bits_addr(nutcore_io_mmio_req_bits_addr),
    .io_mmio_req_bits_size(nutcore_io_mmio_req_bits_size),
    .io_mmio_req_bits_cmd(nutcore_io_mmio_req_bits_cmd),
    .io_mmio_req_bits_wmask(nutcore_io_mmio_req_bits_wmask),
    .io_mmio_req_bits_wdata(nutcore_io_mmio_req_bits_wdata),
    .io_mmio_resp_valid(nutcore_io_mmio_resp_valid),
    .io_mmio_resp_bits_cmd(nutcore_io_mmio_resp_bits_cmd),
    .io_mmio_resp_bits_rdata(nutcore_io_mmio_resp_bits_rdata),
    .io_frontend_req_ready(nutcore_io_frontend_req_ready),
    .io_frontend_req_valid(nutcore_io_frontend_req_valid),
    .io_frontend_req_bits_addr(nutcore_io_frontend_req_bits_addr),
    .io_frontend_req_bits_size(nutcore_io_frontend_req_bits_size),
    .io_frontend_req_bits_cmd(nutcore_io_frontend_req_bits_cmd),
    .io_frontend_req_bits_wmask(nutcore_io_frontend_req_bits_wmask),
    .io_frontend_req_bits_wdata(nutcore_io_frontend_req_bits_wdata),
    .io_frontend_resp_ready(nutcore_io_frontend_resp_ready),
    .io_frontend_resp_valid(nutcore_io_frontend_resp_valid),
    .io_frontend_resp_bits_cmd(nutcore_io_frontend_resp_bits_cmd),
    .io_frontend_resp_bits_rdata(nutcore_io_frontend_resp_bits_rdata),
    .io_extra_meip_0(nutcore_io_extra_meip_0),
    ._WIRE_0(nutcore__WIRE_0),
    .DISPLAY_ENABLE(nutcore_DISPLAY_ENABLE),
    .io_extra_mtip(nutcore_io_extra_mtip),
    .io_extra_msip(nutcore_io_extra_msip)
  );
  CoherenceManager cohMg ( // @[src/main/scala/system/NutShell.scala 54:21]
    .clock(cohMg_clock),
    .reset(cohMg_reset),
    .io_in_req_ready(cohMg_io_in_req_ready),
    .io_in_req_valid(cohMg_io_in_req_valid),
    .io_in_req_bits_addr(cohMg_io_in_req_bits_addr),
    .io_in_req_bits_cmd(cohMg_io_in_req_bits_cmd),
    .io_in_req_bits_wdata(cohMg_io_in_req_bits_wdata),
    .io_in_resp_valid(cohMg_io_in_resp_valid),
    .io_in_resp_bits_cmd(cohMg_io_in_resp_bits_cmd),
    .io_in_resp_bits_rdata(cohMg_io_in_resp_bits_rdata),
    .io_out_mem_req_ready(cohMg_io_out_mem_req_ready),
    .io_out_mem_req_valid(cohMg_io_out_mem_req_valid),
    .io_out_mem_req_bits_addr(cohMg_io_out_mem_req_bits_addr),
    .io_out_mem_req_bits_cmd(cohMg_io_out_mem_req_bits_cmd),
    .io_out_mem_req_bits_wdata(cohMg_io_out_mem_req_bits_wdata),
    .io_out_mem_resp_ready(cohMg_io_out_mem_resp_ready),
    .io_out_mem_resp_valid(cohMg_io_out_mem_resp_valid),
    .io_out_mem_resp_bits_cmd(cohMg_io_out_mem_resp_bits_cmd),
    .io_out_mem_resp_bits_rdata(cohMg_io_out_mem_resp_bits_rdata),
    .io_out_coh_req_ready(cohMg_io_out_coh_req_ready),
    .io_out_coh_req_valid(cohMg_io_out_coh_req_valid),
    .io_out_coh_req_bits_addr(cohMg_io_out_coh_req_bits_addr),
    .io_out_coh_req_bits_wdata(cohMg_io_out_coh_req_bits_wdata),
    .io_out_coh_resp_ready(cohMg_io_out_coh_resp_ready),
    .io_out_coh_resp_valid(cohMg_io_out_coh_resp_valid),
    .io_out_coh_resp_bits_cmd(cohMg_io_out_coh_resp_bits_cmd),
    .io_out_coh_resp_bits_rdata(cohMg_io_out_coh_resp_bits_rdata)
  );
  SimpleBusCrossbarNto1 xbar ( // @[src/main/scala/system/NutShell.scala 55:20]
    .clock(xbar_clock),
    .reset(xbar_reset),
    .io_in_0_req_ready(xbar_io_in_0_req_ready),
    .io_in_0_req_valid(xbar_io_in_0_req_valid),
    .io_in_0_req_bits_addr(xbar_io_in_0_req_bits_addr),
    .io_in_0_req_bits_cmd(xbar_io_in_0_req_bits_cmd),
    .io_in_0_req_bits_wmask(xbar_io_in_0_req_bits_wmask),
    .io_in_0_req_bits_wdata(xbar_io_in_0_req_bits_wdata),
    .io_in_0_resp_valid(xbar_io_in_0_resp_valid),
    .io_in_0_resp_bits_cmd(xbar_io_in_0_resp_bits_cmd),
    .io_in_0_resp_bits_rdata(xbar_io_in_0_resp_bits_rdata),
    .io_in_1_req_ready(xbar_io_in_1_req_ready),
    .io_in_1_req_valid(xbar_io_in_1_req_valid),
    .io_in_1_req_bits_addr(xbar_io_in_1_req_bits_addr),
    .io_in_1_req_bits_size(xbar_io_in_1_req_bits_size),
    .io_in_1_req_bits_cmd(xbar_io_in_1_req_bits_cmd),
    .io_in_1_req_bits_wmask(xbar_io_in_1_req_bits_wmask),
    .io_in_1_req_bits_wdata(xbar_io_in_1_req_bits_wdata),
    .io_in_1_resp_valid(xbar_io_in_1_resp_valid),
    .io_in_1_resp_bits_cmd(xbar_io_in_1_resp_bits_cmd),
    .io_in_1_resp_bits_rdata(xbar_io_in_1_resp_bits_rdata),
    .io_out_req_ready(xbar_io_out_req_ready),
    .io_out_req_valid(xbar_io_out_req_valid),
    .io_out_req_bits_addr(xbar_io_out_req_bits_addr),
    .io_out_req_bits_size(xbar_io_out_req_bits_size),
    .io_out_req_bits_cmd(xbar_io_out_req_bits_cmd),
    .io_out_req_bits_wmask(xbar_io_out_req_bits_wmask),
    .io_out_req_bits_wdata(xbar_io_out_req_bits_wdata),
    .io_out_resp_ready(xbar_io_out_resp_ready),
    .io_out_resp_valid(xbar_io_out_resp_valid),
    .io_out_resp_bits_cmd(xbar_io_out_resp_bits_cmd),
    .io_out_resp_bits_rdata(xbar_io_out_resp_bits_rdata)
  );
  AXI42SimpleBusConverter axi2sb ( // @[src/main/scala/system/NutShell.scala 61:22]
    .clock(axi2sb_clock),
    .reset(axi2sb_reset),
    .io_in_aw_ready(axi2sb_io_in_aw_ready),
    .io_in_aw_valid(axi2sb_io_in_aw_valid),
    .io_in_aw_bits_addr(axi2sb_io_in_aw_bits_addr),
    .io_in_aw_bits_len(axi2sb_io_in_aw_bits_len),
    .io_in_aw_bits_size(axi2sb_io_in_aw_bits_size),
    .io_in_w_ready(axi2sb_io_in_w_ready),
    .io_in_w_valid(axi2sb_io_in_w_valid),
    .io_in_w_bits_data(axi2sb_io_in_w_bits_data),
    .io_in_w_bits_strb(axi2sb_io_in_w_bits_strb),
    .io_in_b_ready(axi2sb_io_in_b_ready),
    .io_in_b_valid(axi2sb_io_in_b_valid),
    .io_in_ar_ready(axi2sb_io_in_ar_ready),
    .io_in_ar_valid(axi2sb_io_in_ar_valid),
    .io_in_ar_bits_addr(axi2sb_io_in_ar_bits_addr),
    .io_in_r_ready(axi2sb_io_in_r_ready),
    .io_in_r_valid(axi2sb_io_in_r_valid),
    .io_in_r_bits_data(axi2sb_io_in_r_bits_data),
    .io_out_req_ready(axi2sb_io_out_req_ready),
    .io_out_req_valid(axi2sb_io_out_req_valid),
    .io_out_req_bits_addr(axi2sb_io_out_req_bits_addr),
    .io_out_req_bits_size(axi2sb_io_out_req_bits_size),
    .io_out_req_bits_cmd(axi2sb_io_out_req_bits_cmd),
    .io_out_req_bits_wmask(axi2sb_io_out_req_bits_wmask),
    .io_out_req_bits_wdata(axi2sb_io_out_req_bits_wdata),
    .io_out_resp_ready(axi2sb_io_out_resp_ready),
    .io_out_resp_valid(axi2sb_io_out_resp_valid),
    .io_out_resp_bits_cmd(axi2sb_io_out_resp_bits_cmd),
    .io_out_resp_bits_rdata(axi2sb_io_out_resp_bits_rdata)
  );
  Prefetcher mem_l2cacheIn_prefetcher ( // @[src/main/scala/system/NutShell.scala 73:30]
    .clock(mem_l2cacheIn_prefetcher_clock),
    .reset(mem_l2cacheIn_prefetcher_reset),
    .io_in_ready(mem_l2cacheIn_prefetcher_io_in_ready),
    .io_in_valid(mem_l2cacheIn_prefetcher_io_in_valid),
    .io_in_bits_addr(mem_l2cacheIn_prefetcher_io_in_bits_addr),
    .io_in_bits_size(mem_l2cacheIn_prefetcher_io_in_bits_size),
    .io_in_bits_cmd(mem_l2cacheIn_prefetcher_io_in_bits_cmd),
    .io_in_bits_wmask(mem_l2cacheIn_prefetcher_io_in_bits_wmask),
    .io_in_bits_wdata(mem_l2cacheIn_prefetcher_io_in_bits_wdata),
    .io_out_ready(mem_l2cacheIn_prefetcher_io_out_ready),
    .io_out_valid(mem_l2cacheIn_prefetcher_io_out_valid),
    .io_out_bits_addr(mem_l2cacheIn_prefetcher_io_out_bits_addr),
    .io_out_bits_size(mem_l2cacheIn_prefetcher_io_out_bits_size),
    .io_out_bits_cmd(mem_l2cacheIn_prefetcher_io_out_bits_cmd),
    .io_out_bits_wmask(mem_l2cacheIn_prefetcher_io_out_bits_wmask),
    .io_out_bits_wdata(mem_l2cacheIn_prefetcher_io_out_bits_wdata),
    .DISPLAY_ENABLE(mem_l2cacheIn_prefetcher_DISPLAY_ENABLE)
  );
  Cache_2 mem_l2cacheOut_cache ( // @[src/main/scala/nutcore/mem/Cache.scala 668:35]
    .clock(mem_l2cacheOut_cache_clock),
    .reset(mem_l2cacheOut_cache_reset),
    .io_in_req_ready(mem_l2cacheOut_cache_io_in_req_ready),
    .io_in_req_valid(mem_l2cacheOut_cache_io_in_req_valid),
    .io_in_req_bits_addr(mem_l2cacheOut_cache_io_in_req_bits_addr),
    .io_in_req_bits_size(mem_l2cacheOut_cache_io_in_req_bits_size),
    .io_in_req_bits_cmd(mem_l2cacheOut_cache_io_in_req_bits_cmd),
    .io_in_req_bits_wmask(mem_l2cacheOut_cache_io_in_req_bits_wmask),
    .io_in_req_bits_wdata(mem_l2cacheOut_cache_io_in_req_bits_wdata),
    .io_in_resp_valid(mem_l2cacheOut_cache_io_in_resp_valid),
    .io_in_resp_bits_cmd(mem_l2cacheOut_cache_io_in_resp_bits_cmd),
    .io_in_resp_bits_rdata(mem_l2cacheOut_cache_io_in_resp_bits_rdata),
    .io_out_mem_req_ready(mem_l2cacheOut_cache_io_out_mem_req_ready),
    .io_out_mem_req_valid(mem_l2cacheOut_cache_io_out_mem_req_valid),
    .io_out_mem_req_bits_addr(mem_l2cacheOut_cache_io_out_mem_req_bits_addr),
    .io_out_mem_req_bits_cmd(mem_l2cacheOut_cache_io_out_mem_req_bits_cmd),
    .io_out_mem_req_bits_wdata(mem_l2cacheOut_cache_io_out_mem_req_bits_wdata),
    .io_out_mem_resp_valid(mem_l2cacheOut_cache_io_out_mem_resp_valid),
    .io_out_mem_resp_bits_cmd(mem_l2cacheOut_cache_io_out_mem_resp_bits_cmd),
    .io_out_mem_resp_bits_rdata(mem_l2cacheOut_cache_io_out_mem_resp_bits_rdata),
    .DISPLAY_ENABLE(mem_l2cacheOut_cache_DISPLAY_ENABLE)
  );
  SimpleBusAddressMapper memAddrMap ( // @[src/main/scala/system/NutShell.scala 93:26]
    .io_in_req_ready(memAddrMap_io_in_req_ready),
    .io_in_req_valid(memAddrMap_io_in_req_valid),
    .io_in_req_bits_addr(memAddrMap_io_in_req_bits_addr),
    .io_in_req_bits_cmd(memAddrMap_io_in_req_bits_cmd),
    .io_in_req_bits_wdata(memAddrMap_io_in_req_bits_wdata),
    .io_in_resp_valid(memAddrMap_io_in_resp_valid),
    .io_in_resp_bits_cmd(memAddrMap_io_in_resp_bits_cmd),
    .io_in_resp_bits_rdata(memAddrMap_io_in_resp_bits_rdata),
    .io_out_req_ready(memAddrMap_io_out_req_ready),
    .io_out_req_valid(memAddrMap_io_out_req_valid),
    .io_out_req_bits_addr(memAddrMap_io_out_req_bits_addr),
    .io_out_req_bits_cmd(memAddrMap_io_out_req_bits_cmd),
    .io_out_req_bits_wdata(memAddrMap_io_out_req_bits_wdata),
    .io_out_resp_valid(memAddrMap_io_out_resp_valid),
    .io_out_resp_bits_cmd(memAddrMap_io_out_resp_bits_cmd),
    .io_out_resp_bits_rdata(memAddrMap_io_out_resp_bits_rdata)
  );
  SimpleBus2AXI4Converter io_mem_bridge ( // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
    .clock(io_mem_bridge_clock),
    .reset(io_mem_bridge_reset),
    .io_in_req_ready(io_mem_bridge_io_in_req_ready),
    .io_in_req_valid(io_mem_bridge_io_in_req_valid),
    .io_in_req_bits_addr(io_mem_bridge_io_in_req_bits_addr),
    .io_in_req_bits_cmd(io_mem_bridge_io_in_req_bits_cmd),
    .io_in_req_bits_wdata(io_mem_bridge_io_in_req_bits_wdata),
    .io_in_resp_valid(io_mem_bridge_io_in_resp_valid),
    .io_in_resp_bits_cmd(io_mem_bridge_io_in_resp_bits_cmd),
    .io_in_resp_bits_rdata(io_mem_bridge_io_in_resp_bits_rdata),
    .io_out_aw_ready(io_mem_bridge_io_out_aw_ready),
    .io_out_aw_valid(io_mem_bridge_io_out_aw_valid),
    .io_out_aw_bits_addr(io_mem_bridge_io_out_aw_bits_addr),
    .io_out_aw_bits_len(io_mem_bridge_io_out_aw_bits_len),
    .io_out_aw_bits_size(io_mem_bridge_io_out_aw_bits_size),
    .io_out_aw_bits_burst(io_mem_bridge_io_out_aw_bits_burst),
    .io_out_w_ready(io_mem_bridge_io_out_w_ready),
    .io_out_w_valid(io_mem_bridge_io_out_w_valid),
    .io_out_w_bits_data(io_mem_bridge_io_out_w_bits_data),
    .io_out_w_bits_last(io_mem_bridge_io_out_w_bits_last),
    .io_out_b_valid(io_mem_bridge_io_out_b_valid),
    .io_out_ar_ready(io_mem_bridge_io_out_ar_ready),
    .io_out_ar_valid(io_mem_bridge_io_out_ar_valid),
    .io_out_ar_bits_addr(io_mem_bridge_io_out_ar_bits_addr),
    .io_out_ar_bits_len(io_mem_bridge_io_out_ar_bits_len),
    .io_out_ar_bits_size(io_mem_bridge_io_out_ar_bits_size),
    .io_out_ar_bits_burst(io_mem_bridge_io_out_ar_bits_burst),
    .io_out_r_valid(io_mem_bridge_io_out_r_valid),
    .io_out_r_bits_data(io_mem_bridge_io_out_r_bits_data),
    .io_out_r_bits_last(io_mem_bridge_io_out_r_bits_last)
  );
  SimpleBusCrossbar1toN mmioXbar ( // @[src/main/scala/system/NutShell.scala 106:24]
    .clock(mmioXbar_clock),
    .reset(mmioXbar_reset),
    .io_in_req_ready(mmioXbar_io_in_req_ready),
    .io_in_req_valid(mmioXbar_io_in_req_valid),
    .io_in_req_bits_addr(mmioXbar_io_in_req_bits_addr),
    .io_in_req_bits_size(mmioXbar_io_in_req_bits_size),
    .io_in_req_bits_cmd(mmioXbar_io_in_req_bits_cmd),
    .io_in_req_bits_wmask(mmioXbar_io_in_req_bits_wmask),
    .io_in_req_bits_wdata(mmioXbar_io_in_req_bits_wdata),
    .io_in_resp_valid(mmioXbar_io_in_resp_valid),
    .io_in_resp_bits_cmd(mmioXbar_io_in_resp_bits_cmd),
    .io_in_resp_bits_rdata(mmioXbar_io_in_resp_bits_rdata),
    .io_out_0_req_ready(mmioXbar_io_out_0_req_ready),
    .io_out_0_req_valid(mmioXbar_io_out_0_req_valid),
    .io_out_0_req_bits_addr(mmioXbar_io_out_0_req_bits_addr),
    .io_out_0_req_bits_cmd(mmioXbar_io_out_0_req_bits_cmd),
    .io_out_0_req_bits_wmask(mmioXbar_io_out_0_req_bits_wmask),
    .io_out_0_req_bits_wdata(mmioXbar_io_out_0_req_bits_wdata),
    .io_out_0_resp_ready(mmioXbar_io_out_0_resp_ready),
    .io_out_0_resp_valid(mmioXbar_io_out_0_resp_valid),
    .io_out_0_resp_bits_rdata(mmioXbar_io_out_0_resp_bits_rdata),
    .io_out_1_req_ready(mmioXbar_io_out_1_req_ready),
    .io_out_1_req_valid(mmioXbar_io_out_1_req_valid),
    .io_out_1_req_bits_addr(mmioXbar_io_out_1_req_bits_addr),
    .io_out_1_req_bits_cmd(mmioXbar_io_out_1_req_bits_cmd),
    .io_out_1_req_bits_wmask(mmioXbar_io_out_1_req_bits_wmask),
    .io_out_1_req_bits_wdata(mmioXbar_io_out_1_req_bits_wdata),
    .io_out_1_resp_ready(mmioXbar_io_out_1_resp_ready),
    .io_out_1_resp_valid(mmioXbar_io_out_1_resp_valid),
    .io_out_1_resp_bits_rdata(mmioXbar_io_out_1_resp_bits_rdata),
    .io_out_2_req_ready(mmioXbar_io_out_2_req_ready),
    .io_out_2_req_valid(mmioXbar_io_out_2_req_valid),
    .io_out_2_req_bits_addr(mmioXbar_io_out_2_req_bits_addr),
    .io_out_2_req_bits_size(mmioXbar_io_out_2_req_bits_size),
    .io_out_2_req_bits_cmd(mmioXbar_io_out_2_req_bits_cmd),
    .io_out_2_req_bits_wmask(mmioXbar_io_out_2_req_bits_wmask),
    .io_out_2_req_bits_wdata(mmioXbar_io_out_2_req_bits_wdata),
    .io_out_2_resp_ready(mmioXbar_io_out_2_resp_ready),
    .io_out_2_resp_valid(mmioXbar_io_out_2_resp_valid),
    .io_out_2_resp_bits_cmd(mmioXbar_io_out_2_resp_bits_cmd),
    .io_out_2_resp_bits_rdata(mmioXbar_io_out_2_resp_bits_rdata),
    .DISPLAY_ENABLE(mmioXbar_DISPLAY_ENABLE)
  );
  AXI4CLINT clint ( // @[src/main/scala/system/NutShell.scala 113:21]
    .clock(clint_clock),
    .reset(clint_reset),
    .io__in_aw_ready(clint_io__in_aw_ready),
    .io__in_aw_valid(clint_io__in_aw_valid),
    .io__in_aw_bits_addr(clint_io__in_aw_bits_addr),
    .io__in_w_ready(clint_io__in_w_ready),
    .io__in_w_valid(clint_io__in_w_valid),
    .io__in_w_bits_data(clint_io__in_w_bits_data),
    .io__in_w_bits_strb(clint_io__in_w_bits_strb),
    .io__in_b_ready(clint_io__in_b_ready),
    .io__in_b_valid(clint_io__in_b_valid),
    .io__in_ar_ready(clint_io__in_ar_ready),
    .io__in_ar_valid(clint_io__in_ar_valid),
    .io__in_ar_bits_addr(clint_io__in_ar_bits_addr),
    .io__in_r_ready(clint_io__in_r_ready),
    .io__in_r_valid(clint_io__in_r_valid),
    .io__in_r_bits_data(clint_io__in_r_bits_data),
    .io__extra_mtip(clint_io__extra_mtip),
    .io__extra_msip(clint_io__extra_msip),
    .isWFI_0(clint_isWFI_0),
    .io_extra_mtip(clint_io_extra_mtip),
    .io_extra_msip(clint_io_extra_msip)
  );
  SimpleBus2AXI4Converter_1 clint_io_in_bridge ( // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
    .clock(clint_io_in_bridge_clock),
    .reset(clint_io_in_bridge_reset),
    .io_in_req_ready(clint_io_in_bridge_io_in_req_ready),
    .io_in_req_valid(clint_io_in_bridge_io_in_req_valid),
    .io_in_req_bits_addr(clint_io_in_bridge_io_in_req_bits_addr),
    .io_in_req_bits_cmd(clint_io_in_bridge_io_in_req_bits_cmd),
    .io_in_req_bits_wmask(clint_io_in_bridge_io_in_req_bits_wmask),
    .io_in_req_bits_wdata(clint_io_in_bridge_io_in_req_bits_wdata),
    .io_in_resp_ready(clint_io_in_bridge_io_in_resp_ready),
    .io_in_resp_valid(clint_io_in_bridge_io_in_resp_valid),
    .io_in_resp_bits_rdata(clint_io_in_bridge_io_in_resp_bits_rdata),
    .io_out_aw_ready(clint_io_in_bridge_io_out_aw_ready),
    .io_out_aw_valid(clint_io_in_bridge_io_out_aw_valid),
    .io_out_aw_bits_addr(clint_io_in_bridge_io_out_aw_bits_addr),
    .io_out_w_ready(clint_io_in_bridge_io_out_w_ready),
    .io_out_w_valid(clint_io_in_bridge_io_out_w_valid),
    .io_out_w_bits_data(clint_io_in_bridge_io_out_w_bits_data),
    .io_out_w_bits_strb(clint_io_in_bridge_io_out_w_bits_strb),
    .io_out_b_ready(clint_io_in_bridge_io_out_b_ready),
    .io_out_b_valid(clint_io_in_bridge_io_out_b_valid),
    .io_out_ar_ready(clint_io_in_bridge_io_out_ar_ready),
    .io_out_ar_valid(clint_io_in_bridge_io_out_ar_valid),
    .io_out_ar_bits_addr(clint_io_in_bridge_io_out_ar_bits_addr),
    .io_out_r_ready(clint_io_in_bridge_io_out_r_ready),
    .io_out_r_valid(clint_io_in_bridge_io_out_r_valid),
    .io_out_r_bits_data(clint_io_in_bridge_io_out_r_bits_data)
  );
  AXI4PLIC plic ( // @[src/main/scala/system/NutShell.scala 120:20]
    .clock(plic_clock),
    .reset(plic_reset),
    .io__in_aw_ready(plic_io__in_aw_ready),
    .io__in_aw_valid(plic_io__in_aw_valid),
    .io__in_aw_bits_addr(plic_io__in_aw_bits_addr),
    .io__in_w_ready(plic_io__in_w_ready),
    .io__in_w_valid(plic_io__in_w_valid),
    .io__in_w_bits_data(plic_io__in_w_bits_data),
    .io__in_w_bits_strb(plic_io__in_w_bits_strb),
    .io__in_b_ready(plic_io__in_b_ready),
    .io__in_b_valid(plic_io__in_b_valid),
    .io__in_ar_ready(plic_io__in_ar_ready),
    .io__in_ar_valid(plic_io__in_ar_valid),
    .io__in_ar_bits_addr(plic_io__in_ar_bits_addr),
    .io__in_r_ready(plic_io__in_r_ready),
    .io__in_r_valid(plic_io__in_r_valid),
    .io__in_r_bits_data(plic_io__in_r_bits_data),
    .io__extra_intrVec(plic_io__extra_intrVec),
    .io__extra_meip_0(plic_io__extra_meip_0),
    .io_extra_meip_0(plic_io_extra_meip_0)
  );
  SimpleBus2AXI4Converter_1 plic_io_in_bridge ( // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
    .clock(plic_io_in_bridge_clock),
    .reset(plic_io_in_bridge_reset),
    .io_in_req_ready(plic_io_in_bridge_io_in_req_ready),
    .io_in_req_valid(plic_io_in_bridge_io_in_req_valid),
    .io_in_req_bits_addr(plic_io_in_bridge_io_in_req_bits_addr),
    .io_in_req_bits_cmd(plic_io_in_bridge_io_in_req_bits_cmd),
    .io_in_req_bits_wmask(plic_io_in_bridge_io_in_req_bits_wmask),
    .io_in_req_bits_wdata(plic_io_in_bridge_io_in_req_bits_wdata),
    .io_in_resp_ready(plic_io_in_bridge_io_in_resp_ready),
    .io_in_resp_valid(plic_io_in_bridge_io_in_resp_valid),
    .io_in_resp_bits_rdata(plic_io_in_bridge_io_in_resp_bits_rdata),
    .io_out_aw_ready(plic_io_in_bridge_io_out_aw_ready),
    .io_out_aw_valid(plic_io_in_bridge_io_out_aw_valid),
    .io_out_aw_bits_addr(plic_io_in_bridge_io_out_aw_bits_addr),
    .io_out_w_ready(plic_io_in_bridge_io_out_w_ready),
    .io_out_w_valid(plic_io_in_bridge_io_out_w_valid),
    .io_out_w_bits_data(plic_io_in_bridge_io_out_w_bits_data),
    .io_out_w_bits_strb(plic_io_in_bridge_io_out_w_bits_strb),
    .io_out_b_ready(plic_io_in_bridge_io_out_b_ready),
    .io_out_b_valid(plic_io_in_bridge_io_out_b_valid),
    .io_out_ar_ready(plic_io_in_bridge_io_out_ar_ready),
    .io_out_ar_valid(plic_io_in_bridge_io_out_ar_valid),
    .io_out_ar_bits_addr(plic_io_in_bridge_io_out_ar_bits_addr),
    .io_out_r_ready(plic_io_in_bridge_io_out_r_ready),
    .io_out_r_valid(plic_io_in_bridge_io_out_r_valid),
    .io_out_r_bits_data(plic_io_in_bridge_io_out_r_bits_data)
  );
  assign io_mem_aw_valid = io_mem_bridge_io_out_aw_valid; // @[src/main/scala/system/NutShell.scala 95:10]
  assign io_mem_aw_bits_addr = io_mem_bridge_io_out_aw_bits_addr; // @[src/main/scala/system/NutShell.scala 95:10]
  assign io_mem_aw_bits_len = io_mem_bridge_io_out_aw_bits_len; // @[src/main/scala/system/NutShell.scala 95:10]
  assign io_mem_aw_bits_size = io_mem_bridge_io_out_aw_bits_size; // @[src/main/scala/system/NutShell.scala 95:10]
  assign io_mem_aw_bits_burst = io_mem_bridge_io_out_aw_bits_burst; // @[src/main/scala/system/NutShell.scala 95:10]
  assign io_mem_w_valid = io_mem_bridge_io_out_w_valid; // @[src/main/scala/system/NutShell.scala 95:10]
  assign io_mem_w_bits_data = io_mem_bridge_io_out_w_bits_data; // @[src/main/scala/system/NutShell.scala 95:10]
  assign io_mem_w_bits_last = io_mem_bridge_io_out_w_bits_last; // @[src/main/scala/system/NutShell.scala 95:10]
  assign io_mem_ar_valid = io_mem_bridge_io_out_ar_valid; // @[src/main/scala/system/NutShell.scala 95:10]
  assign io_mem_ar_bits_addr = io_mem_bridge_io_out_ar_bits_addr; // @[src/main/scala/system/NutShell.scala 95:10]
  assign io_mem_ar_bits_len = io_mem_bridge_io_out_ar_bits_len; // @[src/main/scala/system/NutShell.scala 95:10]
  assign io_mmio_req_valid = mmioXbar_io_out_2_req_valid; // @[src/main/scala/system/NutShell.scala 111:18]
  assign io_mmio_req_bits_addr = mmioXbar_io_out_2_req_bits_addr; // @[src/main/scala/system/NutShell.scala 111:18]
  assign io_mmio_req_bits_size = mmioXbar_io_out_2_req_bits_size; // @[src/main/scala/system/NutShell.scala 111:18]
  assign io_mmio_req_bits_cmd = mmioXbar_io_out_2_req_bits_cmd; // @[src/main/scala/system/NutShell.scala 111:18]
  assign io_mmio_req_bits_wmask = mmioXbar_io_out_2_req_bits_wmask; // @[src/main/scala/system/NutShell.scala 111:18]
  assign io_mmio_req_bits_wdata = mmioXbar_io_out_2_req_bits_wdata; // @[src/main/scala/system/NutShell.scala 111:18]
  assign io_mmio_resp_ready = mmioXbar_io_out_2_resp_ready; // @[src/main/scala/system/NutShell.scala 111:18]
  assign io_frontend_aw_ready = axi2sb_io_in_aw_ready; // @[src/main/scala/system/NutShell.scala 62:16]
  assign io_frontend_w_ready = axi2sb_io_in_w_ready; // @[src/main/scala/system/NutShell.scala 62:16]
  assign io_frontend_b_valid = axi2sb_io_in_b_valid; // @[src/main/scala/system/NutShell.scala 62:16]
  assign io_frontend_ar_ready = axi2sb_io_in_ar_ready; // @[src/main/scala/system/NutShell.scala 62:16]
  assign io_frontend_r_valid = axi2sb_io_in_r_valid; // @[src/main/scala/system/NutShell.scala 62:16]
  assign io_frontend_r_bits_data = axi2sb_io_in_r_bits_data; // @[src/main/scala/system/NutShell.scala 62:16]
  assign nutcore_clock = clock;
  assign nutcore_reset = reset;
  assign nutcore_io_imem_mem_req_ready = cohMg_io_in_req_ready; // @[src/main/scala/system/NutShell.scala 56:15]
  assign nutcore_io_imem_mem_resp_valid = cohMg_io_in_resp_valid; // @[src/main/scala/system/NutShell.scala 56:15]
  assign nutcore_io_imem_mem_resp_bits_cmd = cohMg_io_in_resp_bits_cmd; // @[src/main/scala/system/NutShell.scala 56:15]
  assign nutcore_io_imem_mem_resp_bits_rdata = cohMg_io_in_resp_bits_rdata; // @[src/main/scala/system/NutShell.scala 56:15]
  assign nutcore_io_dmem_mem_req_ready = xbar_io_in_1_req_ready; // @[src/main/scala/system/NutShell.scala 59:17]
  assign nutcore_io_dmem_mem_resp_valid = xbar_io_in_1_resp_valid; // @[src/main/scala/system/NutShell.scala 59:17]
  assign nutcore_io_dmem_mem_resp_bits_cmd = xbar_io_in_1_resp_bits_cmd; // @[src/main/scala/system/NutShell.scala 59:17]
  assign nutcore_io_dmem_mem_resp_bits_rdata = xbar_io_in_1_resp_bits_rdata; // @[src/main/scala/system/NutShell.scala 59:17]
  assign nutcore_io_dmem_coh_req_valid = cohMg_io_out_coh_req_valid; // @[src/main/scala/system/NutShell.scala 57:23]
  assign nutcore_io_dmem_coh_req_bits_addr = cohMg_io_out_coh_req_bits_addr; // @[src/main/scala/system/NutShell.scala 57:23]
  assign nutcore_io_dmem_coh_req_bits_wdata = cohMg_io_out_coh_req_bits_wdata; // @[src/main/scala/system/NutShell.scala 57:23]
  assign nutcore_io_mmio_req_ready = mmioXbar_io_in_req_ready; // @[src/main/scala/system/NutShell.scala 107:18]
  assign nutcore_io_mmio_resp_valid = mmioXbar_io_in_resp_valid; // @[src/main/scala/system/NutShell.scala 107:18]
  assign nutcore_io_mmio_resp_bits_cmd = mmioXbar_io_in_resp_bits_cmd; // @[src/main/scala/system/NutShell.scala 107:18]
  assign nutcore_io_mmio_resp_bits_rdata = mmioXbar_io_in_resp_bits_rdata; // @[src/main/scala/system/NutShell.scala 107:18]
  assign nutcore_io_frontend_req_valid = axi2sb_io_out_req_valid; // @[src/main/scala/system/NutShell.scala 63:23]
  assign nutcore_io_frontend_req_bits_addr = axi2sb_io_out_req_bits_addr; // @[src/main/scala/system/NutShell.scala 63:23]
  assign nutcore_io_frontend_req_bits_size = axi2sb_io_out_req_bits_size; // @[src/main/scala/system/NutShell.scala 63:23]
  assign nutcore_io_frontend_req_bits_cmd = axi2sb_io_out_req_bits_cmd; // @[src/main/scala/system/NutShell.scala 63:23]
  assign nutcore_io_frontend_req_bits_wmask = axi2sb_io_out_req_bits_wmask; // @[src/main/scala/system/NutShell.scala 63:23]
  assign nutcore_io_frontend_req_bits_wdata = axi2sb_io_out_req_bits_wdata; // @[src/main/scala/system/NutShell.scala 63:23]
  assign nutcore_io_frontend_resp_ready = axi2sb_io_out_resp_ready; // @[src/main/scala/system/NutShell.scala 63:23]
  assign nutcore_io_extra_meip_0 = plic_io_extra_meip_0;
  assign nutcore_DISPLAY_ENABLE = _WIRE_4;
  assign nutcore_io_extra_mtip = clint_io_extra_mtip;
  assign nutcore_io_extra_msip = clint_io_extra_msip;
  assign cohMg_clock = clock;
  assign cohMg_reset = reset;
  assign cohMg_io_in_req_valid = nutcore_io_imem_mem_req_valid; // @[src/main/scala/system/NutShell.scala 56:15]
  assign cohMg_io_in_req_bits_addr = nutcore_io_imem_mem_req_bits_addr; // @[src/main/scala/system/NutShell.scala 56:15]
  assign cohMg_io_in_req_bits_cmd = nutcore_io_imem_mem_req_bits_cmd; // @[src/main/scala/system/NutShell.scala 56:15]
  assign cohMg_io_in_req_bits_wdata = nutcore_io_imem_mem_req_bits_wdata; // @[src/main/scala/system/NutShell.scala 56:15]
  assign cohMg_io_out_mem_req_ready = xbar_io_in_0_req_ready; // @[src/main/scala/system/NutShell.scala 58:17]
  assign cohMg_io_out_mem_resp_valid = xbar_io_in_0_resp_valid; // @[src/main/scala/system/NutShell.scala 58:17]
  assign cohMg_io_out_mem_resp_bits_cmd = xbar_io_in_0_resp_bits_cmd; // @[src/main/scala/system/NutShell.scala 58:17]
  assign cohMg_io_out_mem_resp_bits_rdata = xbar_io_in_0_resp_bits_rdata; // @[src/main/scala/system/NutShell.scala 58:17]
  assign cohMg_io_out_coh_req_ready = nutcore_io_dmem_coh_req_ready; // @[src/main/scala/system/NutShell.scala 57:23]
  assign cohMg_io_out_coh_resp_valid = nutcore_io_dmem_coh_resp_valid; // @[src/main/scala/system/NutShell.scala 57:23]
  assign cohMg_io_out_coh_resp_bits_cmd = nutcore_io_dmem_coh_resp_bits_cmd; // @[src/main/scala/system/NutShell.scala 57:23]
  assign cohMg_io_out_coh_resp_bits_rdata = nutcore_io_dmem_coh_resp_bits_rdata; // @[src/main/scala/system/NutShell.scala 57:23]
  assign xbar_clock = clock;
  assign xbar_reset = reset;
  assign xbar_io_in_0_req_valid = cohMg_io_out_mem_req_valid; // @[src/main/scala/system/NutShell.scala 58:17]
  assign xbar_io_in_0_req_bits_addr = cohMg_io_out_mem_req_bits_addr; // @[src/main/scala/system/NutShell.scala 58:17]
  assign xbar_io_in_0_req_bits_cmd = cohMg_io_out_mem_req_bits_cmd; // @[src/main/scala/system/NutShell.scala 58:17]
  assign xbar_io_in_0_req_bits_wmask = 8'hff; // @[src/main/scala/system/NutShell.scala 58:17]
  assign xbar_io_in_0_req_bits_wdata = cohMg_io_out_mem_req_bits_wdata; // @[src/main/scala/system/NutShell.scala 58:17]
  assign xbar_io_in_1_req_valid = nutcore_io_dmem_mem_req_valid; // @[src/main/scala/system/NutShell.scala 59:17]
  assign xbar_io_in_1_req_bits_addr = nutcore_io_dmem_mem_req_bits_addr; // @[src/main/scala/system/NutShell.scala 59:17]
  assign xbar_io_in_1_req_bits_size = 3'h3; // @[src/main/scala/system/NutShell.scala 59:17]
  assign xbar_io_in_1_req_bits_cmd = nutcore_io_dmem_mem_req_bits_cmd; // @[src/main/scala/system/NutShell.scala 59:17]
  assign xbar_io_in_1_req_bits_wmask = 8'hff; // @[src/main/scala/system/NutShell.scala 59:17]
  assign xbar_io_in_1_req_bits_wdata = nutcore_io_dmem_mem_req_bits_wdata; // @[src/main/scala/system/NutShell.scala 59:17]
  assign xbar_io_out_req_ready = mem_l2cacheIn_prefetcher_io_in_ready; // @[src/main/scala/system/NutShell.scala 75:24]
  assign xbar_io_out_resp_valid = mem_l2cacheOut_cache_io_in_resp_valid; // @[src/main/scala/nutcore/mem/Cache.scala 674:17 src/main/scala/system/NutShell.scala 74:27]
  assign xbar_io_out_resp_bits_cmd = mem_l2cacheOut_cache_io_in_resp_bits_cmd; // @[src/main/scala/nutcore/mem/Cache.scala 674:17 src/main/scala/system/NutShell.scala 74:27]
  assign xbar_io_out_resp_bits_rdata = mem_l2cacheOut_cache_io_in_resp_bits_rdata; // @[src/main/scala/nutcore/mem/Cache.scala 674:17 src/main/scala/system/NutShell.scala 74:27]
  assign axi2sb_clock = clock;
  assign axi2sb_reset = reset;
  assign axi2sb_io_in_aw_valid = io_frontend_aw_valid; // @[src/main/scala/system/NutShell.scala 62:16]
  assign axi2sb_io_in_aw_bits_addr = io_frontend_aw_bits_addr; // @[src/main/scala/system/NutShell.scala 62:16]
  assign axi2sb_io_in_aw_bits_len = io_frontend_aw_bits_len; // @[src/main/scala/system/NutShell.scala 62:16]
  assign axi2sb_io_in_aw_bits_size = io_frontend_aw_bits_size; // @[src/main/scala/system/NutShell.scala 62:16]
  assign axi2sb_io_in_w_valid = io_frontend_w_valid; // @[src/main/scala/system/NutShell.scala 62:16]
  assign axi2sb_io_in_w_bits_data = io_frontend_w_bits_data; // @[src/main/scala/system/NutShell.scala 62:16]
  assign axi2sb_io_in_w_bits_strb = io_frontend_w_bits_strb; // @[src/main/scala/system/NutShell.scala 62:16]
  assign axi2sb_io_in_b_ready = io_frontend_b_ready; // @[src/main/scala/system/NutShell.scala 62:16]
  assign axi2sb_io_in_ar_valid = io_frontend_ar_valid; // @[src/main/scala/system/NutShell.scala 62:16]
  assign axi2sb_io_in_ar_bits_addr = io_frontend_ar_bits_addr; // @[src/main/scala/system/NutShell.scala 62:16]
  assign axi2sb_io_in_r_ready = io_frontend_r_ready; // @[src/main/scala/system/NutShell.scala 62:16]
  assign axi2sb_io_out_req_ready = nutcore_io_frontend_req_ready; // @[src/main/scala/system/NutShell.scala 63:23]
  assign axi2sb_io_out_resp_valid = nutcore_io_frontend_resp_valid; // @[src/main/scala/system/NutShell.scala 63:23]
  assign axi2sb_io_out_resp_bits_cmd = nutcore_io_frontend_resp_bits_cmd; // @[src/main/scala/system/NutShell.scala 63:23]
  assign axi2sb_io_out_resp_bits_rdata = nutcore_io_frontend_resp_bits_rdata; // @[src/main/scala/system/NutShell.scala 63:23]
  assign mem_l2cacheIn_prefetcher_clock = clock;
  assign mem_l2cacheIn_prefetcher_reset = reset;
  assign mem_l2cacheIn_prefetcher_io_in_valid = xbar_io_out_req_valid; // @[src/main/scala/system/NutShell.scala 75:24]
  assign mem_l2cacheIn_prefetcher_io_in_bits_addr = xbar_io_out_req_bits_addr; // @[src/main/scala/system/NutShell.scala 75:24]
  assign mem_l2cacheIn_prefetcher_io_in_bits_size = xbar_io_out_req_bits_size; // @[src/main/scala/system/NutShell.scala 75:24]
  assign mem_l2cacheIn_prefetcher_io_in_bits_cmd = xbar_io_out_req_bits_cmd; // @[src/main/scala/system/NutShell.scala 75:24]
  assign mem_l2cacheIn_prefetcher_io_in_bits_wmask = xbar_io_out_req_bits_wmask; // @[src/main/scala/system/NutShell.scala 75:24]
  assign mem_l2cacheIn_prefetcher_io_in_bits_wdata = xbar_io_out_req_bits_wdata; // @[src/main/scala/system/NutShell.scala 75:24]
  assign mem_l2cacheIn_prefetcher_io_out_ready = mem_l2cacheOut_cache_io_in_req_ready; // @[src/main/scala/nutcore/mem/Cache.scala 674:17 src/main/scala/system/NutShell.scala 74:27]
  assign mem_l2cacheIn_prefetcher_DISPLAY_ENABLE = _WIRE_4;
  assign mem_l2cacheOut_cache_clock = clock;
  assign mem_l2cacheOut_cache_reset = reset;
  assign mem_l2cacheOut_cache_io_in_req_valid = mem_l2cacheIn_prefetcher_io_out_valid; // @[src/main/scala/system/NutShell.scala 74:27 76:21]
  assign mem_l2cacheOut_cache_io_in_req_bits_addr = mem_l2cacheIn_prefetcher_io_out_bits_addr; // @[src/main/scala/system/NutShell.scala 74:27 76:21]
  assign mem_l2cacheOut_cache_io_in_req_bits_size = mem_l2cacheIn_prefetcher_io_out_bits_size; // @[src/main/scala/system/NutShell.scala 74:27 76:21]
  assign mem_l2cacheOut_cache_io_in_req_bits_cmd = mem_l2cacheIn_prefetcher_io_out_bits_cmd; // @[src/main/scala/system/NutShell.scala 74:27 76:21]
  assign mem_l2cacheOut_cache_io_in_req_bits_wmask = mem_l2cacheIn_prefetcher_io_out_bits_wmask; // @[src/main/scala/system/NutShell.scala 74:27 76:21]
  assign mem_l2cacheOut_cache_io_in_req_bits_wdata = mem_l2cacheIn_prefetcher_io_out_bits_wdata; // @[src/main/scala/system/NutShell.scala 74:27 76:21]
  assign mem_l2cacheOut_cache_io_out_mem_req_ready = memAddrMap_io_in_req_ready; // @[src/main/scala/system/NutShell.scala 71:26 94:20]
  assign mem_l2cacheOut_cache_io_out_mem_resp_valid = memAddrMap_io_in_resp_valid; // @[src/main/scala/system/NutShell.scala 71:26 94:20]
  assign mem_l2cacheOut_cache_io_out_mem_resp_bits_cmd = memAddrMap_io_in_resp_bits_cmd; // @[src/main/scala/system/NutShell.scala 71:26 94:20]
  assign mem_l2cacheOut_cache_io_out_mem_resp_bits_rdata = memAddrMap_io_in_resp_bits_rdata; // @[src/main/scala/system/NutShell.scala 71:26 94:20]
  assign mem_l2cacheOut_cache_DISPLAY_ENABLE = _WIRE_4;
  assign memAddrMap_io_in_req_valid = mem_l2cacheOut_cache_io_out_mem_req_valid; // @[src/main/scala/system/NutShell.scala 71:26 81:16]
  assign memAddrMap_io_in_req_bits_addr = mem_l2cacheOut_cache_io_out_mem_req_bits_addr; // @[src/main/scala/system/NutShell.scala 71:26 81:16]
  assign memAddrMap_io_in_req_bits_cmd = mem_l2cacheOut_cache_io_out_mem_req_bits_cmd; // @[src/main/scala/system/NutShell.scala 71:26 81:16]
  assign memAddrMap_io_in_req_bits_wdata = mem_l2cacheOut_cache_io_out_mem_req_bits_wdata; // @[src/main/scala/system/NutShell.scala 71:26 81:16]
  assign memAddrMap_io_out_req_ready = io_mem_bridge_io_in_req_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign memAddrMap_io_out_resp_valid = io_mem_bridge_io_in_resp_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign memAddrMap_io_out_resp_bits_cmd = io_mem_bridge_io_in_resp_bits_cmd; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign memAddrMap_io_out_resp_bits_rdata = io_mem_bridge_io_in_resp_bits_rdata; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign io_mem_bridge_clock = clock;
  assign io_mem_bridge_reset = reset;
  assign io_mem_bridge_io_in_req_valid = memAddrMap_io_out_req_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign io_mem_bridge_io_in_req_bits_addr = memAddrMap_io_out_req_bits_addr; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign io_mem_bridge_io_in_req_bits_cmd = memAddrMap_io_out_req_bits_cmd; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign io_mem_bridge_io_in_req_bits_wdata = memAddrMap_io_out_req_bits_wdata; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign io_mem_bridge_io_out_aw_ready = io_mem_aw_ready; // @[src/main/scala/system/NutShell.scala 95:10]
  assign io_mem_bridge_io_out_w_ready = io_mem_w_ready; // @[src/main/scala/system/NutShell.scala 95:10]
  assign io_mem_bridge_io_out_b_valid = io_mem_b_valid; // @[src/main/scala/system/NutShell.scala 95:10]
  assign io_mem_bridge_io_out_ar_ready = io_mem_ar_ready; // @[src/main/scala/system/NutShell.scala 95:10]
  assign io_mem_bridge_io_out_r_valid = io_mem_r_valid; // @[src/main/scala/system/NutShell.scala 95:10]
  assign io_mem_bridge_io_out_r_bits_data = io_mem_r_bits_data; // @[src/main/scala/system/NutShell.scala 95:10]
  assign io_mem_bridge_io_out_r_bits_last = io_mem_r_bits_last; // @[src/main/scala/system/NutShell.scala 95:10]
  assign mmioXbar_clock = clock;
  assign mmioXbar_reset = reset;
  assign mmioXbar_io_in_req_valid = nutcore_io_mmio_req_valid; // @[src/main/scala/system/NutShell.scala 107:18]
  assign mmioXbar_io_in_req_bits_addr = nutcore_io_mmio_req_bits_addr; // @[src/main/scala/system/NutShell.scala 107:18]
  assign mmioXbar_io_in_req_bits_size = nutcore_io_mmio_req_bits_size; // @[src/main/scala/system/NutShell.scala 107:18]
  assign mmioXbar_io_in_req_bits_cmd = nutcore_io_mmio_req_bits_cmd; // @[src/main/scala/system/NutShell.scala 107:18]
  assign mmioXbar_io_in_req_bits_wmask = nutcore_io_mmio_req_bits_wmask; // @[src/main/scala/system/NutShell.scala 107:18]
  assign mmioXbar_io_in_req_bits_wdata = nutcore_io_mmio_req_bits_wdata; // @[src/main/scala/system/NutShell.scala 107:18]
  assign mmioXbar_io_out_0_req_ready = clint_io_in_bridge_io_in_req_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign mmioXbar_io_out_0_resp_valid = clint_io_in_bridge_io_in_resp_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign mmioXbar_io_out_0_resp_bits_rdata = clint_io_in_bridge_io_in_resp_bits_rdata; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign mmioXbar_io_out_1_req_ready = plic_io_in_bridge_io_in_req_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign mmioXbar_io_out_1_resp_valid = plic_io_in_bridge_io_in_resp_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign mmioXbar_io_out_1_resp_bits_rdata = plic_io_in_bridge_io_in_resp_bits_rdata; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign mmioXbar_io_out_2_req_ready = io_mmio_req_ready; // @[src/main/scala/system/NutShell.scala 111:18]
  assign mmioXbar_io_out_2_resp_valid = io_mmio_resp_valid; // @[src/main/scala/system/NutShell.scala 111:18]
  assign mmioXbar_io_out_2_resp_bits_cmd = io_mmio_resp_bits_cmd; // @[src/main/scala/system/NutShell.scala 111:18]
  assign mmioXbar_io_out_2_resp_bits_rdata = io_mmio_resp_bits_rdata; // @[src/main/scala/system/NutShell.scala 111:18]
  assign mmioXbar_DISPLAY_ENABLE = _WIRE_4;
  assign clint_clock = clock;
  assign clint_reset = reset;
  assign clint_io__in_aw_valid = clint_io_in_bridge_io_out_aw_valid; // @[src/main/scala/system/NutShell.scala 114:15]
  assign clint_io__in_aw_bits_addr = clint_io_in_bridge_io_out_aw_bits_addr; // @[src/main/scala/system/NutShell.scala 114:15]
  assign clint_io__in_w_valid = clint_io_in_bridge_io_out_w_valid; // @[src/main/scala/system/NutShell.scala 114:15]
  assign clint_io__in_w_bits_data = clint_io_in_bridge_io_out_w_bits_data; // @[src/main/scala/system/NutShell.scala 114:15]
  assign clint_io__in_w_bits_strb = clint_io_in_bridge_io_out_w_bits_strb; // @[src/main/scala/system/NutShell.scala 114:15]
  assign clint_io__in_b_ready = clint_io_in_bridge_io_out_b_ready; // @[src/main/scala/system/NutShell.scala 114:15]
  assign clint_io__in_ar_valid = clint_io_in_bridge_io_out_ar_valid; // @[src/main/scala/system/NutShell.scala 114:15]
  assign clint_io__in_ar_bits_addr = clint_io_in_bridge_io_out_ar_bits_addr; // @[src/main/scala/system/NutShell.scala 114:15]
  assign clint_io__in_r_ready = clint_io_in_bridge_io_out_r_ready; // @[src/main/scala/system/NutShell.scala 114:15]
  assign clint_isWFI_0 = nutcore__WIRE_0;
  assign clint_io_in_bridge_clock = clock;
  assign clint_io_in_bridge_reset = reset;
  assign clint_io_in_bridge_io_in_req_valid = mmioXbar_io_out_0_req_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign clint_io_in_bridge_io_in_req_bits_addr = mmioXbar_io_out_0_req_bits_addr; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign clint_io_in_bridge_io_in_req_bits_cmd = mmioXbar_io_out_0_req_bits_cmd; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign clint_io_in_bridge_io_in_req_bits_wmask = mmioXbar_io_out_0_req_bits_wmask; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign clint_io_in_bridge_io_in_req_bits_wdata = mmioXbar_io_out_0_req_bits_wdata; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign clint_io_in_bridge_io_in_resp_ready = mmioXbar_io_out_0_resp_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign clint_io_in_bridge_io_out_aw_ready = clint_io__in_aw_ready; // @[src/main/scala/system/NutShell.scala 114:15]
  assign clint_io_in_bridge_io_out_w_ready = clint_io__in_w_ready; // @[src/main/scala/system/NutShell.scala 114:15]
  assign clint_io_in_bridge_io_out_b_valid = clint_io__in_b_valid; // @[src/main/scala/system/NutShell.scala 114:15]
  assign clint_io_in_bridge_io_out_ar_ready = clint_io__in_ar_ready; // @[src/main/scala/system/NutShell.scala 114:15]
  assign clint_io_in_bridge_io_out_r_valid = clint_io__in_r_valid; // @[src/main/scala/system/NutShell.scala 114:15]
  assign clint_io_in_bridge_io_out_r_bits_data = clint_io__in_r_bits_data; // @[src/main/scala/system/NutShell.scala 114:15]
  assign plic_clock = clock;
  assign plic_reset = reset;
  assign plic_io__in_aw_valid = plic_io_in_bridge_io_out_aw_valid; // @[src/main/scala/system/NutShell.scala 121:14]
  assign plic_io__in_aw_bits_addr = plic_io_in_bridge_io_out_aw_bits_addr; // @[src/main/scala/system/NutShell.scala 121:14]
  assign plic_io__in_w_valid = plic_io_in_bridge_io_out_w_valid; // @[src/main/scala/system/NutShell.scala 121:14]
  assign plic_io__in_w_bits_data = plic_io_in_bridge_io_out_w_bits_data; // @[src/main/scala/system/NutShell.scala 121:14]
  assign plic_io__in_w_bits_strb = plic_io_in_bridge_io_out_w_bits_strb; // @[src/main/scala/system/NutShell.scala 121:14]
  assign plic_io__in_b_ready = plic_io_in_bridge_io_out_b_ready; // @[src/main/scala/system/NutShell.scala 121:14]
  assign plic_io__in_ar_valid = plic_io_in_bridge_io_out_ar_valid; // @[src/main/scala/system/NutShell.scala 121:14]
  assign plic_io__in_ar_bits_addr = plic_io_in_bridge_io_out_ar_bits_addr; // @[src/main/scala/system/NutShell.scala 121:14]
  assign plic_io__in_r_ready = plic_io_in_bridge_io_out_r_ready; // @[src/main/scala/system/NutShell.scala 121:14]
  assign plic_io__extra_intrVec = plic_io_extra_intrVec_REG_1; // @[src/main/scala/system/NutShell.scala 122:29]
  assign plic_io_in_bridge_clock = clock;
  assign plic_io_in_bridge_reset = reset;
  assign plic_io_in_bridge_io_in_req_valid = mmioXbar_io_out_1_req_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign plic_io_in_bridge_io_in_req_bits_addr = mmioXbar_io_out_1_req_bits_addr; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign plic_io_in_bridge_io_in_req_bits_cmd = mmioXbar_io_out_1_req_bits_cmd; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign plic_io_in_bridge_io_in_req_bits_wmask = mmioXbar_io_out_1_req_bits_wmask; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign plic_io_in_bridge_io_in_req_bits_wdata = mmioXbar_io_out_1_req_bits_wdata; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign plic_io_in_bridge_io_in_resp_ready = mmioXbar_io_out_1_resp_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign plic_io_in_bridge_io_out_aw_ready = plic_io__in_aw_ready; // @[src/main/scala/system/NutShell.scala 121:14]
  assign plic_io_in_bridge_io_out_w_ready = plic_io__in_w_ready; // @[src/main/scala/system/NutShell.scala 121:14]
  assign plic_io_in_bridge_io_out_b_valid = plic_io__in_b_valid; // @[src/main/scala/system/NutShell.scala 121:14]
  assign plic_io_in_bridge_io_out_ar_ready = plic_io__in_ar_ready; // @[src/main/scala/system/NutShell.scala 121:14]
  assign plic_io_in_bridge_io_out_r_valid = plic_io__in_r_valid; // @[src/main/scala/system/NutShell.scala 121:14]
  assign plic_io_in_bridge_io_out_r_bits_data = plic_io__in_r_bits_data; // @[src/main/scala/system/NutShell.scala 121:14]
  always @(posedge clock) begin
    plic_io_extra_intrVec_REG <= io_meip; // @[src/main/scala/system/NutShell.scala 122:47]
    plic_io_extra_intrVec_REG_1 <= plic_io_extra_intrVec_REG; // @[src/main/scala/system/NutShell.scala 122:39]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  plic_io_extra_intrVec_REG = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  plic_io_extra_intrVec_REG_1 = _RAND_1[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module SynthesizableDifftestMem(
  input         clock,
  input         read_valid, // @[difftest/src/main/scala/common/Mem.scala 160:16]
  input  [63:0] read_index, // @[difftest/src/main/scala/common/Mem.scala 160:16]
  output [63:0] read_data_0, // @[difftest/src/main/scala/common/Mem.scala 160:16]
  input         write_valid, // @[difftest/src/main/scala/common/Mem.scala 165:17]
  input  [63:0] write_index, // @[difftest/src/main/scala/common/Mem.scala 165:17]
  input  [63:0] write_data_0 // @[difftest/src/main/scala/common/Mem.scala 165:17]
);
`ifdef RANDOMIZE_MEM_INIT
  reg [63:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg /* sparse */ [63:0] mem [0:16777215]; // @[difftest/src/main/scala/common/Mem.scala 273:16]
  wire  mem_read_data_0_MPORT_en; // @[difftest/src/main/scala/common/Mem.scala 273:16]
  wire [23:0] mem_read_data_0_MPORT_addr; // @[difftest/src/main/scala/common/Mem.scala 273:16]
  wire [63:0] mem_read_data_0_MPORT_data; // @[difftest/src/main/scala/common/Mem.scala 273:16]
  wire  mem_MPORT_1_en; // @[difftest/src/main/scala/common/Mem.scala 273:16]
  wire [23:0] mem_MPORT_1_addr; // @[difftest/src/main/scala/common/Mem.scala 273:16]
  wire [63:0] mem_MPORT_1_data; // @[difftest/src/main/scala/common/Mem.scala 273:16]
  wire [63:0] mem_MPORT_data; // @[difftest/src/main/scala/common/Mem.scala 273:16]
  wire [23:0] mem_MPORT_addr; // @[difftest/src/main/scala/common/Mem.scala 273:16]
  wire  mem_MPORT_mask; // @[difftest/src/main/scala/common/Mem.scala 273:16]
  wire  mem_MPORT_en; // @[difftest/src/main/scala/common/Mem.scala 273:16]
  wire [64:0] _r_index_T = read_index * 1'h1; // @[difftest/src/main/scala/common/Mem.scala 276:30]
  wire [65:0] _r_index_T_1 = {{1'd0}, _r_index_T}; // @[difftest/src/main/scala/common/Mem.scala 276:43]
  wire [64:0] r_index = _r_index_T_1[64:0]; // @[difftest/src/main/scala/common/Mem.scala 276:43]
  reg [63:0] read_data_0_r; // @[difftest/src/main/scala/common/Mem.scala 277:30]
  wire [64:0] _w_index_T = write_index * 1'h1; // @[difftest/src/main/scala/common/Mem.scala 279:31]
  wire [65:0] _w_index_T_1 = {{1'd0}, _w_index_T}; // @[difftest/src/main/scala/common/Mem.scala 279:44]
  wire [64:0] w_index = _w_index_T_1[64:0]; // @[difftest/src/main/scala/common/Mem.scala 279:44]
  DifftestMemInitializer initializer ( // @[difftest/src/main/scala/common/Mem.scala 285:27]
  );
  assign mem_read_data_0_MPORT_en = 1'h1;
  assign mem_read_data_0_MPORT_addr = r_index[23:0];
  assign mem_read_data_0_MPORT_data = mem[mem_read_data_0_MPORT_addr]; // @[difftest/src/main/scala/common/Mem.scala 273:16]
  assign mem_MPORT_1_en = write_valid;
  assign mem_MPORT_1_addr = w_index[23:0];
  assign mem_MPORT_1_data = mem[mem_MPORT_1_addr]; // @[difftest/src/main/scala/common/Mem.scala 273:16]
  assign mem_MPORT_data = write_data_0;
  assign mem_MPORT_addr = w_index[23:0];
  assign mem_MPORT_mask = 1'h1;
  assign mem_MPORT_en = write_valid;
  assign read_data_0 = read_data_0_r; // @[difftest/src/main/scala/common/Mem.scala 277:18]
  always @(posedge clock) begin
    if (mem_MPORT_en & mem_MPORT_mask) begin
      mem[mem_MPORT_addr] <= mem_MPORT_data; // @[difftest/src/main/scala/common/Mem.scala 273:16]
    end
    if (read_valid) begin // @[difftest/src/main/scala/common/Mem.scala 277:30]
      read_data_0_r <= mem_read_data_0_MPORT_data; // @[difftest/src/main/scala/common/Mem.scala 277:30]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {2{`RANDOM}};
  for (initvar = 0; initvar < 16777216; initvar = initvar+1)
    mem[initvar] = _RAND_0[63:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {2{`RANDOM}};
  read_data_0_r = _RAND_1[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module AXI4RAM(
  input         clock,
  input         reset,
  output        io_in_aw_ready, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input         io_in_aw_valid, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input  [31:0] io_in_aw_bits_addr, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output        io_in_w_ready, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input         io_in_w_valid, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input  [63:0] io_in_w_bits_data, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input         io_in_w_bits_last, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output        io_in_b_valid, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output        io_in_ar_ready, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input         io_in_ar_valid, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input  [31:0] io_in_ar_bits_addr, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input  [7:0]  io_in_ar_bits_len, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input  [2:0]  io_in_ar_bits_size, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input  [1:0]  io_in_ar_bits_burst, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output        io_in_r_valid, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output [63:0] io_in_r_bits_data, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output        io_in_r_bits_last // @[src/main/scala/device/AXI4Slave.scala 28:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [63:0] _RAND_14;
`endif // RANDOMIZE_REG_INIT
  wire  rdata_mem_clock; // @[difftest/src/main/scala/common/Mem.scala 305:31]
  wire  rdata_mem_read_valid; // @[difftest/src/main/scala/common/Mem.scala 305:31]
  wire [63:0] rdata_mem_read_index; // @[difftest/src/main/scala/common/Mem.scala 305:31]
  wire [63:0] rdata_mem_read_data_0; // @[difftest/src/main/scala/common/Mem.scala 305:31]
  wire  rdata_mem_write_valid; // @[difftest/src/main/scala/common/Mem.scala 305:31]
  wire [63:0] rdata_mem_write_index; // @[difftest/src/main/scala/common/Mem.scala 305:31]
  wire [63:0] rdata_mem_write_data_0; // @[difftest/src/main/scala/common/Mem.scala 305:31]
  reg [7:0] c_value; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
  reg [7:0] readBeatCnt; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
  wire  _len_T = io_in_ar_ready & io_in_ar_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  reg [7:0] len_r; // @[src/main/scala/utils/Hold.scala 23:65]
  wire [7:0] _GEN_0 = _len_T ? io_in_ar_bits_len : len_r; // @[src/main/scala/utils/Hold.scala 23:{65,65,65}]
  reg [1:0] burst_r; // @[src/main/scala/utils/Hold.scala 23:65]
  wire [1:0] _GEN_1 = _len_T ? io_in_ar_bits_burst : burst_r; // @[src/main/scala/utils/Hold.scala 23:{65,65,65}]
  wire [31:0] _wrapAddr_WIRE = {{24'd0}, io_in_ar_bits_len}; // @[src/main/scala/device/AXI4Slave.scala 45:{69,69}]
  wire [38:0] _GEN_19 = {{7'd0}, _wrapAddr_WIRE}; // @[src/main/scala/device/AXI4Slave.scala 45:89]
  wire [38:0] _wrapAddr_T = _GEN_19 << io_in_ar_bits_size; // @[src/main/scala/device/AXI4Slave.scala 45:89]
  wire [38:0] _wrapAddr_T_1 = ~_wrapAddr_T; // @[src/main/scala/device/AXI4Slave.scala 45:42]
  wire [38:0] _GEN_28 = {{7'd0}, io_in_ar_bits_addr}; // @[src/main/scala/device/AXI4Slave.scala 45:40]
  wire [38:0] wrapAddr = _GEN_28 & _wrapAddr_T_1; // @[src/main/scala/device/AXI4Slave.scala 45:40]
  reg [38:0] raddr_r; // @[src/main/scala/utils/Hold.scala 23:65]
  wire [38:0] _GEN_2 = _len_T ? wrapAddr : raddr_r; // @[src/main/scala/utils/Hold.scala 23:{65,65,65}]
  wire [7:0] _value_T_1 = readBeatCnt + 8'h1; // @[src/main/scala/chisel3/util/Counter.scala 77:24]
  wire [7:0] _GEN_3 = _GEN_1 == 2'h2 & readBeatCnt == _GEN_0 ? 8'h0 : _value_T_1; // @[src/main/scala/device/AXI4Slave.scala 50:{77,93} src/main/scala/chisel3/util/Counter.scala 77:15]
  reg  ren_REG; // @[src/main/scala/device/AXI4Slave.scala 73:17]
  wire  ren = ren_REG | io_in_r_valid & ~io_in_r_bits_last; // @[src/main/scala/device/AXI4Slave.scala 73:44]
  wire [7:0] _GEN_4 = ren ? _GEN_3 : readBeatCnt; // @[src/main/scala/device/AXI4Slave.scala 48:18 src/main/scala/chisel3/util/Counter.scala 61:40]
  wire [7:0] _value_T_3 = c_value + 8'h1; // @[src/main/scala/chisel3/util/Counter.scala 77:24]
  wire [31:0] _value_T_4 = io_in_ar_bits_addr >> io_in_ar_bits_size; // @[src/main/scala/device/AXI4Slave.scala 57:45]
  wire [31:0] _value_T_5 = _value_T_4 & _wrapAddr_WIRE; // @[src/main/scala/device/AXI4Slave.scala 57:67]
  wire  _T_7 = io_in_ar_bits_len != 8'h0 & io_in_ar_bits_burst == 2'h2; // @[src/main/scala/device/AXI4Slave.scala 58:40]
  wire  _T_11 = io_in_ar_bits_len == 8'h7; // @[src/main/scala/device/AXI4Slave.scala 60:30]
  wire  _T_12 = io_in_ar_bits_len == 8'h1 | io_in_ar_bits_len == 8'h3 | _T_11; // @[src/main/scala/device/AXI4Slave.scala 59:71]
  wire  _T_14 = _T_12 | io_in_ar_bits_len == 8'hf; // @[src/main/scala/device/AXI4Slave.scala 60:38]
  wire [31:0] _GEN_7 = _len_T ? _value_T_5 : {{24'd0}, _GEN_4}; // @[src/main/scala/device/AXI4Slave.scala 56:27 57:23]
  wire  _r_busy_T_2 = io_in_r_valid & io_in_r_bits_last; // @[src/main/scala/device/AXI4Slave.scala 70:52]
  reg  r_busy; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  _GEN_8 = _r_busy_T_2 ? 1'h0 : r_busy; // @[src/main/scala/utils/StopWatch.scala 26:19 24:20 26:23]
  wire  _GEN_9 = _len_T | _GEN_8; // @[src/main/scala/utils/StopWatch.scala 27:{20,24}]
  wire  _io_in_r_valid_T_2 = ren & (_len_T | r_busy); // @[src/main/scala/device/AXI4Slave.scala 74:35]
  reg  io_in_r_valid_r; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  _GEN_10 = io_in_r_valid ? 1'h0 : io_in_r_valid_r; // @[src/main/scala/utils/StopWatch.scala 26:19 24:20 26:23]
  wire  _GEN_11 = _io_in_r_valid_T_2 | _GEN_10; // @[src/main/scala/utils/StopWatch.scala 27:{20,24}]
  reg [7:0] writeBeatCnt; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
  wire  _waddr_T = io_in_aw_ready & io_in_aw_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  reg [31:0] waddr_r; // @[src/main/scala/utils/Hold.scala 23:65]
  wire [31:0] _GEN_12 = _waddr_T ? io_in_aw_bits_addr : waddr_r; // @[src/main/scala/utils/Hold.scala 23:{65,65,65}]
  wire  _T_18 = io_in_w_ready & io_in_w_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  wire [7:0] _value_T_7 = writeBeatCnt + 8'h1; // @[src/main/scala/chisel3/util/Counter.scala 77:24]
  reg  w_busy; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  _GEN_15 = io_in_b_valid ? 1'h0 : w_busy; // @[src/main/scala/utils/StopWatch.scala 26:19 24:20 26:23]
  wire  _GEN_16 = _waddr_T | _GEN_15; // @[src/main/scala/utils/StopWatch.scala 27:{20,24}]
  wire  _io_in_b_valid_T_1 = _T_18 & io_in_w_bits_last; // @[src/main/scala/device/AXI4Slave.scala 97:41]
  reg  io_in_b_valid_r; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  _GEN_17 = io_in_b_valid ? 1'h0 : io_in_b_valid_r; // @[src/main/scala/utils/StopWatch.scala 26:19 24:20 26:23]
  wire  _GEN_18 = _io_in_b_valid_T_1 | _GEN_17; // @[src/main/scala/utils/StopWatch.scala 27:{20,24}]
  wire [31:0] _wIdx_T = _GEN_12 & 32'h7ffffff; // @[src/main/scala/device/AXI4RAM.scala 33:33]
  wire [28:0] _GEN_30 = {{21'd0}, writeBeatCnt}; // @[src/main/scala/device/AXI4RAM.scala 36:27]
  wire [28:0] wIdx = _wIdx_T[31:3] + _GEN_30; // @[src/main/scala/device/AXI4RAM.scala 36:27]
  wire [38:0] _rIdx_T = _GEN_2 & 39'h7ffffff; // @[src/main/scala/device/AXI4RAM.scala 33:33]
  wire [35:0] _GEN_31 = {{28'd0}, readBeatCnt}; // @[src/main/scala/device/AXI4RAM.scala 37:27]
  wire [35:0] rIdx = _rIdx_T[38:3] + _GEN_31; // @[src/main/scala/device/AXI4RAM.scala 37:27]
  wire  _wen_T_1 = wIdx < 29'h1000000; // @[src/main/scala/device/AXI4RAM.scala 34:32]
  wire [31:0] rdata_lo = {io_in_w_bits_data[31:24],io_in_w_bits_data[23:16],io_in_w_bits_data[15:8],io_in_w_bits_data[7:
    0]}; // @[difftest/src/main/scala/common/Mem.scala 187:42]
  wire [31:0] rdata_hi = {io_in_w_bits_data[63:56],io_in_w_bits_data[55:48],io_in_w_bits_data[47:40],io_in_w_bits_data[
    39:32]}; // @[difftest/src/main/scala/common/Mem.scala 187:42]
  reg  rdata_REG; // @[difftest/src/main/scala/common/Mem.scala 181:16]
  reg  rdata_REG_1; // @[difftest/src/main/scala/common/Mem.scala 181:61]
  reg [63:0] rdata_r_0; // @[difftest/src/main/scala/common/Mem.scala 181:42]
  wire [63:0] _rdata_T_36_0 = rdata_REG ? rdata_mem_read_data_0 : rdata_r_0; // @[difftest/src/main/scala/common/Mem.scala 181:8]
  wire [31:0] rdata_lo_2 = {_rdata_T_36_0[31:24],_rdata_T_36_0[23:16],_rdata_T_36_0[15:8],_rdata_T_36_0[7:0]}; // @[src/main/scala/device/AXI4RAM.scala 49:32]
  wire [31:0] rdata_hi_2 = {_rdata_T_36_0[63:56],_rdata_T_36_0[55:48],_rdata_T_36_0[47:40],_rdata_T_36_0[39:32]}; // @[src/main/scala/device/AXI4RAM.scala 49:32]
  wire [31:0] _GEN_32 = reset ? 32'h0 : _GEN_7; // @[src/main/scala/chisel3/util/Counter.scala 61:{40,40}]
  SynthesizableDifftestMem rdata_mem ( // @[difftest/src/main/scala/common/Mem.scala 305:31]
    .clock(rdata_mem_clock),
    .read_valid(rdata_mem_read_valid),
    .read_index(rdata_mem_read_index),
    .read_data_0(rdata_mem_read_data_0),
    .write_valid(rdata_mem_write_valid),
    .write_index(rdata_mem_write_index),
    .write_data_0(rdata_mem_write_data_0)
  );
  assign io_in_aw_ready = ~w_busy; // @[src/main/scala/device/AXI4Slave.scala 94:18]
  assign io_in_w_ready = io_in_aw_valid | w_busy; // @[src/main/scala/device/AXI4Slave.scala 95:30]
  assign io_in_b_valid = io_in_b_valid_r; // @[src/main/scala/device/AXI4Slave.scala 97:14]
  assign io_in_ar_ready = 1'h1; // @[src/main/scala/device/AXI4Slave.scala 71:29]
  assign io_in_r_valid = io_in_r_valid_r; // @[src/main/scala/device/AXI4Slave.scala 74:14]
  assign io_in_r_bits_data = {rdata_hi_2,rdata_lo_2}; // @[src/main/scala/device/AXI4RAM.scala 49:32]
  assign io_in_r_bits_last = c_value == _GEN_0; // @[src/main/scala/device/AXI4Slave.scala 47:36]
  assign rdata_mem_clock = clock;
  assign rdata_mem_read_valid = ren_REG | io_in_r_valid & ~io_in_r_bits_last; // @[src/main/scala/device/AXI4Slave.scala 73:44]
  assign rdata_mem_read_index = {{28'd0}, rIdx}; // @[difftest/src/main/scala/common/Mem.scala 180:16]
  assign rdata_mem_write_valid = _T_18 & _wen_T_1; // @[src/main/scala/device/AXI4RAM.scala 38:23]
  assign rdata_mem_write_index = {{35'd0}, wIdx};
  assign rdata_mem_write_data_0 = {rdata_hi,rdata_lo}; // @[difftest/src/main/scala/common/Mem.scala 187:42]
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/chisel3/util/Counter.scala 61:40]
      c_value <= 8'h0; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end else if (io_in_r_valid) begin // @[src/main/scala/device/AXI4Slave.scala 52:26]
      if (io_in_r_bits_last) begin // @[src/main/scala/device/AXI4Slave.scala 54:33]
        c_value <= 8'h0; // @[src/main/scala/device/AXI4Slave.scala 54:43]
      end else begin
        c_value <= _value_T_3; // @[src/main/scala/chisel3/util/Counter.scala 77:15]
      end
    end
    readBeatCnt <= _GEN_32[7:0]; // @[src/main/scala/chisel3/util/Counter.scala 61:{40,40}]
    if (reset) begin // @[src/main/scala/utils/Hold.scala 23:65]
      len_r <= 8'h0; // @[src/main/scala/utils/Hold.scala 23:65]
    end else if (_len_T) begin // @[src/main/scala/utils/Hold.scala 23:65]
      len_r <= io_in_ar_bits_len; // @[src/main/scala/utils/Hold.scala 23:65]
    end
    if (reset) begin // @[src/main/scala/utils/Hold.scala 23:65]
      burst_r <= 2'h0; // @[src/main/scala/utils/Hold.scala 23:65]
    end else if (_len_T) begin // @[src/main/scala/utils/Hold.scala 23:65]
      burst_r <= io_in_ar_bits_burst; // @[src/main/scala/utils/Hold.scala 23:65]
    end
    if (reset) begin // @[src/main/scala/utils/Hold.scala 23:65]
      raddr_r <= 39'h0; // @[src/main/scala/utils/Hold.scala 23:65]
    end else if (_len_T) begin // @[src/main/scala/utils/Hold.scala 23:65]
      raddr_r <= wrapAddr; // @[src/main/scala/utils/Hold.scala 23:65]
    end
    if (reset) begin // @[src/main/scala/device/AXI4Slave.scala 73:17]
      ren_REG <= 1'h0; // @[src/main/scala/device/AXI4Slave.scala 73:17]
    end else begin
      ren_REG <= _len_T; // @[src/main/scala/device/AXI4Slave.scala 73:17]
    end
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      r_busy <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else begin
      r_busy <= _GEN_9;
    end
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      io_in_r_valid_r <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else begin
      io_in_r_valid_r <= _GEN_11;
    end
    if (reset) begin // @[src/main/scala/chisel3/util/Counter.scala 61:40]
      writeBeatCnt <= 8'h0; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end else if (_T_18) begin // @[src/main/scala/device/AXI4Slave.scala 82:26]
      if (io_in_w_bits_last) begin // @[src/main/scala/device/AXI4Slave.scala 84:33]
        writeBeatCnt <= 8'h0; // @[src/main/scala/device/AXI4Slave.scala 84:43]
      end else begin
        writeBeatCnt <= _value_T_7; // @[src/main/scala/chisel3/util/Counter.scala 77:15]
      end
    end
    if (reset) begin // @[src/main/scala/utils/Hold.scala 23:65]
      waddr_r <= 32'h0; // @[src/main/scala/utils/Hold.scala 23:65]
    end else if (_waddr_T) begin // @[src/main/scala/utils/Hold.scala 23:65]
      waddr_r <= io_in_aw_bits_addr; // @[src/main/scala/utils/Hold.scala 23:65]
    end
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      w_busy <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else begin
      w_busy <= _GEN_16;
    end
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      io_in_b_valid_r <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else begin
      io_in_b_valid_r <= _GEN_18;
    end
    rdata_REG <= ren_REG | io_in_r_valid & ~io_in_r_bits_last; // @[src/main/scala/device/AXI4Slave.scala 73:44]
    rdata_REG_1 <= ren_REG | io_in_r_valid & ~io_in_r_bits_last; // @[src/main/scala/device/AXI4Slave.scala 73:44]
    if (rdata_REG_1) begin // @[difftest/src/main/scala/common/Mem.scala 181:42]
      rdata_r_0 <= rdata_mem_read_data_0; // @[difftest/src/main/scala/common/Mem.scala 181:42]
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_len_T & _T_7 & ~reset & ~_T_14) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at AXI4Slave.scala:59 assert(axi4.ar.bits.len === 1.U || axi4.ar.bits.len === 3.U ||\n"
            ); // @[src/main/scala/device/AXI4Slave.scala 59:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~_T_14 & (_len_T & _T_7 & ~reset)) begin
          $fatal; // @[src/main/scala/device/AXI4Slave.scala 59:17]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  c_value = _RAND_0[7:0];
  _RAND_1 = {1{`RANDOM}};
  readBeatCnt = _RAND_1[7:0];
  _RAND_2 = {1{`RANDOM}};
  len_r = _RAND_2[7:0];
  _RAND_3 = {1{`RANDOM}};
  burst_r = _RAND_3[1:0];
  _RAND_4 = {2{`RANDOM}};
  raddr_r = _RAND_4[38:0];
  _RAND_5 = {1{`RANDOM}};
  ren_REG = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  r_busy = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  io_in_r_valid_r = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  writeBeatCnt = _RAND_8[7:0];
  _RAND_9 = {1{`RANDOM}};
  waddr_r = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  w_busy = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  io_in_b_valid_r = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  rdata_REG = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  rdata_REG_1 = _RAND_13[0:0];
  _RAND_14 = {2{`RANDOM}};
  rdata_r_0 = _RAND_14[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module LatencyPipe(
  output        io_in_ready, // @[src/main/scala/utils/LatencyPipe.scala 9:14]
  input         io_in_valid, // @[src/main/scala/utils/LatencyPipe.scala 9:14]
  input  [31:0] io_in_bits_addr, // @[src/main/scala/utils/LatencyPipe.scala 9:14]
  input  [7:0]  io_in_bits_len, // @[src/main/scala/utils/LatencyPipe.scala 9:14]
  input  [2:0]  io_in_bits_size, // @[src/main/scala/utils/LatencyPipe.scala 9:14]
  input  [1:0]  io_in_bits_burst, // @[src/main/scala/utils/LatencyPipe.scala 9:14]
  input         io_out_ready, // @[src/main/scala/utils/LatencyPipe.scala 9:14]
  output        io_out_valid, // @[src/main/scala/utils/LatencyPipe.scala 9:14]
  output [31:0] io_out_bits_addr, // @[src/main/scala/utils/LatencyPipe.scala 9:14]
  output [7:0]  io_out_bits_len, // @[src/main/scala/utils/LatencyPipe.scala 9:14]
  output [2:0]  io_out_bits_size, // @[src/main/scala/utils/LatencyPipe.scala 9:14]
  output [1:0]  io_out_bits_burst // @[src/main/scala/utils/LatencyPipe.scala 9:14]
);
  assign io_in_ready = io_out_ready; // @[src/main/scala/utils/LatencyPipe.scala 17:10]
  assign io_out_valid = io_in_valid; // @[src/main/scala/utils/LatencyPipe.scala 17:10]
  assign io_out_bits_addr = io_in_bits_addr; // @[src/main/scala/utils/LatencyPipe.scala 17:10]
  assign io_out_bits_len = io_in_bits_len; // @[src/main/scala/utils/LatencyPipe.scala 17:10]
  assign io_out_bits_size = io_in_bits_size; // @[src/main/scala/utils/LatencyPipe.scala 17:10]
  assign io_out_bits_burst = io_in_bits_burst; // @[src/main/scala/utils/LatencyPipe.scala 17:10]
endmodule
module AXI4Delayer(
  output        io_in_aw_ready, // @[src/main/scala/bus/axi4/Delayer.scala 10:14]
  input         io_in_aw_valid, // @[src/main/scala/bus/axi4/Delayer.scala 10:14]
  input  [31:0] io_in_aw_bits_addr, // @[src/main/scala/bus/axi4/Delayer.scala 10:14]
  input  [7:0]  io_in_aw_bits_len, // @[src/main/scala/bus/axi4/Delayer.scala 10:14]
  input  [2:0]  io_in_aw_bits_size, // @[src/main/scala/bus/axi4/Delayer.scala 10:14]
  input  [1:0]  io_in_aw_bits_burst, // @[src/main/scala/bus/axi4/Delayer.scala 10:14]
  output        io_in_w_ready, // @[src/main/scala/bus/axi4/Delayer.scala 10:14]
  input         io_in_w_valid, // @[src/main/scala/bus/axi4/Delayer.scala 10:14]
  input  [63:0] io_in_w_bits_data, // @[src/main/scala/bus/axi4/Delayer.scala 10:14]
  input         io_in_w_bits_last, // @[src/main/scala/bus/axi4/Delayer.scala 10:14]
  output        io_in_b_valid, // @[src/main/scala/bus/axi4/Delayer.scala 10:14]
  output        io_in_ar_ready, // @[src/main/scala/bus/axi4/Delayer.scala 10:14]
  input         io_in_ar_valid, // @[src/main/scala/bus/axi4/Delayer.scala 10:14]
  input  [31:0] io_in_ar_bits_addr, // @[src/main/scala/bus/axi4/Delayer.scala 10:14]
  input  [7:0]  io_in_ar_bits_len, // @[src/main/scala/bus/axi4/Delayer.scala 10:14]
  output        io_in_r_valid, // @[src/main/scala/bus/axi4/Delayer.scala 10:14]
  output [63:0] io_in_r_bits_data, // @[src/main/scala/bus/axi4/Delayer.scala 10:14]
  output        io_in_r_bits_last, // @[src/main/scala/bus/axi4/Delayer.scala 10:14]
  input         io_out_aw_ready, // @[src/main/scala/bus/axi4/Delayer.scala 10:14]
  output        io_out_aw_valid, // @[src/main/scala/bus/axi4/Delayer.scala 10:14]
  output [31:0] io_out_aw_bits_addr, // @[src/main/scala/bus/axi4/Delayer.scala 10:14]
  input         io_out_w_ready, // @[src/main/scala/bus/axi4/Delayer.scala 10:14]
  output        io_out_w_valid, // @[src/main/scala/bus/axi4/Delayer.scala 10:14]
  output [63:0] io_out_w_bits_data, // @[src/main/scala/bus/axi4/Delayer.scala 10:14]
  output        io_out_w_bits_last, // @[src/main/scala/bus/axi4/Delayer.scala 10:14]
  input         io_out_b_valid, // @[src/main/scala/bus/axi4/Delayer.scala 10:14]
  output        io_out_ar_valid, // @[src/main/scala/bus/axi4/Delayer.scala 10:14]
  output [31:0] io_out_ar_bits_addr, // @[src/main/scala/bus/axi4/Delayer.scala 10:14]
  output [7:0]  io_out_ar_bits_len, // @[src/main/scala/bus/axi4/Delayer.scala 10:14]
  output [2:0]  io_out_ar_bits_size, // @[src/main/scala/bus/axi4/Delayer.scala 10:14]
  output [1:0]  io_out_ar_bits_burst, // @[src/main/scala/bus/axi4/Delayer.scala 10:14]
  input         io_out_r_valid, // @[src/main/scala/bus/axi4/Delayer.scala 10:14]
  input  [63:0] io_out_r_bits_data, // @[src/main/scala/bus/axi4/Delayer.scala 10:14]
  input         io_out_r_bits_last // @[src/main/scala/bus/axi4/Delayer.scala 10:14]
);
  wire  io_out_ar_pipe_io_in_ready; // @[src/main/scala/utils/LatencyPipe.scala 22:22]
  wire  io_out_ar_pipe_io_in_valid; // @[src/main/scala/utils/LatencyPipe.scala 22:22]
  wire [31:0] io_out_ar_pipe_io_in_bits_addr; // @[src/main/scala/utils/LatencyPipe.scala 22:22]
  wire [7:0] io_out_ar_pipe_io_in_bits_len; // @[src/main/scala/utils/LatencyPipe.scala 22:22]
  wire [2:0] io_out_ar_pipe_io_in_bits_size; // @[src/main/scala/utils/LatencyPipe.scala 22:22]
  wire [1:0] io_out_ar_pipe_io_in_bits_burst; // @[src/main/scala/utils/LatencyPipe.scala 22:22]
  wire  io_out_ar_pipe_io_out_ready; // @[src/main/scala/utils/LatencyPipe.scala 22:22]
  wire  io_out_ar_pipe_io_out_valid; // @[src/main/scala/utils/LatencyPipe.scala 22:22]
  wire [31:0] io_out_ar_pipe_io_out_bits_addr; // @[src/main/scala/utils/LatencyPipe.scala 22:22]
  wire [7:0] io_out_ar_pipe_io_out_bits_len; // @[src/main/scala/utils/LatencyPipe.scala 22:22]
  wire [2:0] io_out_ar_pipe_io_out_bits_size; // @[src/main/scala/utils/LatencyPipe.scala 22:22]
  wire [1:0] io_out_ar_pipe_io_out_bits_burst; // @[src/main/scala/utils/LatencyPipe.scala 22:22]
  wire  io_out_aw_pipe_io_in_ready; // @[src/main/scala/utils/LatencyPipe.scala 22:22]
  wire  io_out_aw_pipe_io_in_valid; // @[src/main/scala/utils/LatencyPipe.scala 22:22]
  wire [31:0] io_out_aw_pipe_io_in_bits_addr; // @[src/main/scala/utils/LatencyPipe.scala 22:22]
  wire [7:0] io_out_aw_pipe_io_in_bits_len; // @[src/main/scala/utils/LatencyPipe.scala 22:22]
  wire [2:0] io_out_aw_pipe_io_in_bits_size; // @[src/main/scala/utils/LatencyPipe.scala 22:22]
  wire [1:0] io_out_aw_pipe_io_in_bits_burst; // @[src/main/scala/utils/LatencyPipe.scala 22:22]
  wire  io_out_aw_pipe_io_out_ready; // @[src/main/scala/utils/LatencyPipe.scala 22:22]
  wire  io_out_aw_pipe_io_out_valid; // @[src/main/scala/utils/LatencyPipe.scala 22:22]
  wire [31:0] io_out_aw_pipe_io_out_bits_addr; // @[src/main/scala/utils/LatencyPipe.scala 22:22]
  wire [7:0] io_out_aw_pipe_io_out_bits_len; // @[src/main/scala/utils/LatencyPipe.scala 22:22]
  wire [2:0] io_out_aw_pipe_io_out_bits_size; // @[src/main/scala/utils/LatencyPipe.scala 22:22]
  wire [1:0] io_out_aw_pipe_io_out_bits_burst; // @[src/main/scala/utils/LatencyPipe.scala 22:22]
  LatencyPipe io_out_ar_pipe ( // @[src/main/scala/utils/LatencyPipe.scala 22:22]
    .io_in_ready(io_out_ar_pipe_io_in_ready),
    .io_in_valid(io_out_ar_pipe_io_in_valid),
    .io_in_bits_addr(io_out_ar_pipe_io_in_bits_addr),
    .io_in_bits_len(io_out_ar_pipe_io_in_bits_len),
    .io_in_bits_size(io_out_ar_pipe_io_in_bits_size),
    .io_in_bits_burst(io_out_ar_pipe_io_in_bits_burst),
    .io_out_ready(io_out_ar_pipe_io_out_ready),
    .io_out_valid(io_out_ar_pipe_io_out_valid),
    .io_out_bits_addr(io_out_ar_pipe_io_out_bits_addr),
    .io_out_bits_len(io_out_ar_pipe_io_out_bits_len),
    .io_out_bits_size(io_out_ar_pipe_io_out_bits_size),
    .io_out_bits_burst(io_out_ar_pipe_io_out_bits_burst)
  );
  LatencyPipe io_out_aw_pipe ( // @[src/main/scala/utils/LatencyPipe.scala 22:22]
    .io_in_ready(io_out_aw_pipe_io_in_ready),
    .io_in_valid(io_out_aw_pipe_io_in_valid),
    .io_in_bits_addr(io_out_aw_pipe_io_in_bits_addr),
    .io_in_bits_len(io_out_aw_pipe_io_in_bits_len),
    .io_in_bits_size(io_out_aw_pipe_io_in_bits_size),
    .io_in_bits_burst(io_out_aw_pipe_io_in_bits_burst),
    .io_out_ready(io_out_aw_pipe_io_out_ready),
    .io_out_valid(io_out_aw_pipe_io_out_valid),
    .io_out_bits_addr(io_out_aw_pipe_io_out_bits_addr),
    .io_out_bits_len(io_out_aw_pipe_io_out_bits_len),
    .io_out_bits_size(io_out_aw_pipe_io_out_bits_size),
    .io_out_bits_burst(io_out_aw_pipe_io_out_bits_burst)
  );
  assign io_in_aw_ready = io_out_aw_pipe_io_in_ready; // @[src/main/scala/utils/LatencyPipe.scala 23:16]
  assign io_in_w_ready = io_out_w_ready; // @[src/main/scala/bus/axi4/Delayer.scala 17:13]
  assign io_in_b_valid = io_out_b_valid; // @[src/main/scala/bus/axi4/Delayer.scala 18:13]
  assign io_in_ar_ready = io_out_ar_pipe_io_in_ready; // @[src/main/scala/utils/LatencyPipe.scala 23:16]
  assign io_in_r_valid = io_out_r_valid; // @[src/main/scala/bus/axi4/Delayer.scala 19:13]
  assign io_in_r_bits_data = io_out_r_bits_data; // @[src/main/scala/bus/axi4/Delayer.scala 19:13]
  assign io_in_r_bits_last = io_out_r_bits_last; // @[src/main/scala/bus/axi4/Delayer.scala 19:13]
  assign io_out_aw_valid = io_out_aw_pipe_io_out_valid; // @[src/main/scala/bus/axi4/Delayer.scala 16:13]
  assign io_out_aw_bits_addr = io_out_aw_pipe_io_out_bits_addr; // @[src/main/scala/bus/axi4/Delayer.scala 16:13]
  assign io_out_w_valid = io_in_w_valid; // @[src/main/scala/bus/axi4/Delayer.scala 17:13]
  assign io_out_w_bits_data = io_in_w_bits_data; // @[src/main/scala/bus/axi4/Delayer.scala 17:13]
  assign io_out_w_bits_last = io_in_w_bits_last; // @[src/main/scala/bus/axi4/Delayer.scala 17:13]
  assign io_out_ar_valid = io_out_ar_pipe_io_out_valid; // @[src/main/scala/bus/axi4/Delayer.scala 15:13]
  assign io_out_ar_bits_addr = io_out_ar_pipe_io_out_bits_addr; // @[src/main/scala/bus/axi4/Delayer.scala 15:13]
  assign io_out_ar_bits_len = io_out_ar_pipe_io_out_bits_len; // @[src/main/scala/bus/axi4/Delayer.scala 15:13]
  assign io_out_ar_bits_size = io_out_ar_pipe_io_out_bits_size; // @[src/main/scala/bus/axi4/Delayer.scala 15:13]
  assign io_out_ar_bits_burst = io_out_ar_pipe_io_out_bits_burst; // @[src/main/scala/bus/axi4/Delayer.scala 15:13]
  assign io_out_ar_pipe_io_in_valid = io_in_ar_valid; // @[src/main/scala/utils/LatencyPipe.scala 23:16]
  assign io_out_ar_pipe_io_in_bits_addr = io_in_ar_bits_addr; // @[src/main/scala/utils/LatencyPipe.scala 23:16]
  assign io_out_ar_pipe_io_in_bits_len = io_in_ar_bits_len; // @[src/main/scala/utils/LatencyPipe.scala 23:16]
  assign io_out_ar_pipe_io_in_bits_size = 3'h3; // @[src/main/scala/utils/LatencyPipe.scala 23:16]
  assign io_out_ar_pipe_io_in_bits_burst = 2'h2; // @[src/main/scala/utils/LatencyPipe.scala 23:16]
  assign io_out_ar_pipe_io_out_ready = 1'h1; // @[src/main/scala/bus/axi4/Delayer.scala 15:13]
  assign io_out_aw_pipe_io_in_valid = io_in_aw_valid; // @[src/main/scala/utils/LatencyPipe.scala 23:16]
  assign io_out_aw_pipe_io_in_bits_addr = io_in_aw_bits_addr; // @[src/main/scala/utils/LatencyPipe.scala 23:16]
  assign io_out_aw_pipe_io_in_bits_len = io_in_aw_bits_len; // @[src/main/scala/utils/LatencyPipe.scala 23:16]
  assign io_out_aw_pipe_io_in_bits_size = io_in_aw_bits_size; // @[src/main/scala/utils/LatencyPipe.scala 23:16]
  assign io_out_aw_pipe_io_in_bits_burst = io_in_aw_bits_burst; // @[src/main/scala/utils/LatencyPipe.scala 23:16]
  assign io_out_aw_pipe_io_out_ready = io_out_aw_ready; // @[src/main/scala/bus/axi4/Delayer.scala 16:13]
endmodule
module SimpleBusCrossbar1toN_1(
  input         clock,
  input         reset,
  output        io_in_req_ready, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  input         io_in_req_valid, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  input  [31:0] io_in_req_bits_addr, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  input  [2:0]  io_in_req_bits_size, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  input  [3:0]  io_in_req_bits_cmd, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  input  [7:0]  io_in_req_bits_wmask, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  input  [63:0] io_in_req_bits_wdata, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  input         io_in_resp_ready, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output        io_in_resp_valid, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output [3:0]  io_in_resp_bits_cmd, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output [63:0] io_in_resp_bits_rdata, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  input         io_out_0_req_ready, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output        io_out_0_req_valid, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output [31:0] io_out_0_req_bits_addr, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output [3:0]  io_out_0_req_bits_cmd, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output [7:0]  io_out_0_req_bits_wmask, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output [63:0] io_out_0_req_bits_wdata, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output        io_out_0_resp_ready, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  input         io_out_0_resp_valid, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  input  [63:0] io_out_0_resp_bits_rdata, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  input         io_out_1_req_ready, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output        io_out_1_req_valid, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output [31:0] io_out_1_req_bits_addr, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output [3:0]  io_out_1_req_bits_cmd, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output [7:0]  io_out_1_req_bits_wmask, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output [63:0] io_out_1_req_bits_wdata, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output        io_out_1_resp_ready, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  input         io_out_1_resp_valid, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  input  [63:0] io_out_1_resp_bits_rdata, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  input         io_out_2_req_ready, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output        io_out_2_req_valid, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output [31:0] io_out_2_req_bits_addr, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output [3:0]  io_out_2_req_bits_cmd, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output [7:0]  io_out_2_req_bits_wmask, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output [63:0] io_out_2_req_bits_wdata, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output        io_out_2_resp_ready, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  input         io_out_2_resp_valid, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  input  [63:0] io_out_2_resp_bits_rdata, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  input         io_out_3_req_ready, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output        io_out_3_req_valid, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output [31:0] io_out_3_req_bits_addr, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output [3:0]  io_out_3_req_bits_cmd, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output [7:0]  io_out_3_req_bits_wmask, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output [63:0] io_out_3_req_bits_wdata, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output        io_out_3_resp_ready, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  input         io_out_3_resp_valid, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  input  [63:0] io_out_3_resp_bits_rdata, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  input         DISPLAY_ENABLE
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
`endif // RANDOMIZE_REG_INIT
  reg [1:0] state; // @[src/main/scala/bus/simplebus/Crossbar.scala 32:22]
  wire  outMatchVec_0 = io_in_req_bits_addr >= 32'h40600000 & io_in_req_bits_addr < 32'h40600010; // @[src/main/scala/bus/simplebus/Crossbar.scala 37:34]
  wire  outMatchVec_1 = io_in_req_bits_addr >= 32'h40000000 & io_in_req_bits_addr < 32'h40001000; // @[src/main/scala/bus/simplebus/Crossbar.scala 37:34]
  wire  outMatchVec_2 = io_in_req_bits_addr >= 32'h40004000 & io_in_req_bits_addr < 32'h40005000; // @[src/main/scala/bus/simplebus/Crossbar.scala 37:34]
  wire  outMatchVec_3 = io_in_req_bits_addr >= 32'h40003000 & io_in_req_bits_addr < 32'h40004000; // @[src/main/scala/bus/simplebus/Crossbar.scala 37:34]
  wire [3:0] _outSelVec_enc_T = outMatchVec_3 ? 4'h8 : 4'h0; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [3:0] _outSelVec_enc_T_1 = outMatchVec_2 ? 4'h4 : _outSelVec_enc_T; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [3:0] _outSelVec_enc_T_2 = outMatchVec_1 ? 4'h2 : _outSelVec_enc_T_1; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [3:0] outSelVec_enc = outMatchVec_0 ? 4'h1 : _outSelVec_enc_T_2; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire  outSelVec_0 = outSelVec_enc[0]; // @[src/main/scala/chisel3/util/OneHot.scala 83:30]
  wire  outSelVec_1 = outSelVec_enc[1]; // @[src/main/scala/chisel3/util/OneHot.scala 83:30]
  wire  outSelVec_2 = outSelVec_enc[2]; // @[src/main/scala/chisel3/util/OneHot.scala 83:30]
  wire  outSelVec_3 = outSelVec_enc[3]; // @[src/main/scala/chisel3/util/OneHot.scala 83:30]
  wire  _outSelRespVec_T = io_in_req_ready & io_in_req_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  wire  _outSelRespVec_T_1 = state == 2'h0; // @[src/main/scala/bus/simplebus/Crossbar.scala 41:57]
  wire  _outSelRespVec_T_2 = _outSelRespVec_T & state == 2'h0; // @[src/main/scala/bus/simplebus/Crossbar.scala 41:48]
  reg  outSelRespVec_0; // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
  reg  outSelRespVec_1; // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
  reg  outSelRespVec_2; // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
  reg  outSelRespVec_3; // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
  wire [3:0] _reqInvalidAddr_T = {outSelVec_3,outSelVec_2,outSelVec_1,outSelVec_0}; // @[src/main/scala/bus/simplebus/Crossbar.scala 42:54]
  wire  reqInvalidAddr = io_in_req_valid & ~(|_reqInvalidAddr_T); // @[src/main/scala/bus/simplebus/Crossbar.scala 42:40]
  reg [63:0] c; // @[src/main/scala/utils/GTimer.scala 24:20]
  wire [63:0] _c_T_1 = c + 64'h1; // @[src/main/scala/utils/GTimer.scala 25:12]
  wire  _T_2 = ~reset; // @[src/main/scala/bus/simplebus/Crossbar.scala 46:13]
  wire  _T_10 = io_in_resp_ready & io_in_resp_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  wire [1:0] _GEN_6 = _T_10 ? 2'h0 : state; // @[src/main/scala/bus/simplebus/Crossbar.scala 32:22 56:{42,50}]
  wire  _io_in_req_ready_T_6 = outSelVec_0 & io_out_0_req_ready | outSelVec_1 & io_out_1_req_ready | outSelVec_2 &
    io_out_2_req_ready | outSelVec_3 & io_out_3_req_ready; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _io_in_resp_valid_T_6 = outSelRespVec_0 & io_out_0_resp_valid | outSelRespVec_1 & io_out_1_resp_valid |
    outSelRespVec_2 & io_out_2_resp_valid | outSelRespVec_3 & io_out_3_resp_valid; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_in_resp_bits_T = outSelRespVec_0 ? io_out_0_resp_bits_rdata : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_in_resp_bits_T_1 = outSelRespVec_1 ? io_out_1_resp_bits_rdata : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_in_resp_bits_T_2 = outSelRespVec_2 ? io_out_2_resp_bits_rdata : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_in_resp_bits_T_3 = outSelRespVec_3 ? io_out_3_resp_bits_rdata : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_in_resp_bits_T_4 = _io_in_resp_bits_T | _io_in_resp_bits_T_1; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_in_resp_bits_T_5 = _io_in_resp_bits_T_4 | _io_in_resp_bits_T_2; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [3:0] _io_in_resp_bits_T_7 = outSelRespVec_0 ? 4'h6 : 4'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [3:0] _io_in_resp_bits_T_8 = outSelRespVec_1 ? 4'h6 : 4'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [3:0] _io_in_resp_bits_T_9 = outSelRespVec_2 ? 4'h6 : 4'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [3:0] _io_in_resp_bits_T_10 = outSelRespVec_3 ? 4'h6 : 4'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [3:0] _io_in_resp_bits_T_11 = _io_in_resp_bits_T_7 | _io_in_resp_bits_T_8; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [3:0] _io_in_resp_bits_T_12 = _io_in_resp_bits_T_11 | _io_in_resp_bits_T_9; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  reg [63:0] c_1; // @[src/main/scala/utils/GTimer.scala 24:20]
  wire [63:0] _c_T_3 = c_1 + 64'h1; // @[src/main/scala/utils/GTimer.scala 25:12]
  reg [63:0] c_2; // @[src/main/scala/utils/GTimer.scala 24:20]
  wire [63:0] _c_T_5 = c_2 + 64'h1; // @[src/main/scala/utils/GTimer.scala 25:12]
  assign io_in_req_ready = _io_in_req_ready_T_6 | reqInvalidAddr; // @[src/main/scala/bus/simplebus/Crossbar.scala 61:64]
  assign io_in_resp_valid = _io_in_resp_valid_T_6 | state == 2'h2; // @[src/main/scala/bus/simplebus/Crossbar.scala 71:70]
  assign io_in_resp_bits_cmd = _io_in_resp_bits_T_12 | _io_in_resp_bits_T_10; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign io_in_resp_bits_rdata = _io_in_resp_bits_T_5 | _io_in_resp_bits_T_3; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign io_out_0_req_valid = outSelVec_0 & io_in_req_valid & _outSelRespVec_T_1; // @[src/main/scala/bus/simplebus/Crossbar.scala 63:60]
  assign io_out_0_req_bits_addr = io_in_req_bits_addr; // @[src/main/scala/bus/simplebus/Crossbar.scala 64:24]
  assign io_out_0_req_bits_cmd = io_in_req_bits_cmd; // @[src/main/scala/bus/simplebus/Crossbar.scala 64:24]
  assign io_out_0_req_bits_wmask = io_in_req_bits_wmask; // @[src/main/scala/bus/simplebus/Crossbar.scala 64:24]
  assign io_out_0_req_bits_wdata = io_in_req_bits_wdata; // @[src/main/scala/bus/simplebus/Crossbar.scala 64:24]
  assign io_out_0_resp_ready = outSelRespVec_0 & io_in_resp_ready & state == 2'h1; // @[src/main/scala/bus/simplebus/Crossbar.scala 69:66]
  assign io_out_1_req_valid = outSelVec_1 & io_in_req_valid & _outSelRespVec_T_1; // @[src/main/scala/bus/simplebus/Crossbar.scala 63:60]
  assign io_out_1_req_bits_addr = io_in_req_bits_addr; // @[src/main/scala/bus/simplebus/Crossbar.scala 64:24]
  assign io_out_1_req_bits_cmd = io_in_req_bits_cmd; // @[src/main/scala/bus/simplebus/Crossbar.scala 64:24]
  assign io_out_1_req_bits_wmask = io_in_req_bits_wmask; // @[src/main/scala/bus/simplebus/Crossbar.scala 64:24]
  assign io_out_1_req_bits_wdata = io_in_req_bits_wdata; // @[src/main/scala/bus/simplebus/Crossbar.scala 64:24]
  assign io_out_1_resp_ready = outSelRespVec_1 & io_in_resp_ready & state == 2'h1; // @[src/main/scala/bus/simplebus/Crossbar.scala 69:66]
  assign io_out_2_req_valid = outSelVec_2 & io_in_req_valid & _outSelRespVec_T_1; // @[src/main/scala/bus/simplebus/Crossbar.scala 63:60]
  assign io_out_2_req_bits_addr = io_in_req_bits_addr; // @[src/main/scala/bus/simplebus/Crossbar.scala 64:24]
  assign io_out_2_req_bits_cmd = io_in_req_bits_cmd; // @[src/main/scala/bus/simplebus/Crossbar.scala 64:24]
  assign io_out_2_req_bits_wmask = io_in_req_bits_wmask; // @[src/main/scala/bus/simplebus/Crossbar.scala 64:24]
  assign io_out_2_req_bits_wdata = io_in_req_bits_wdata; // @[src/main/scala/bus/simplebus/Crossbar.scala 64:24]
  assign io_out_2_resp_ready = outSelRespVec_2 & io_in_resp_ready & state == 2'h1; // @[src/main/scala/bus/simplebus/Crossbar.scala 69:66]
  assign io_out_3_req_valid = outSelVec_3 & io_in_req_valid & _outSelRespVec_T_1; // @[src/main/scala/bus/simplebus/Crossbar.scala 63:60]
  assign io_out_3_req_bits_addr = io_in_req_bits_addr; // @[src/main/scala/bus/simplebus/Crossbar.scala 64:24]
  assign io_out_3_req_bits_cmd = io_in_req_bits_cmd; // @[src/main/scala/bus/simplebus/Crossbar.scala 64:24]
  assign io_out_3_req_bits_wmask = io_in_req_bits_wmask; // @[src/main/scala/bus/simplebus/Crossbar.scala 64:24]
  assign io_out_3_req_bits_wdata = io_in_req_bits_wdata; // @[src/main/scala/bus/simplebus/Crossbar.scala 64:24]
  assign io_out_3_resp_ready = outSelRespVec_3 & io_in_resp_ready & state == 2'h1; // @[src/main/scala/bus/simplebus/Crossbar.scala 69:66]
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 32:22]
      state <= 2'h0; // @[src/main/scala/bus/simplebus/Crossbar.scala 32:22]
    end else if (2'h0 == state) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 51:18]
      if (reqInvalidAddr) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 54:29]
        state <= 2'h2; // @[src/main/scala/bus/simplebus/Crossbar.scala 54:37]
      end else if (_outSelRespVec_T) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 53:29]
        state <= 2'h1; // @[src/main/scala/bus/simplebus/Crossbar.scala 53:37]
      end
    end else if (2'h1 == state) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 51:18]
      state <= _GEN_6;
    end else if (2'h2 == state) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 51:18]
      state <= _GEN_6;
    end
    if (reset) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
      outSelRespVec_0 <= 1'h0; // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
    end else if (_outSelRespVec_T_2) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
      outSelRespVec_0 <= outSelVec_0; // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
    end
    if (reset) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
      outSelRespVec_1 <= 1'h0; // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
    end else if (_outSelRespVec_T_2) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
      outSelRespVec_1 <= outSelVec_1; // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
    end
    if (reset) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
      outSelRespVec_2 <= 1'h0; // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
    end else if (_outSelRespVec_T_2) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
      outSelRespVec_2 <= outSelVec_2; // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
    end
    if (reset) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
      outSelRespVec_3 <= 1'h0; // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
    end else if (_outSelRespVec_T_2) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
      outSelRespVec_3 <= outSelVec_3; // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
    end
    if (reset) begin // @[src/main/scala/utils/GTimer.scala 24:20]
      c <= 64'h0; // @[src/main/scala/utils/GTimer.scala 24:20]
    end else begin
      c <= _c_T_1; // @[src/main/scala/utils/GTimer.scala 25:7]
    end
    if (reset) begin // @[src/main/scala/utils/GTimer.scala 24:20]
      c_1 <= 64'h0; // @[src/main/scala/utils/GTimer.scala 24:20]
    end else begin
      c_1 <= _c_T_3; // @[src/main/scala/utils/GTimer.scala 25:7]
    end
    if (reset) begin // @[src/main/scala/utils/GTimer.scala 24:20]
      c_2 <= 64'h0; // @[src/main/scala/utils/GTimer.scala 24:20]
    end else begin
      c_2 <= _c_T_5; // @[src/main/scala/utils/GTimer.scala 25:7]
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (reqInvalidAddr & DISPLAY_ENABLE & ~reset) begin
          $fwrite(32'h80000002,"crossbar access bad addr %x, time %d\n",io_in_req_bits_addr,c); // @[src/main/scala/bus/simplebus/Crossbar.scala 46:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2 & ~(~reqInvalidAddr)) begin
          $fwrite(32'h80000002,
            "Assertion failed: address decode error, bad addr = 0x%x\n\n    at Crossbar.scala:49 assert(!reqInvalidAddr, \"address decode error, bad addr = 0x%%%%x\\n\", addr)\n"
            ,io_in_req_bits_addr); // @[src/main/scala/bus/simplebus/Crossbar.scala 49:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~reqInvalidAddr) & _T_2) begin
          $fatal; // @[src/main/scala/bus/simplebus/Crossbar.scala 49:9]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _outSelRespVec_T & _T_2) begin
          $fwrite(32'h80000002,
            "%d: xbar: outSelVec = Vec(%d, %d, %d, %d), outSel.req: addr = 0x%x, cmd = %d, size = %d, wmask = 0x%x, wdata = 0x%x\n"
            ,c_1,outSelVec_0,outSelVec_1,outSelVec_2,outSelVec_3,io_in_req_bits_addr,io_in_req_bits_cmd,
            io_in_req_bits_size,io_in_req_bits_wmask,io_in_req_bits_wdata); // @[src/main/scala/bus/simplebus/Crossbar.scala 77:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_10 & _T_2) begin
          $fwrite(32'h80000002,"%d: xbar: outSelVec = Vec(%d, %d, %d, %d), outSel.resp: rdata = %x, cmd = %d\n",c_2,
            outSelVec_0,outSelVec_1,outSelVec_2,outSelVec_3,io_in_resp_bits_rdata,io_in_resp_bits_cmd); // @[src/main/scala/bus/simplebus/Crossbar.scala 80:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  outSelRespVec_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  outSelRespVec_1 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  outSelRespVec_2 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  outSelRespVec_3 = _RAND_4[0:0];
  _RAND_5 = {2{`RANDOM}};
  c = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  c_1 = _RAND_6[63:0];
  _RAND_7 = {2{`RANDOM}};
  c_2 = _RAND_7[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module AXI4UART(
  input         clock,
  input         reset,
  output        io_in_aw_ready, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input         io_in_aw_valid, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input  [31:0] io_in_aw_bits_addr, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output        io_in_w_ready, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input         io_in_w_valid, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input  [63:0] io_in_w_bits_data, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input  [7:0]  io_in_w_bits_strb, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input         io_in_b_ready, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output        io_in_b_valid, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output        io_in_ar_ready, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input         io_in_ar_valid, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input  [31:0] io_in_ar_bits_addr, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input         io_in_r_ready, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output        io_in_r_valid, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output [63:0] io_in_r_bits_data, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output        io_extra_out_valid, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output [7:0]  io_extra_out_ch, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output        io_extra_in_valid, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input  [7:0]  io_extra_in_ch // @[src/main/scala/device/AXI4Slave.scala 28:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
`endif // RANDOMIZE_REG_INIT
  wire  _r_busy_T = io_in_ar_ready & io_in_ar_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  wire  _r_busy_T_1 = io_in_r_ready & io_in_r_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  reg  r_busy; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  _GEN_0 = _r_busy_T_1 ? 1'h0 : r_busy; // @[src/main/scala/utils/StopWatch.scala 26:19 24:20 26:23]
  wire  _GEN_1 = _r_busy_T | _GEN_0; // @[src/main/scala/utils/StopWatch.scala 27:{20,24}]
  reg  ren_REG; // @[src/main/scala/device/AXI4Slave.scala 73:17]
  wire  _io_in_r_valid_T_2 = ren_REG & (_r_busy_T | r_busy); // @[src/main/scala/device/AXI4Slave.scala 74:35]
  reg  io_in_r_valid_r; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  _GEN_2 = _r_busy_T_1 ? 1'h0 : io_in_r_valid_r; // @[src/main/scala/utils/StopWatch.scala 26:19 24:20 26:23]
  wire  _GEN_3 = _io_in_r_valid_T_2 | _GEN_2; // @[src/main/scala/utils/StopWatch.scala 27:{20,24}]
  wire  _w_busy_T = io_in_aw_ready & io_in_aw_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  wire  _w_busy_T_1 = io_in_b_ready & io_in_b_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  reg  w_busy; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  _GEN_4 = _w_busy_T_1 ? 1'h0 : w_busy; // @[src/main/scala/utils/StopWatch.scala 26:19 24:20 26:23]
  wire  _GEN_5 = _w_busy_T | _GEN_4; // @[src/main/scala/utils/StopWatch.scala 27:{20,24}]
  wire  _io_in_b_valid_T = io_in_w_ready & io_in_w_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  reg  io_in_b_valid_r; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  _GEN_6 = _w_busy_T_1 ? 1'h0 : io_in_b_valid_r; // @[src/main/scala/utils/StopWatch.scala 26:19 24:20 26:23]
  wire  _GEN_7 = _io_in_b_valid_T | _GEN_6; // @[src/main/scala/utils/StopWatch.scala 27:{20,24}]
  reg [31:0] txfifo; // @[src/main/scala/device/AXI4UART.scala 29:19]
  reg [31:0] stat; // @[src/main/scala/device/AXI4UART.scala 30:21]
  reg [31:0] ctrl; // @[src/main/scala/device/AXI4UART.scala 31:21]
  wire  _io_extra_out_valid_T_1 = io_in_aw_bits_addr[3:0] == 4'h4; // @[src/main/scala/device/AXI4UART.scala 33:41]
  wire [7:0] _T_5 = io_in_w_bits_strb >> io_in_aw_bits_addr[2:0]; // @[src/main/scala/device/AXI4UART.scala 45:77]
  wire [7:0] _T_15 = _T_5[0] ? 8'hff : 8'h0; // @[src/main/scala/utils/BitUtils.scala 27:45]
  wire [7:0] _T_17 = _T_5[1] ? 8'hff : 8'h0; // @[src/main/scala/utils/BitUtils.scala 27:45]
  wire [7:0] _T_19 = _T_5[2] ? 8'hff : 8'h0; // @[src/main/scala/utils/BitUtils.scala 27:45]
  wire [7:0] _T_21 = _T_5[3] ? 8'hff : 8'h0; // @[src/main/scala/utils/BitUtils.scala 27:45]
  wire [7:0] _T_23 = _T_5[4] ? 8'hff : 8'h0; // @[src/main/scala/utils/BitUtils.scala 27:45]
  wire [7:0] _T_25 = _T_5[5] ? 8'hff : 8'h0; // @[src/main/scala/utils/BitUtils.scala 27:45]
  wire [7:0] _T_27 = _T_5[6] ? 8'hff : 8'h0; // @[src/main/scala/utils/BitUtils.scala 27:45]
  wire [7:0] _T_29 = _T_5[7] ? 8'hff : 8'h0; // @[src/main/scala/utils/BitUtils.scala 27:45]
  wire [63:0] _T_30 = {_T_29,_T_27,_T_25,_T_23,_T_21,_T_19,_T_17,_T_15}; // @[src/main/scala/utils/BitUtils.scala 27:26]
  wire  _io_in_r_bits_data_T = 4'h0 == io_in_ar_bits_addr[3:0]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _io_in_r_bits_data_T_1 = 4'h4 == io_in_ar_bits_addr[3:0]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _io_in_r_bits_data_T_2 = 4'h8 == io_in_ar_bits_addr[3:0]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _io_in_r_bits_data_T_3 = 4'hc == io_in_ar_bits_addr[3:0]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [7:0] _io_in_r_bits_data_T_4 = _io_in_r_bits_data_T ? io_extra_in_ch : 8'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] _io_in_r_bits_data_T_5 = _io_in_r_bits_data_T_1 ? txfifo : 32'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] _io_in_r_bits_data_T_6 = _io_in_r_bits_data_T_2 ? stat : 32'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] _io_in_r_bits_data_T_7 = _io_in_r_bits_data_T_3 ? ctrl : 32'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] _GEN_11 = {{24'd0}, _io_in_r_bits_data_T_4}; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] _io_in_r_bits_data_T_8 = _GEN_11 | _io_in_r_bits_data_T_5; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] _io_in_r_bits_data_T_9 = _io_in_r_bits_data_T_8 | _io_in_r_bits_data_T_6; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] _io_in_r_bits_data_T_10 = _io_in_r_bits_data_T_9 | _io_in_r_bits_data_T_7; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] _txfifo_T = io_in_w_bits_data[31:0] & _T_30[31:0]; // @[src/main/scala/utils/BitUtils.scala 34:14]
  wire [31:0] _txfifo_T_1 = ~_T_30[31:0]; // @[src/main/scala/utils/BitUtils.scala 34:39]
  wire [31:0] _txfifo_T_2 = txfifo & _txfifo_T_1; // @[src/main/scala/utils/BitUtils.scala 34:37]
  wire [31:0] _txfifo_T_3 = _txfifo_T | _txfifo_T_2; // @[src/main/scala/utils/BitUtils.scala 34:26]
  wire [31:0] _stat_T_2 = stat & _txfifo_T_1; // @[src/main/scala/utils/BitUtils.scala 34:37]
  wire [31:0] _stat_T_3 = _txfifo_T | _stat_T_2; // @[src/main/scala/utils/BitUtils.scala 34:26]
  wire [31:0] _ctrl_T_2 = ctrl & _txfifo_T_1; // @[src/main/scala/utils/BitUtils.scala 34:37]
  wire [31:0] _ctrl_T_3 = _txfifo_T | _ctrl_T_2; // @[src/main/scala/utils/BitUtils.scala 34:26]
  assign io_in_aw_ready = ~w_busy; // @[src/main/scala/device/AXI4Slave.scala 94:18]
  assign io_in_w_ready = io_in_aw_valid | w_busy; // @[src/main/scala/device/AXI4Slave.scala 95:30]
  assign io_in_b_valid = io_in_b_valid_r; // @[src/main/scala/device/AXI4Slave.scala 97:14]
  assign io_in_ar_ready = io_in_r_ready | ~r_busy; // @[src/main/scala/device/AXI4Slave.scala 71:29]
  assign io_in_r_valid = io_in_r_valid_r; // @[src/main/scala/device/AXI4Slave.scala 74:14]
  assign io_in_r_bits_data = {{32'd0}, _io_in_r_bits_data_T_10}; // @[src/main/scala/utils/RegMap.scala 30:11]
  assign io_extra_out_valid = io_in_aw_bits_addr[3:0] == 4'h4 & _io_in_b_valid_T; // @[src/main/scala/device/AXI4UART.scala 33:49]
  assign io_extra_out_ch = io_in_w_bits_data[7:0]; // @[src/main/scala/device/AXI4UART.scala 34:40]
  assign io_extra_in_valid = io_in_ar_bits_addr[3:0] == 4'h0 & _r_busy_T_1; // @[src/main/scala/device/AXI4UART.scala 35:48]
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      r_busy <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else begin
      r_busy <= _GEN_1;
    end
    if (reset) begin // @[src/main/scala/device/AXI4Slave.scala 73:17]
      ren_REG <= 1'h0; // @[src/main/scala/device/AXI4Slave.scala 73:17]
    end else begin
      ren_REG <= _r_busy_T; // @[src/main/scala/device/AXI4Slave.scala 73:17]
    end
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      io_in_r_valid_r <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else begin
      io_in_r_valid_r <= _GEN_3;
    end
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      w_busy <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else begin
      w_busy <= _GEN_5;
    end
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      io_in_b_valid_r <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else begin
      io_in_b_valid_r <= _GEN_7;
    end
    if (_io_in_b_valid_T & _io_extra_out_valid_T_1) begin // @[src/main/scala/utils/RegMap.scala 32:48]
      txfifo <= _txfifo_T_3; // @[src/main/scala/utils/RegMap.scala 32:52]
    end
    if (reset) begin // @[src/main/scala/device/AXI4UART.scala 30:21]
      stat <= 32'h1; // @[src/main/scala/device/AXI4UART.scala 30:21]
    end else if (_io_in_b_valid_T & io_in_aw_bits_addr[3:0] == 4'h8) begin // @[src/main/scala/utils/RegMap.scala 32:48]
      stat <= _stat_T_3; // @[src/main/scala/utils/RegMap.scala 32:52]
    end
    if (reset) begin // @[src/main/scala/device/AXI4UART.scala 31:21]
      ctrl <= 32'h0; // @[src/main/scala/device/AXI4UART.scala 31:21]
    end else if (_io_in_b_valid_T & io_in_aw_bits_addr[3:0] == 4'hc) begin // @[src/main/scala/utils/RegMap.scala 32:48]
      ctrl <= _ctrl_T_3; // @[src/main/scala/utils/RegMap.scala 32:52]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  r_busy = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  ren_REG = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  io_in_r_valid_r = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  w_busy = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  io_in_b_valid_r = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  txfifo = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  stat = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  ctrl = _RAND_7[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module AXI4Flash(
  input         clock,
  input         reset,
  output        io_in_aw_ready, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input         io_in_aw_valid, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output        io_in_w_ready, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input         io_in_w_valid, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input         io_in_b_ready, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output        io_in_b_valid, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output        io_in_ar_ready, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input         io_in_ar_valid, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input  [31:0] io_in_ar_bits_addr, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input         io_in_r_ready, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output        io_in_r_valid, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output [63:0] io_in_r_bits_data // @[src/main/scala/device/AXI4Slave.scala 28:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
`endif // RANDOMIZE_REG_INIT
  wire  _r_busy_T = io_in_ar_ready & io_in_ar_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  wire  _r_busy_T_1 = io_in_r_ready & io_in_r_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  reg  r_busy; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  _GEN_0 = _r_busy_T_1 ? 1'h0 : r_busy; // @[src/main/scala/utils/StopWatch.scala 26:19 24:20 26:23]
  wire  _GEN_1 = _r_busy_T | _GEN_0; // @[src/main/scala/utils/StopWatch.scala 27:{20,24}]
  reg  ren_REG; // @[src/main/scala/device/AXI4Slave.scala 73:17]
  wire  _io_in_r_valid_T_2 = ren_REG & (_r_busy_T | r_busy); // @[src/main/scala/device/AXI4Slave.scala 74:35]
  reg  io_in_r_valid_r; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  _GEN_2 = _r_busy_T_1 ? 1'h0 : io_in_r_valid_r; // @[src/main/scala/utils/StopWatch.scala 26:19 24:20 26:23]
  wire  _GEN_3 = _io_in_r_valid_T_2 | _GEN_2; // @[src/main/scala/utils/StopWatch.scala 27:{20,24}]
  wire  _w_busy_T = io_in_aw_ready & io_in_aw_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  wire  _w_busy_T_1 = io_in_b_ready & io_in_b_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  reg  w_busy; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  _GEN_4 = _w_busy_T_1 ? 1'h0 : w_busy; // @[src/main/scala/utils/StopWatch.scala 26:19 24:20 26:23]
  wire  _GEN_5 = _w_busy_T | _GEN_4; // @[src/main/scala/utils/StopWatch.scala 27:{20,24}]
  wire  _io_in_b_valid_T = io_in_w_ready & io_in_w_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  reg  io_in_b_valid_r; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  _GEN_6 = _w_busy_T_1 ? 1'h0 : io_in_b_valid_r; // @[src/main/scala/utils/StopWatch.scala 26:19 24:20 26:23]
  wire  _GEN_7 = _io_in_b_valid_T | _GEN_6; // @[src/main/scala/utils/StopWatch.scala 27:{20,24}]
  wire  _rdata_T = 13'h0 == io_in_ar_bits_addr[12:0]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _rdata_T_1 = 13'h4 == io_in_ar_bits_addr[12:0]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _rdata_T_2 = 13'h8 == io_in_ar_bits_addr[12:0]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [20:0] _rdata_T_3 = _rdata_T ? 21'h10029b : 21'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [24:0] _rdata_T_4 = _rdata_T_1 ? 25'h1f29293 : 25'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [17:0] _rdata_T_5 = _rdata_T_2 ? 18'h28067 : 18'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [24:0] _GEN_9 = {{4'd0}, _rdata_T_3}; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [24:0] _rdata_T_6 = _GEN_9 | _rdata_T_4; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [24:0] _GEN_10 = {{7'd0}, _rdata_T_5}; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [24:0] _rdata_T_7 = _rdata_T_6 | _GEN_10; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] rdata = {{39'd0}, _rdata_T_7}; // @[src/main/scala/device/AXI4Flash.scala 37:19 src/main/scala/utils/RegMap.scala 30:11]
  reg [63:0] io_in_r_bits_data_REG; // @[src/main/scala/device/AXI4Flash.scala 41:38]
  reg [63:0] io_in_r_bits_data_r; // @[src/main/scala/device/AXI4Flash.scala 41:30]
  assign io_in_aw_ready = ~w_busy; // @[src/main/scala/device/AXI4Slave.scala 94:18]
  assign io_in_w_ready = io_in_aw_valid | w_busy; // @[src/main/scala/device/AXI4Slave.scala 95:30]
  assign io_in_b_valid = io_in_b_valid_r; // @[src/main/scala/device/AXI4Slave.scala 97:14]
  assign io_in_ar_ready = io_in_r_ready | ~r_busy; // @[src/main/scala/device/AXI4Slave.scala 71:29]
  assign io_in_r_valid = io_in_r_valid_r; // @[src/main/scala/device/AXI4Slave.scala 74:14]
  assign io_in_r_bits_data = io_in_r_bits_data_r; // @[src/main/scala/device/AXI4Flash.scala 41:18]
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      r_busy <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else begin
      r_busy <= _GEN_1;
    end
    if (reset) begin // @[src/main/scala/device/AXI4Slave.scala 73:17]
      ren_REG <= 1'h0; // @[src/main/scala/device/AXI4Slave.scala 73:17]
    end else begin
      ren_REG <= _r_busy_T; // @[src/main/scala/device/AXI4Slave.scala 73:17]
    end
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      io_in_r_valid_r <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else begin
      io_in_r_valid_r <= _GEN_3;
    end
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      w_busy <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else begin
      w_busy <= _GEN_5;
    end
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      io_in_b_valid_r <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else begin
      io_in_b_valid_r <= _GEN_7;
    end
    io_in_r_bits_data_REG <= {rdata[31:0],rdata[31:0]}; // @[src/main/scala/device/AXI4Flash.scala 41:43]
    if (ren_REG) begin // @[src/main/scala/device/AXI4Flash.scala 41:30]
      io_in_r_bits_data_r <= io_in_r_bits_data_REG; // @[src/main/scala/device/AXI4Flash.scala 41:30]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  r_busy = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  ren_REG = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  io_in_r_valid_r = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  w_busy = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  io_in_b_valid_r = _RAND_4[0:0];
  _RAND_5 = {2{`RANDOM}};
  io_in_r_bits_data_REG = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  io_in_r_bits_data_r = _RAND_6[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module AXI4MeipGen(
  input         clock,
  input         reset,
  output        io_in_aw_ready, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input         io_in_aw_valid, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input  [31:0] io_in_aw_bits_addr, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output        io_in_w_ready, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input         io_in_w_valid, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input  [63:0] io_in_w_bits_data, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input  [7:0]  io_in_w_bits_strb, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input         io_in_b_ready, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output        io_in_b_valid, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output        io_in_ar_ready, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input         io_in_ar_valid, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input         io_in_r_ready, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output        io_in_r_valid, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output [63:0] io_in_r_bits_data, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output        io_extra_meip // @[src/main/scala/device/AXI4Slave.scala 28:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
`endif // RANDOMIZE_REG_INIT
  wire [7:0] _fullMask_T_9 = io_in_w_bits_strb[0] ? 8'hff : 8'h0; // @[src/main/scala/utils/BitUtils.scala 27:45]
  wire [7:0] _fullMask_T_11 = io_in_w_bits_strb[1] ? 8'hff : 8'h0; // @[src/main/scala/utils/BitUtils.scala 27:45]
  wire [7:0] _fullMask_T_13 = io_in_w_bits_strb[2] ? 8'hff : 8'h0; // @[src/main/scala/utils/BitUtils.scala 27:45]
  wire [7:0] _fullMask_T_15 = io_in_w_bits_strb[3] ? 8'hff : 8'h0; // @[src/main/scala/utils/BitUtils.scala 27:45]
  wire [7:0] _fullMask_T_17 = io_in_w_bits_strb[4] ? 8'hff : 8'h0; // @[src/main/scala/utils/BitUtils.scala 27:45]
  wire [7:0] _fullMask_T_19 = io_in_w_bits_strb[5] ? 8'hff : 8'h0; // @[src/main/scala/utils/BitUtils.scala 27:45]
  wire [7:0] _fullMask_T_21 = io_in_w_bits_strb[6] ? 8'hff : 8'h0; // @[src/main/scala/utils/BitUtils.scala 27:45]
  wire [7:0] _fullMask_T_23 = io_in_w_bits_strb[7] ? 8'hff : 8'h0; // @[src/main/scala/utils/BitUtils.scala 27:45]
  wire [63:0] fullMask = {_fullMask_T_23,_fullMask_T_21,_fullMask_T_19,_fullMask_T_17,_fullMask_T_15,_fullMask_T_13,
    _fullMask_T_11,_fullMask_T_9}; // @[src/main/scala/utils/BitUtils.scala 27:26]
  wire  _r_busy_T = io_in_ar_ready & io_in_ar_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  wire  _r_busy_T_1 = io_in_r_ready & io_in_r_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  reg  r_busy; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  _GEN_0 = _r_busy_T_1 ? 1'h0 : r_busy; // @[src/main/scala/utils/StopWatch.scala 26:19 24:20 26:23]
  wire  _GEN_1 = _r_busy_T | _GEN_0; // @[src/main/scala/utils/StopWatch.scala 27:{20,24}]
  reg  ren_REG; // @[src/main/scala/device/AXI4Slave.scala 73:17]
  wire  _io_in_r_valid_T_2 = ren_REG & (_r_busy_T | r_busy); // @[src/main/scala/device/AXI4Slave.scala 74:35]
  reg  io_in_r_valid_r; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  _GEN_2 = _r_busy_T_1 ? 1'h0 : io_in_r_valid_r; // @[src/main/scala/utils/StopWatch.scala 26:19 24:20 26:23]
  wire  _GEN_3 = _io_in_r_valid_T_2 | _GEN_2; // @[src/main/scala/utils/StopWatch.scala 27:{20,24}]
  wire  _w_busy_T = io_in_aw_ready & io_in_aw_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  wire  _w_busy_T_1 = io_in_b_ready & io_in_b_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  reg  w_busy; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  _GEN_4 = _w_busy_T_1 ? 1'h0 : w_busy; // @[src/main/scala/utils/StopWatch.scala 26:19 24:20 26:23]
  wire  _GEN_5 = _w_busy_T | _GEN_4; // @[src/main/scala/utils/StopWatch.scala 27:{20,24}]
  wire  _io_in_b_valid_T = io_in_w_ready & io_in_w_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  reg  io_in_b_valid_r; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  _GEN_6 = _w_busy_T_1 ? 1'h0 : io_in_b_valid_r; // @[src/main/scala/utils/StopWatch.scala 26:19 24:20 26:23]
  wire  _GEN_7 = _io_in_b_valid_T | _GEN_6; // @[src/main/scala/utils/StopWatch.scala 27:{20,24}]
  reg  meip; // @[src/main/scala/sim/MeipGen.scala 31:21]
  wire  _meip_T_3 = io_in_w_bits_data[0] & fullMask[0] | meip & ~fullMask[0]; // @[src/main/scala/utils/BitUtils.scala 34:26]
  assign io_in_aw_ready = ~w_busy; // @[src/main/scala/device/AXI4Slave.scala 94:18]
  assign io_in_w_ready = io_in_aw_valid | w_busy; // @[src/main/scala/device/AXI4Slave.scala 95:30]
  assign io_in_b_valid = io_in_b_valid_r; // @[src/main/scala/device/AXI4Slave.scala 97:14]
  assign io_in_ar_ready = io_in_r_ready | ~r_busy; // @[src/main/scala/device/AXI4Slave.scala 71:29]
  assign io_in_r_valid = io_in_r_valid_r; // @[src/main/scala/device/AXI4Slave.scala 74:14]
  assign io_in_r_bits_data = {{63'd0}, meip}; // @[src/main/scala/utils/RegMap.scala 30:11]
  assign io_extra_meip = meip; // @[src/main/scala/sim/MeipGen.scala 41:21]
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      r_busy <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else begin
      r_busy <= _GEN_1;
    end
    if (reset) begin // @[src/main/scala/device/AXI4Slave.scala 73:17]
      ren_REG <= 1'h0; // @[src/main/scala/device/AXI4Slave.scala 73:17]
    end else begin
      ren_REG <= _r_busy_T; // @[src/main/scala/device/AXI4Slave.scala 73:17]
    end
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      io_in_r_valid_r <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else begin
      io_in_r_valid_r <= _GEN_3;
    end
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      w_busy <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else begin
      w_busy <= _GEN_5;
    end
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      io_in_b_valid_r <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else begin
      io_in_b_valid_r <= _GEN_7;
    end
    if (reset) begin // @[src/main/scala/sim/MeipGen.scala 31:21]
      meip <= 1'h0; // @[src/main/scala/sim/MeipGen.scala 31:21]
    end else if (_io_in_b_valid_T & io_in_aw_bits_addr[3:0] == 4'h0) begin // @[src/main/scala/utils/RegMap.scala 32:48]
      meip <= _meip_T_3; // @[src/main/scala/utils/RegMap.scala 32:52]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  r_busy = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  ren_REG = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  io_in_r_valid_r = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  w_busy = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  io_in_b_valid_r = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  meip = _RAND_5[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module AXI4DMA(
  input         clock,
  input         reset,
  output        io_in_aw_ready, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input         io_in_aw_valid, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input  [31:0] io_in_aw_bits_addr, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output        io_in_w_ready, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input         io_in_w_valid, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input  [63:0] io_in_w_bits_data, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input  [7:0]  io_in_w_bits_strb, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input         io_in_b_ready, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output        io_in_b_valid, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output        io_in_ar_ready, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input         io_in_ar_valid, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input  [31:0] io_in_ar_bits_addr, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input         io_in_r_ready, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output        io_in_r_valid, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output [63:0] io_in_r_bits_data, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input         io_extra_dma_aw_ready, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output        io_extra_dma_aw_valid, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output [31:0] io_extra_dma_aw_bits_addr, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output [7:0]  io_extra_dma_aw_bits_len, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output [2:0]  io_extra_dma_aw_bits_size, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input         io_extra_dma_w_ready, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output        io_extra_dma_w_valid, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output [63:0] io_extra_dma_w_bits_data, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output [7:0]  io_extra_dma_w_bits_strb, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output        io_extra_dma_w_bits_last, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output        io_extra_dma_b_ready, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input         io_extra_dma_b_valid, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input         io_extra_dma_ar_ready, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output        io_extra_dma_ar_valid, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output [31:0] io_extra_dma_ar_bits_addr, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output [7:0]  io_extra_dma_ar_bits_len, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output [2:0]  io_extra_dma_ar_bits_size, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output        io_extra_dma_r_ready, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input         io_extra_dma_r_valid, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input  [63:0] io_extra_dma_r_bits_data // @[src/main/scala/device/AXI4Slave.scala 28:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
`endif // RANDOMIZE_REG_INIT
  wire  _r_busy_T = io_in_ar_ready & io_in_ar_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  wire  _r_busy_T_1 = io_in_r_ready & io_in_r_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  reg  r_busy; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  _GEN_0 = _r_busy_T_1 ? 1'h0 : r_busy; // @[src/main/scala/utils/StopWatch.scala 26:19 24:20 26:23]
  wire  _GEN_1 = _r_busy_T | _GEN_0; // @[src/main/scala/utils/StopWatch.scala 27:{20,24}]
  reg  ren_REG; // @[src/main/scala/device/AXI4Slave.scala 73:17]
  wire  _io_in_r_valid_T_2 = ren_REG & (_r_busy_T | r_busy); // @[src/main/scala/device/AXI4Slave.scala 74:35]
  reg  io_in_r_valid_r; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  _GEN_2 = _r_busy_T_1 ? 1'h0 : io_in_r_valid_r; // @[src/main/scala/utils/StopWatch.scala 26:19 24:20 26:23]
  wire  _GEN_3 = _io_in_r_valid_T_2 | _GEN_2; // @[src/main/scala/utils/StopWatch.scala 27:{20,24}]
  wire  _w_busy_T = io_in_aw_ready & io_in_aw_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  wire  _w_busy_T_1 = io_in_b_ready & io_in_b_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  reg  w_busy; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  _GEN_4 = _w_busy_T_1 ? 1'h0 : w_busy; // @[src/main/scala/utils/StopWatch.scala 26:19 24:20 26:23]
  wire  _GEN_5 = _w_busy_T | _GEN_4; // @[src/main/scala/utils/StopWatch.scala 27:{20,24}]
  wire  _io_in_b_valid_T = io_in_w_ready & io_in_w_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  reg  io_in_b_valid_r; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  _GEN_6 = _w_busy_T_1 ? 1'h0 : io_in_b_valid_r; // @[src/main/scala/utils/StopWatch.scala 26:19 24:20 26:23]
  wire  _GEN_7 = _io_in_b_valid_T | _GEN_6; // @[src/main/scala/utils/StopWatch.scala 27:{20,24}]
  reg [31:0] dest; // @[src/main/scala/device/AXI4DMA.scala 34:17]
  reg [31:0] src; // @[src/main/scala/device/AXI4DMA.scala 35:16]
  reg [31:0] len; // @[src/main/scala/device/AXI4DMA.scala 36:20]
  reg [31:0] data; // @[src/main/scala/device/AXI4DMA.scala 39:17]
  reg [2:0] state; // @[src/main/scala/device/AXI4DMA.scala 42:22]
  wire [2:0] _GEN_8 = state == 3'h0 & len != 32'h0 ? 3'h1 : state; // @[src/main/scala/device/AXI4DMA.scala 42:22 52:{42,50}]
  wire  _T_4 = io_extra_dma_ar_ready & io_extra_dma_ar_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  wire [2:0] _GEN_9 = state == 3'h1 & _T_4 ? 3'h2 : _GEN_8; // @[src/main/scala/device/AXI4DMA.scala 53:{46,54}]
  wire  _T_7 = io_extra_dma_r_ready & io_extra_dma_r_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  wire  _awAck_T = io_extra_dma_aw_ready & io_extra_dma_aw_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  reg  awAck; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  _GEN_14 = _awAck_T | awAck; // @[src/main/scala/utils/StopWatch.scala 24:20 30:{20,24}]
  wire  _wSend_T_1 = io_extra_dma_w_ready & io_extra_dma_w_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  reg  wAck; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  wSend = _awAck_T & _wSend_T_1 & io_extra_dma_w_bits_last | awAck & wAck; // @[src/main/scala/device/AXI4DMA.scala 63:49]
  wire  _wAck_T_1 = _wSend_T_1 & io_extra_dma_w_bits_last; // @[src/main/scala/device/AXI4DMA.scala 62:39]
  wire  _GEN_16 = _wAck_T_1 | wAck; // @[src/main/scala/utils/StopWatch.scala 24:20 30:{20,24}]
  wire  _T_9 = state == 3'h3; // @[src/main/scala/device/AXI4DMA.scala 65:15]
  wire  _T_12 = io_extra_dma_b_ready & io_extra_dma_b_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  wire [31:0] _len_T_1 = len - 32'h4; // @[src/main/scala/device/AXI4DMA.scala 67:16]
  wire [31:0] _dest_T_1 = dest + 32'h4; // @[src/main/scala/device/AXI4DMA.scala 68:18]
  wire [31:0] _src_T_1 = src + 32'h4; // @[src/main/scala/device/AXI4DMA.scala 69:16]
  wire [3:0] _io_extra_dma_w_bits_strb_T_2 = dest[2] * 3'h4; // @[src/main/scala/device/AXI4DMA.scala 91:68]
  wire [18:0] _io_extra_dma_w_bits_strb_T_3 = 19'hf << _io_extra_dma_w_bits_strb_T_2; // @[src/main/scala/device/AXI4DMA.scala 91:41]
  wire [7:0] _T_19 = io_in_w_bits_strb >> io_in_aw_bits_addr[2:0]; // @[src/main/scala/device/AXI4DMA.scala 102:77]
  wire [7:0] _T_29 = _T_19[0] ? 8'hff : 8'h0; // @[src/main/scala/utils/BitUtils.scala 27:45]
  wire [7:0] _T_31 = _T_19[1] ? 8'hff : 8'h0; // @[src/main/scala/utils/BitUtils.scala 27:45]
  wire [7:0] _T_33 = _T_19[2] ? 8'hff : 8'h0; // @[src/main/scala/utils/BitUtils.scala 27:45]
  wire [7:0] _T_35 = _T_19[3] ? 8'hff : 8'h0; // @[src/main/scala/utils/BitUtils.scala 27:45]
  wire [7:0] _T_37 = _T_19[4] ? 8'hff : 8'h0; // @[src/main/scala/utils/BitUtils.scala 27:45]
  wire [7:0] _T_39 = _T_19[5] ? 8'hff : 8'h0; // @[src/main/scala/utils/BitUtils.scala 27:45]
  wire [7:0] _T_41 = _T_19[6] ? 8'hff : 8'h0; // @[src/main/scala/utils/BitUtils.scala 27:45]
  wire [7:0] _T_43 = _T_19[7] ? 8'hff : 8'h0; // @[src/main/scala/utils/BitUtils.scala 27:45]
  wire [63:0] _T_44 = {_T_43,_T_41,_T_39,_T_37,_T_35,_T_33,_T_31,_T_29}; // @[src/main/scala/utils/BitUtils.scala 27:26]
  wire  _io_in_r_bits_data_T = 4'h0 == io_in_ar_bits_addr[3:0]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _io_in_r_bits_data_T_1 = 4'h4 == io_in_ar_bits_addr[3:0]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _io_in_r_bits_data_T_2 = 4'h8 == io_in_ar_bits_addr[3:0]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [31:0] _io_in_r_bits_data_T_3 = _io_in_r_bits_data_T ? dest : 32'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] _io_in_r_bits_data_T_4 = _io_in_r_bits_data_T_1 ? src : 32'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] _io_in_r_bits_data_T_5 = _io_in_r_bits_data_T_2 ? len : 32'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] _io_in_r_bits_data_T_6 = _io_in_r_bits_data_T_3 | _io_in_r_bits_data_T_4; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] _io_in_r_bits_data_T_7 = _io_in_r_bits_data_T_6 | _io_in_r_bits_data_T_5; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] _dest_T_2 = io_in_w_bits_data[31:0] & _T_44[31:0]; // @[src/main/scala/utils/BitUtils.scala 34:14]
  wire [31:0] _dest_T_3 = ~_T_44[31:0]; // @[src/main/scala/utils/BitUtils.scala 34:39]
  wire [31:0] _dest_T_4 = dest & _dest_T_3; // @[src/main/scala/utils/BitUtils.scala 34:37]
  wire [31:0] _dest_T_5 = _dest_T_2 | _dest_T_4; // @[src/main/scala/utils/BitUtils.scala 34:26]
  wire [31:0] _src_T_4 = src & _dest_T_3; // @[src/main/scala/utils/BitUtils.scala 34:37]
  wire [31:0] _src_T_5 = _dest_T_2 | _src_T_4; // @[src/main/scala/utils/BitUtils.scala 34:26]
  wire [31:0] _len_T_4 = len & _dest_T_3; // @[src/main/scala/utils/BitUtils.scala 34:37]
  wire [31:0] _len_T_5 = _dest_T_2 | _len_T_4; // @[src/main/scala/utils/BitUtils.scala 34:26]
  assign io_in_aw_ready = ~w_busy; // @[src/main/scala/device/AXI4Slave.scala 94:18]
  assign io_in_w_ready = io_in_aw_valid | w_busy; // @[src/main/scala/device/AXI4Slave.scala 95:30]
  assign io_in_b_valid = io_in_b_valid_r; // @[src/main/scala/device/AXI4Slave.scala 97:14]
  assign io_in_ar_ready = io_in_r_ready | ~r_busy; // @[src/main/scala/device/AXI4Slave.scala 71:29]
  assign io_in_r_valid = io_in_r_valid_r; // @[src/main/scala/device/AXI4Slave.scala 74:14]
  assign io_in_r_bits_data = {{32'd0}, _io_in_r_bits_data_T_7}; // @[src/main/scala/utils/RegMap.scala 30:11]
  assign io_extra_dma_aw_valid = _T_9 & ~awAck; // @[src/main/scala/device/AXI4DMA.scala 88:43]
  assign io_extra_dma_aw_bits_addr = dest; // @[src/main/scala/device/AXI4DMA.scala 87:20]
  assign io_extra_dma_aw_bits_len = io_extra_dma_ar_bits_len; // @[src/main/scala/device/AXI4DMA.scala 86:15]
  assign io_extra_dma_aw_bits_size = io_extra_dma_ar_bits_size; // @[src/main/scala/device/AXI4DMA.scala 86:15]
  assign io_extra_dma_w_valid = _T_9 & ~wAck; // @[src/main/scala/device/AXI4DMA.scala 89:42]
  assign io_extra_dma_w_bits_data = {data,data}; // @[src/main/scala/device/AXI4DMA.scala 90:26]
  assign io_extra_dma_w_bits_strb = _io_extra_dma_w_bits_strb_T_3[7:0]; // @[src/main/scala/device/AXI4DMA.scala 91:19]
  assign io_extra_dma_w_bits_last = 1'h1; // @[src/main/scala/device/AXI4DMA.scala 92:19]
  assign io_extra_dma_b_ready = state == 3'h4; // @[src/main/scala/device/AXI4DMA.scala 93:25]
  assign io_extra_dma_ar_valid = state == 3'h1; // @[src/main/scala/device/AXI4DMA.scala 83:26]
  assign io_extra_dma_ar_bits_addr = src; // @[src/main/scala/device/AXI4DMA.scala 82:20]
  assign io_extra_dma_ar_bits_len = 8'h0; // @[src/main/scala/device/AXI4DMA.scala 81:19]
  assign io_extra_dma_ar_bits_size = 3'h2; // @[src/main/scala/device/AXI4DMA.scala 75:20]
  assign io_extra_dma_r_ready = state == 3'h2; // @[src/main/scala/device/AXI4DMA.scala 84:25]
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      r_busy <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else begin
      r_busy <= _GEN_1;
    end
    if (reset) begin // @[src/main/scala/device/AXI4Slave.scala 73:17]
      ren_REG <= 1'h0; // @[src/main/scala/device/AXI4Slave.scala 73:17]
    end else begin
      ren_REG <= _r_busy_T; // @[src/main/scala/device/AXI4Slave.scala 73:17]
    end
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      io_in_r_valid_r <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else begin
      io_in_r_valid_r <= _GEN_3;
    end
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      w_busy <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else begin
      w_busy <= _GEN_5;
    end
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      io_in_b_valid_r <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else begin
      io_in_b_valid_r <= _GEN_7;
    end
    if (_io_in_b_valid_T & io_in_aw_bits_addr[3:0] == 4'h0) begin // @[src/main/scala/utils/RegMap.scala 32:48]
      dest <= _dest_T_5; // @[src/main/scala/utils/RegMap.scala 32:52]
    end else if (state == 3'h4 & _T_12) begin // @[src/main/scala/device/AXI4DMA.scala 66:52]
      dest <= _dest_T_1; // @[src/main/scala/device/AXI4DMA.scala 68:10]
    end
    if (_io_in_b_valid_T & io_in_aw_bits_addr[3:0] == 4'h4) begin // @[src/main/scala/utils/RegMap.scala 32:48]
      src <= _src_T_5; // @[src/main/scala/utils/RegMap.scala 32:52]
    end else if (state == 3'h4 & _T_12) begin // @[src/main/scala/device/AXI4DMA.scala 66:52]
      src <= _src_T_1; // @[src/main/scala/device/AXI4DMA.scala 69:9]
    end
    if (reset) begin // @[src/main/scala/device/AXI4DMA.scala 36:20]
      len <= 32'h0; // @[src/main/scala/device/AXI4DMA.scala 36:20]
    end else if (_io_in_b_valid_T & io_in_aw_bits_addr[3:0] == 4'h8) begin // @[src/main/scala/utils/RegMap.scala 32:48]
      len <= _len_T_5; // @[src/main/scala/utils/RegMap.scala 32:52]
    end else if (state == 3'h4 & _T_12) begin // @[src/main/scala/device/AXI4DMA.scala 66:52]
      len <= _len_T_1; // @[src/main/scala/device/AXI4DMA.scala 67:9]
    end
    if (state == 3'h2 & _T_7) begin // @[src/main/scala/device/AXI4DMA.scala 54:51]
      if (src[2]) begin // @[src/main/scala/device/AXI4DMA.scala 55:10]
        data <= io_extra_dma_r_bits_data[63:32]; // @[src/main/scala/device/AXI4DMA.scala 55:10]
      end else begin
        data <= io_extra_dma_r_bits_data[31:0];
      end
    end
    if (reset) begin // @[src/main/scala/device/AXI4DMA.scala 42:22]
      state <= 3'h0; // @[src/main/scala/device/AXI4DMA.scala 42:22]
    end else if (state == 3'h4 & _T_12) begin // @[src/main/scala/device/AXI4DMA.scala 66:52]
      if (len <= 32'h4) begin // @[src/main/scala/device/AXI4DMA.scala 70:17]
        state <= 3'h0;
      end else begin
        state <= 3'h1;
      end
    end else if (state == 3'h3 & wSend) begin // @[src/main/scala/device/AXI4DMA.scala 65:41]
      state <= 3'h4; // @[src/main/scala/device/AXI4DMA.scala 65:49]
    end else if (state == 3'h2 & _T_7) begin // @[src/main/scala/device/AXI4DMA.scala 54:51]
      state <= 3'h3; // @[src/main/scala/device/AXI4DMA.scala 56:11]
    end else begin
      state <= _GEN_9;
    end
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      awAck <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else if (wSend) begin // @[src/main/scala/utils/StopWatch.scala 31:19]
      awAck <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 31:23]
    end else begin
      awAck <= _GEN_14;
    end
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      wAck <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else if (wSend) begin // @[src/main/scala/utils/StopWatch.scala 31:19]
      wAck <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 31:23]
    end else begin
      wAck <= _GEN_16;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  r_busy = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  ren_REG = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  io_in_r_valid_r = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  w_busy = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  io_in_b_valid_r = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  dest = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  src = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  len = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  data = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  state = _RAND_9[2:0];
  _RAND_10 = {1{`RANDOM}};
  awAck = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  wAck = _RAND_11[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module SimMMIO(
  input         clock,
  input         reset,
  output        io_rw_req_ready, // @[src/main/scala/sim/SimMMIO.scala 28:14]
  input         io_rw_req_valid, // @[src/main/scala/sim/SimMMIO.scala 28:14]
  input  [31:0] io_rw_req_bits_addr, // @[src/main/scala/sim/SimMMIO.scala 28:14]
  input  [2:0]  io_rw_req_bits_size, // @[src/main/scala/sim/SimMMIO.scala 28:14]
  input  [3:0]  io_rw_req_bits_cmd, // @[src/main/scala/sim/SimMMIO.scala 28:14]
  input  [7:0]  io_rw_req_bits_wmask, // @[src/main/scala/sim/SimMMIO.scala 28:14]
  input  [63:0] io_rw_req_bits_wdata, // @[src/main/scala/sim/SimMMIO.scala 28:14]
  input         io_rw_resp_ready, // @[src/main/scala/sim/SimMMIO.scala 28:14]
  output        io_rw_resp_valid, // @[src/main/scala/sim/SimMMIO.scala 28:14]
  output [3:0]  io_rw_resp_bits_cmd, // @[src/main/scala/sim/SimMMIO.scala 28:14]
  output [63:0] io_rw_resp_bits_rdata, // @[src/main/scala/sim/SimMMIO.scala 28:14]
  output        io_meip, // @[src/main/scala/sim/SimMMIO.scala 28:14]
  input         io_dma_aw_ready, // @[src/main/scala/sim/SimMMIO.scala 28:14]
  output        io_dma_aw_valid, // @[src/main/scala/sim/SimMMIO.scala 28:14]
  output [31:0] io_dma_aw_bits_addr, // @[src/main/scala/sim/SimMMIO.scala 28:14]
  output [7:0]  io_dma_aw_bits_len, // @[src/main/scala/sim/SimMMIO.scala 28:14]
  output [2:0]  io_dma_aw_bits_size, // @[src/main/scala/sim/SimMMIO.scala 28:14]
  input         io_dma_w_ready, // @[src/main/scala/sim/SimMMIO.scala 28:14]
  output        io_dma_w_valid, // @[src/main/scala/sim/SimMMIO.scala 28:14]
  output [63:0] io_dma_w_bits_data, // @[src/main/scala/sim/SimMMIO.scala 28:14]
  output [7:0]  io_dma_w_bits_strb, // @[src/main/scala/sim/SimMMIO.scala 28:14]
  output        io_dma_b_ready, // @[src/main/scala/sim/SimMMIO.scala 28:14]
  input         io_dma_b_valid, // @[src/main/scala/sim/SimMMIO.scala 28:14]
  input         io_dma_ar_ready, // @[src/main/scala/sim/SimMMIO.scala 28:14]
  output        io_dma_ar_valid, // @[src/main/scala/sim/SimMMIO.scala 28:14]
  output [31:0] io_dma_ar_bits_addr, // @[src/main/scala/sim/SimMMIO.scala 28:14]
  output        io_dma_r_ready, // @[src/main/scala/sim/SimMMIO.scala 28:14]
  input         io_dma_r_valid, // @[src/main/scala/sim/SimMMIO.scala 28:14]
  input  [63:0] io_dma_r_bits_data, // @[src/main/scala/sim/SimMMIO.scala 28:14]
  output        io_uart_out_valid, // @[src/main/scala/sim/SimMMIO.scala 28:14]
  output [7:0]  io_uart_out_ch, // @[src/main/scala/sim/SimMMIO.scala 28:14]
  output        io_uart_in_valid, // @[src/main/scala/sim/SimMMIO.scala 28:14]
  input  [7:0]  io_uart_in_ch, // @[src/main/scala/sim/SimMMIO.scala 28:14]
  input         _WIRE_4
);
  wire  xbar_clock; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire  xbar_reset; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire  xbar_io_in_req_ready; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire  xbar_io_in_req_valid; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire [31:0] xbar_io_in_req_bits_addr; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire [2:0] xbar_io_in_req_bits_size; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire [3:0] xbar_io_in_req_bits_cmd; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire [7:0] xbar_io_in_req_bits_wmask; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire [63:0] xbar_io_in_req_bits_wdata; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire  xbar_io_in_resp_ready; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire  xbar_io_in_resp_valid; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire [3:0] xbar_io_in_resp_bits_cmd; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire [63:0] xbar_io_in_resp_bits_rdata; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire  xbar_io_out_0_req_ready; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire  xbar_io_out_0_req_valid; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire [31:0] xbar_io_out_0_req_bits_addr; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire [3:0] xbar_io_out_0_req_bits_cmd; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire [7:0] xbar_io_out_0_req_bits_wmask; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire [63:0] xbar_io_out_0_req_bits_wdata; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire  xbar_io_out_0_resp_ready; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire  xbar_io_out_0_resp_valid; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire [63:0] xbar_io_out_0_resp_bits_rdata; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire  xbar_io_out_1_req_ready; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire  xbar_io_out_1_req_valid; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire [31:0] xbar_io_out_1_req_bits_addr; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire [3:0] xbar_io_out_1_req_bits_cmd; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire [7:0] xbar_io_out_1_req_bits_wmask; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire [63:0] xbar_io_out_1_req_bits_wdata; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire  xbar_io_out_1_resp_ready; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire  xbar_io_out_1_resp_valid; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire [63:0] xbar_io_out_1_resp_bits_rdata; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire  xbar_io_out_2_req_ready; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire  xbar_io_out_2_req_valid; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire [31:0] xbar_io_out_2_req_bits_addr; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire [3:0] xbar_io_out_2_req_bits_cmd; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire [7:0] xbar_io_out_2_req_bits_wmask; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire [63:0] xbar_io_out_2_req_bits_wdata; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire  xbar_io_out_2_resp_ready; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire  xbar_io_out_2_resp_valid; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire [63:0] xbar_io_out_2_resp_bits_rdata; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire  xbar_io_out_3_req_ready; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire  xbar_io_out_3_req_valid; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire [31:0] xbar_io_out_3_req_bits_addr; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire [3:0] xbar_io_out_3_req_bits_cmd; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire [7:0] xbar_io_out_3_req_bits_wmask; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire [63:0] xbar_io_out_3_req_bits_wdata; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire  xbar_io_out_3_resp_ready; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire  xbar_io_out_3_resp_valid; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire [63:0] xbar_io_out_3_resp_bits_rdata; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire  xbar_DISPLAY_ENABLE; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire  uart_clock; // @[src/main/scala/sim/SimMMIO.scala 48:20]
  wire  uart_reset; // @[src/main/scala/sim/SimMMIO.scala 48:20]
  wire  uart_io_in_aw_ready; // @[src/main/scala/sim/SimMMIO.scala 48:20]
  wire  uart_io_in_aw_valid; // @[src/main/scala/sim/SimMMIO.scala 48:20]
  wire [31:0] uart_io_in_aw_bits_addr; // @[src/main/scala/sim/SimMMIO.scala 48:20]
  wire  uart_io_in_w_ready; // @[src/main/scala/sim/SimMMIO.scala 48:20]
  wire  uart_io_in_w_valid; // @[src/main/scala/sim/SimMMIO.scala 48:20]
  wire [63:0] uart_io_in_w_bits_data; // @[src/main/scala/sim/SimMMIO.scala 48:20]
  wire [7:0] uart_io_in_w_bits_strb; // @[src/main/scala/sim/SimMMIO.scala 48:20]
  wire  uart_io_in_b_ready; // @[src/main/scala/sim/SimMMIO.scala 48:20]
  wire  uart_io_in_b_valid; // @[src/main/scala/sim/SimMMIO.scala 48:20]
  wire  uart_io_in_ar_ready; // @[src/main/scala/sim/SimMMIO.scala 48:20]
  wire  uart_io_in_ar_valid; // @[src/main/scala/sim/SimMMIO.scala 48:20]
  wire [31:0] uart_io_in_ar_bits_addr; // @[src/main/scala/sim/SimMMIO.scala 48:20]
  wire  uart_io_in_r_ready; // @[src/main/scala/sim/SimMMIO.scala 48:20]
  wire  uart_io_in_r_valid; // @[src/main/scala/sim/SimMMIO.scala 48:20]
  wire [63:0] uart_io_in_r_bits_data; // @[src/main/scala/sim/SimMMIO.scala 48:20]
  wire  uart_io_extra_out_valid; // @[src/main/scala/sim/SimMMIO.scala 48:20]
  wire [7:0] uart_io_extra_out_ch; // @[src/main/scala/sim/SimMMIO.scala 48:20]
  wire  uart_io_extra_in_valid; // @[src/main/scala/sim/SimMMIO.scala 48:20]
  wire [7:0] uart_io_extra_in_ch; // @[src/main/scala/sim/SimMMIO.scala 48:20]
  wire  flash_clock; // @[src/main/scala/sim/SimMMIO.scala 50:21]
  wire  flash_reset; // @[src/main/scala/sim/SimMMIO.scala 50:21]
  wire  flash_io_in_aw_ready; // @[src/main/scala/sim/SimMMIO.scala 50:21]
  wire  flash_io_in_aw_valid; // @[src/main/scala/sim/SimMMIO.scala 50:21]
  wire  flash_io_in_w_ready; // @[src/main/scala/sim/SimMMIO.scala 50:21]
  wire  flash_io_in_w_valid; // @[src/main/scala/sim/SimMMIO.scala 50:21]
  wire  flash_io_in_b_ready; // @[src/main/scala/sim/SimMMIO.scala 50:21]
  wire  flash_io_in_b_valid; // @[src/main/scala/sim/SimMMIO.scala 50:21]
  wire  flash_io_in_ar_ready; // @[src/main/scala/sim/SimMMIO.scala 50:21]
  wire  flash_io_in_ar_valid; // @[src/main/scala/sim/SimMMIO.scala 50:21]
  wire [31:0] flash_io_in_ar_bits_addr; // @[src/main/scala/sim/SimMMIO.scala 50:21]
  wire  flash_io_in_r_ready; // @[src/main/scala/sim/SimMMIO.scala 50:21]
  wire  flash_io_in_r_valid; // @[src/main/scala/sim/SimMMIO.scala 50:21]
  wire [63:0] flash_io_in_r_bits_data; // @[src/main/scala/sim/SimMMIO.scala 50:21]
  wire  meipGen_clock; // @[src/main/scala/sim/SimMMIO.scala 52:23]
  wire  meipGen_reset; // @[src/main/scala/sim/SimMMIO.scala 52:23]
  wire  meipGen_io_in_aw_ready; // @[src/main/scala/sim/SimMMIO.scala 52:23]
  wire  meipGen_io_in_aw_valid; // @[src/main/scala/sim/SimMMIO.scala 52:23]
  wire [31:0] meipGen_io_in_aw_bits_addr; // @[src/main/scala/sim/SimMMIO.scala 52:23]
  wire  meipGen_io_in_w_ready; // @[src/main/scala/sim/SimMMIO.scala 52:23]
  wire  meipGen_io_in_w_valid; // @[src/main/scala/sim/SimMMIO.scala 52:23]
  wire [63:0] meipGen_io_in_w_bits_data; // @[src/main/scala/sim/SimMMIO.scala 52:23]
  wire [7:0] meipGen_io_in_w_bits_strb; // @[src/main/scala/sim/SimMMIO.scala 52:23]
  wire  meipGen_io_in_b_ready; // @[src/main/scala/sim/SimMMIO.scala 52:23]
  wire  meipGen_io_in_b_valid; // @[src/main/scala/sim/SimMMIO.scala 52:23]
  wire  meipGen_io_in_ar_ready; // @[src/main/scala/sim/SimMMIO.scala 52:23]
  wire  meipGen_io_in_ar_valid; // @[src/main/scala/sim/SimMMIO.scala 52:23]
  wire  meipGen_io_in_r_ready; // @[src/main/scala/sim/SimMMIO.scala 52:23]
  wire  meipGen_io_in_r_valid; // @[src/main/scala/sim/SimMMIO.scala 52:23]
  wire [63:0] meipGen_io_in_r_bits_data; // @[src/main/scala/sim/SimMMIO.scala 52:23]
  wire  meipGen_io_extra_meip; // @[src/main/scala/sim/SimMMIO.scala 52:23]
  wire  dma_clock; // @[src/main/scala/sim/SimMMIO.scala 53:19]
  wire  dma_reset; // @[src/main/scala/sim/SimMMIO.scala 53:19]
  wire  dma_io_in_aw_ready; // @[src/main/scala/sim/SimMMIO.scala 53:19]
  wire  dma_io_in_aw_valid; // @[src/main/scala/sim/SimMMIO.scala 53:19]
  wire [31:0] dma_io_in_aw_bits_addr; // @[src/main/scala/sim/SimMMIO.scala 53:19]
  wire  dma_io_in_w_ready; // @[src/main/scala/sim/SimMMIO.scala 53:19]
  wire  dma_io_in_w_valid; // @[src/main/scala/sim/SimMMIO.scala 53:19]
  wire [63:0] dma_io_in_w_bits_data; // @[src/main/scala/sim/SimMMIO.scala 53:19]
  wire [7:0] dma_io_in_w_bits_strb; // @[src/main/scala/sim/SimMMIO.scala 53:19]
  wire  dma_io_in_b_ready; // @[src/main/scala/sim/SimMMIO.scala 53:19]
  wire  dma_io_in_b_valid; // @[src/main/scala/sim/SimMMIO.scala 53:19]
  wire  dma_io_in_ar_ready; // @[src/main/scala/sim/SimMMIO.scala 53:19]
  wire  dma_io_in_ar_valid; // @[src/main/scala/sim/SimMMIO.scala 53:19]
  wire [31:0] dma_io_in_ar_bits_addr; // @[src/main/scala/sim/SimMMIO.scala 53:19]
  wire  dma_io_in_r_ready; // @[src/main/scala/sim/SimMMIO.scala 53:19]
  wire  dma_io_in_r_valid; // @[src/main/scala/sim/SimMMIO.scala 53:19]
  wire [63:0] dma_io_in_r_bits_data; // @[src/main/scala/sim/SimMMIO.scala 53:19]
  wire  dma_io_extra_dma_aw_ready; // @[src/main/scala/sim/SimMMIO.scala 53:19]
  wire  dma_io_extra_dma_aw_valid; // @[src/main/scala/sim/SimMMIO.scala 53:19]
  wire [31:0] dma_io_extra_dma_aw_bits_addr; // @[src/main/scala/sim/SimMMIO.scala 53:19]
  wire [7:0] dma_io_extra_dma_aw_bits_len; // @[src/main/scala/sim/SimMMIO.scala 53:19]
  wire [2:0] dma_io_extra_dma_aw_bits_size; // @[src/main/scala/sim/SimMMIO.scala 53:19]
  wire  dma_io_extra_dma_w_ready; // @[src/main/scala/sim/SimMMIO.scala 53:19]
  wire  dma_io_extra_dma_w_valid; // @[src/main/scala/sim/SimMMIO.scala 53:19]
  wire [63:0] dma_io_extra_dma_w_bits_data; // @[src/main/scala/sim/SimMMIO.scala 53:19]
  wire [7:0] dma_io_extra_dma_w_bits_strb; // @[src/main/scala/sim/SimMMIO.scala 53:19]
  wire  dma_io_extra_dma_w_bits_last; // @[src/main/scala/sim/SimMMIO.scala 53:19]
  wire  dma_io_extra_dma_b_ready; // @[src/main/scala/sim/SimMMIO.scala 53:19]
  wire  dma_io_extra_dma_b_valid; // @[src/main/scala/sim/SimMMIO.scala 53:19]
  wire  dma_io_extra_dma_ar_ready; // @[src/main/scala/sim/SimMMIO.scala 53:19]
  wire  dma_io_extra_dma_ar_valid; // @[src/main/scala/sim/SimMMIO.scala 53:19]
  wire [31:0] dma_io_extra_dma_ar_bits_addr; // @[src/main/scala/sim/SimMMIO.scala 53:19]
  wire [7:0] dma_io_extra_dma_ar_bits_len; // @[src/main/scala/sim/SimMMIO.scala 53:19]
  wire [2:0] dma_io_extra_dma_ar_bits_size; // @[src/main/scala/sim/SimMMIO.scala 53:19]
  wire  dma_io_extra_dma_r_ready; // @[src/main/scala/sim/SimMMIO.scala 53:19]
  wire  dma_io_extra_dma_r_valid; // @[src/main/scala/sim/SimMMIO.scala 53:19]
  wire [63:0] dma_io_extra_dma_r_bits_data; // @[src/main/scala/sim/SimMMIO.scala 53:19]
  wire  uart_io_in_bridge_clock; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  uart_io_in_bridge_reset; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  uart_io_in_bridge_io_in_req_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  uart_io_in_bridge_io_in_req_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [31:0] uart_io_in_bridge_io_in_req_bits_addr; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [3:0] uart_io_in_bridge_io_in_req_bits_cmd; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [7:0] uart_io_in_bridge_io_in_req_bits_wmask; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [63:0] uart_io_in_bridge_io_in_req_bits_wdata; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  uart_io_in_bridge_io_in_resp_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  uart_io_in_bridge_io_in_resp_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [63:0] uart_io_in_bridge_io_in_resp_bits_rdata; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  uart_io_in_bridge_io_out_aw_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  uart_io_in_bridge_io_out_aw_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [31:0] uart_io_in_bridge_io_out_aw_bits_addr; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  uart_io_in_bridge_io_out_w_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  uart_io_in_bridge_io_out_w_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [63:0] uart_io_in_bridge_io_out_w_bits_data; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [7:0] uart_io_in_bridge_io_out_w_bits_strb; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  uart_io_in_bridge_io_out_b_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  uart_io_in_bridge_io_out_b_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  uart_io_in_bridge_io_out_ar_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  uart_io_in_bridge_io_out_ar_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [31:0] uart_io_in_bridge_io_out_ar_bits_addr; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  uart_io_in_bridge_io_out_r_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  uart_io_in_bridge_io_out_r_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [63:0] uart_io_in_bridge_io_out_r_bits_data; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  flash_io_in_bridge_clock; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  flash_io_in_bridge_reset; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  flash_io_in_bridge_io_in_req_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  flash_io_in_bridge_io_in_req_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [31:0] flash_io_in_bridge_io_in_req_bits_addr; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [3:0] flash_io_in_bridge_io_in_req_bits_cmd; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [7:0] flash_io_in_bridge_io_in_req_bits_wmask; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [63:0] flash_io_in_bridge_io_in_req_bits_wdata; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  flash_io_in_bridge_io_in_resp_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  flash_io_in_bridge_io_in_resp_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [63:0] flash_io_in_bridge_io_in_resp_bits_rdata; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  flash_io_in_bridge_io_out_aw_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  flash_io_in_bridge_io_out_aw_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [31:0] flash_io_in_bridge_io_out_aw_bits_addr; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  flash_io_in_bridge_io_out_w_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  flash_io_in_bridge_io_out_w_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [63:0] flash_io_in_bridge_io_out_w_bits_data; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [7:0] flash_io_in_bridge_io_out_w_bits_strb; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  flash_io_in_bridge_io_out_b_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  flash_io_in_bridge_io_out_b_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  flash_io_in_bridge_io_out_ar_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  flash_io_in_bridge_io_out_ar_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [31:0] flash_io_in_bridge_io_out_ar_bits_addr; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  flash_io_in_bridge_io_out_r_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  flash_io_in_bridge_io_out_r_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [63:0] flash_io_in_bridge_io_out_r_bits_data; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  meipGen_io_in_bridge_clock; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  meipGen_io_in_bridge_reset; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  meipGen_io_in_bridge_io_in_req_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  meipGen_io_in_bridge_io_in_req_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [31:0] meipGen_io_in_bridge_io_in_req_bits_addr; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [3:0] meipGen_io_in_bridge_io_in_req_bits_cmd; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [7:0] meipGen_io_in_bridge_io_in_req_bits_wmask; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [63:0] meipGen_io_in_bridge_io_in_req_bits_wdata; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  meipGen_io_in_bridge_io_in_resp_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  meipGen_io_in_bridge_io_in_resp_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [63:0] meipGen_io_in_bridge_io_in_resp_bits_rdata; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  meipGen_io_in_bridge_io_out_aw_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  meipGen_io_in_bridge_io_out_aw_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [31:0] meipGen_io_in_bridge_io_out_aw_bits_addr; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  meipGen_io_in_bridge_io_out_w_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  meipGen_io_in_bridge_io_out_w_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [63:0] meipGen_io_in_bridge_io_out_w_bits_data; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [7:0] meipGen_io_in_bridge_io_out_w_bits_strb; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  meipGen_io_in_bridge_io_out_b_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  meipGen_io_in_bridge_io_out_b_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  meipGen_io_in_bridge_io_out_ar_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  meipGen_io_in_bridge_io_out_ar_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [31:0] meipGen_io_in_bridge_io_out_ar_bits_addr; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  meipGen_io_in_bridge_io_out_r_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  meipGen_io_in_bridge_io_out_r_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [63:0] meipGen_io_in_bridge_io_out_r_bits_data; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  dma_io_in_bridge_clock; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  dma_io_in_bridge_reset; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  dma_io_in_bridge_io_in_req_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  dma_io_in_bridge_io_in_req_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [31:0] dma_io_in_bridge_io_in_req_bits_addr; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [3:0] dma_io_in_bridge_io_in_req_bits_cmd; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [7:0] dma_io_in_bridge_io_in_req_bits_wmask; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [63:0] dma_io_in_bridge_io_in_req_bits_wdata; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  dma_io_in_bridge_io_in_resp_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  dma_io_in_bridge_io_in_resp_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [63:0] dma_io_in_bridge_io_in_resp_bits_rdata; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  dma_io_in_bridge_io_out_aw_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  dma_io_in_bridge_io_out_aw_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [31:0] dma_io_in_bridge_io_out_aw_bits_addr; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  dma_io_in_bridge_io_out_w_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  dma_io_in_bridge_io_out_w_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [63:0] dma_io_in_bridge_io_out_w_bits_data; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [7:0] dma_io_in_bridge_io_out_w_bits_strb; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  dma_io_in_bridge_io_out_b_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  dma_io_in_bridge_io_out_b_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  dma_io_in_bridge_io_out_ar_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  dma_io_in_bridge_io_out_ar_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [31:0] dma_io_in_bridge_io_out_ar_bits_addr; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  dma_io_in_bridge_io_out_r_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  dma_io_in_bridge_io_out_r_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [63:0] dma_io_in_bridge_io_out_r_bits_data; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  SimpleBusCrossbar1toN_1 xbar ( // @[src/main/scala/sim/SimMMIO.scala 45:20]
    .clock(xbar_clock),
    .reset(xbar_reset),
    .io_in_req_ready(xbar_io_in_req_ready),
    .io_in_req_valid(xbar_io_in_req_valid),
    .io_in_req_bits_addr(xbar_io_in_req_bits_addr),
    .io_in_req_bits_size(xbar_io_in_req_bits_size),
    .io_in_req_bits_cmd(xbar_io_in_req_bits_cmd),
    .io_in_req_bits_wmask(xbar_io_in_req_bits_wmask),
    .io_in_req_bits_wdata(xbar_io_in_req_bits_wdata),
    .io_in_resp_ready(xbar_io_in_resp_ready),
    .io_in_resp_valid(xbar_io_in_resp_valid),
    .io_in_resp_bits_cmd(xbar_io_in_resp_bits_cmd),
    .io_in_resp_bits_rdata(xbar_io_in_resp_bits_rdata),
    .io_out_0_req_ready(xbar_io_out_0_req_ready),
    .io_out_0_req_valid(xbar_io_out_0_req_valid),
    .io_out_0_req_bits_addr(xbar_io_out_0_req_bits_addr),
    .io_out_0_req_bits_cmd(xbar_io_out_0_req_bits_cmd),
    .io_out_0_req_bits_wmask(xbar_io_out_0_req_bits_wmask),
    .io_out_0_req_bits_wdata(xbar_io_out_0_req_bits_wdata),
    .io_out_0_resp_ready(xbar_io_out_0_resp_ready),
    .io_out_0_resp_valid(xbar_io_out_0_resp_valid),
    .io_out_0_resp_bits_rdata(xbar_io_out_0_resp_bits_rdata),
    .io_out_1_req_ready(xbar_io_out_1_req_ready),
    .io_out_1_req_valid(xbar_io_out_1_req_valid),
    .io_out_1_req_bits_addr(xbar_io_out_1_req_bits_addr),
    .io_out_1_req_bits_cmd(xbar_io_out_1_req_bits_cmd),
    .io_out_1_req_bits_wmask(xbar_io_out_1_req_bits_wmask),
    .io_out_1_req_bits_wdata(xbar_io_out_1_req_bits_wdata),
    .io_out_1_resp_ready(xbar_io_out_1_resp_ready),
    .io_out_1_resp_valid(xbar_io_out_1_resp_valid),
    .io_out_1_resp_bits_rdata(xbar_io_out_1_resp_bits_rdata),
    .io_out_2_req_ready(xbar_io_out_2_req_ready),
    .io_out_2_req_valid(xbar_io_out_2_req_valid),
    .io_out_2_req_bits_addr(xbar_io_out_2_req_bits_addr),
    .io_out_2_req_bits_cmd(xbar_io_out_2_req_bits_cmd),
    .io_out_2_req_bits_wmask(xbar_io_out_2_req_bits_wmask),
    .io_out_2_req_bits_wdata(xbar_io_out_2_req_bits_wdata),
    .io_out_2_resp_ready(xbar_io_out_2_resp_ready),
    .io_out_2_resp_valid(xbar_io_out_2_resp_valid),
    .io_out_2_resp_bits_rdata(xbar_io_out_2_resp_bits_rdata),
    .io_out_3_req_ready(xbar_io_out_3_req_ready),
    .io_out_3_req_valid(xbar_io_out_3_req_valid),
    .io_out_3_req_bits_addr(xbar_io_out_3_req_bits_addr),
    .io_out_3_req_bits_cmd(xbar_io_out_3_req_bits_cmd),
    .io_out_3_req_bits_wmask(xbar_io_out_3_req_bits_wmask),
    .io_out_3_req_bits_wdata(xbar_io_out_3_req_bits_wdata),
    .io_out_3_resp_ready(xbar_io_out_3_resp_ready),
    .io_out_3_resp_valid(xbar_io_out_3_resp_valid),
    .io_out_3_resp_bits_rdata(xbar_io_out_3_resp_bits_rdata),
    .DISPLAY_ENABLE(xbar_DISPLAY_ENABLE)
  );
  AXI4UART uart ( // @[src/main/scala/sim/SimMMIO.scala 48:20]
    .clock(uart_clock),
    .reset(uart_reset),
    .io_in_aw_ready(uart_io_in_aw_ready),
    .io_in_aw_valid(uart_io_in_aw_valid),
    .io_in_aw_bits_addr(uart_io_in_aw_bits_addr),
    .io_in_w_ready(uart_io_in_w_ready),
    .io_in_w_valid(uart_io_in_w_valid),
    .io_in_w_bits_data(uart_io_in_w_bits_data),
    .io_in_w_bits_strb(uart_io_in_w_bits_strb),
    .io_in_b_ready(uart_io_in_b_ready),
    .io_in_b_valid(uart_io_in_b_valid),
    .io_in_ar_ready(uart_io_in_ar_ready),
    .io_in_ar_valid(uart_io_in_ar_valid),
    .io_in_ar_bits_addr(uart_io_in_ar_bits_addr),
    .io_in_r_ready(uart_io_in_r_ready),
    .io_in_r_valid(uart_io_in_r_valid),
    .io_in_r_bits_data(uart_io_in_r_bits_data),
    .io_extra_out_valid(uart_io_extra_out_valid),
    .io_extra_out_ch(uart_io_extra_out_ch),
    .io_extra_in_valid(uart_io_extra_in_valid),
    .io_extra_in_ch(uart_io_extra_in_ch)
  );
  AXI4Flash flash ( // @[src/main/scala/sim/SimMMIO.scala 50:21]
    .clock(flash_clock),
    .reset(flash_reset),
    .io_in_aw_ready(flash_io_in_aw_ready),
    .io_in_aw_valid(flash_io_in_aw_valid),
    .io_in_w_ready(flash_io_in_w_ready),
    .io_in_w_valid(flash_io_in_w_valid),
    .io_in_b_ready(flash_io_in_b_ready),
    .io_in_b_valid(flash_io_in_b_valid),
    .io_in_ar_ready(flash_io_in_ar_ready),
    .io_in_ar_valid(flash_io_in_ar_valid),
    .io_in_ar_bits_addr(flash_io_in_ar_bits_addr),
    .io_in_r_ready(flash_io_in_r_ready),
    .io_in_r_valid(flash_io_in_r_valid),
    .io_in_r_bits_data(flash_io_in_r_bits_data)
  );
  AXI4MeipGen meipGen ( // @[src/main/scala/sim/SimMMIO.scala 52:23]
    .clock(meipGen_clock),
    .reset(meipGen_reset),
    .io_in_aw_ready(meipGen_io_in_aw_ready),
    .io_in_aw_valid(meipGen_io_in_aw_valid),
    .io_in_aw_bits_addr(meipGen_io_in_aw_bits_addr),
    .io_in_w_ready(meipGen_io_in_w_ready),
    .io_in_w_valid(meipGen_io_in_w_valid),
    .io_in_w_bits_data(meipGen_io_in_w_bits_data),
    .io_in_w_bits_strb(meipGen_io_in_w_bits_strb),
    .io_in_b_ready(meipGen_io_in_b_ready),
    .io_in_b_valid(meipGen_io_in_b_valid),
    .io_in_ar_ready(meipGen_io_in_ar_ready),
    .io_in_ar_valid(meipGen_io_in_ar_valid),
    .io_in_r_ready(meipGen_io_in_r_ready),
    .io_in_r_valid(meipGen_io_in_r_valid),
    .io_in_r_bits_data(meipGen_io_in_r_bits_data),
    .io_extra_meip(meipGen_io_extra_meip)
  );
  AXI4DMA dma ( // @[src/main/scala/sim/SimMMIO.scala 53:19]
    .clock(dma_clock),
    .reset(dma_reset),
    .io_in_aw_ready(dma_io_in_aw_ready),
    .io_in_aw_valid(dma_io_in_aw_valid),
    .io_in_aw_bits_addr(dma_io_in_aw_bits_addr),
    .io_in_w_ready(dma_io_in_w_ready),
    .io_in_w_valid(dma_io_in_w_valid),
    .io_in_w_bits_data(dma_io_in_w_bits_data),
    .io_in_w_bits_strb(dma_io_in_w_bits_strb),
    .io_in_b_ready(dma_io_in_b_ready),
    .io_in_b_valid(dma_io_in_b_valid),
    .io_in_ar_ready(dma_io_in_ar_ready),
    .io_in_ar_valid(dma_io_in_ar_valid),
    .io_in_ar_bits_addr(dma_io_in_ar_bits_addr),
    .io_in_r_ready(dma_io_in_r_ready),
    .io_in_r_valid(dma_io_in_r_valid),
    .io_in_r_bits_data(dma_io_in_r_bits_data),
    .io_extra_dma_aw_ready(dma_io_extra_dma_aw_ready),
    .io_extra_dma_aw_valid(dma_io_extra_dma_aw_valid),
    .io_extra_dma_aw_bits_addr(dma_io_extra_dma_aw_bits_addr),
    .io_extra_dma_aw_bits_len(dma_io_extra_dma_aw_bits_len),
    .io_extra_dma_aw_bits_size(dma_io_extra_dma_aw_bits_size),
    .io_extra_dma_w_ready(dma_io_extra_dma_w_ready),
    .io_extra_dma_w_valid(dma_io_extra_dma_w_valid),
    .io_extra_dma_w_bits_data(dma_io_extra_dma_w_bits_data),
    .io_extra_dma_w_bits_strb(dma_io_extra_dma_w_bits_strb),
    .io_extra_dma_w_bits_last(dma_io_extra_dma_w_bits_last),
    .io_extra_dma_b_ready(dma_io_extra_dma_b_ready),
    .io_extra_dma_b_valid(dma_io_extra_dma_b_valid),
    .io_extra_dma_ar_ready(dma_io_extra_dma_ar_ready),
    .io_extra_dma_ar_valid(dma_io_extra_dma_ar_valid),
    .io_extra_dma_ar_bits_addr(dma_io_extra_dma_ar_bits_addr),
    .io_extra_dma_ar_bits_len(dma_io_extra_dma_ar_bits_len),
    .io_extra_dma_ar_bits_size(dma_io_extra_dma_ar_bits_size),
    .io_extra_dma_r_ready(dma_io_extra_dma_r_ready),
    .io_extra_dma_r_valid(dma_io_extra_dma_r_valid),
    .io_extra_dma_r_bits_data(dma_io_extra_dma_r_bits_data)
  );
  SimpleBus2AXI4Converter_1 uart_io_in_bridge ( // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
    .clock(uart_io_in_bridge_clock),
    .reset(uart_io_in_bridge_reset),
    .io_in_req_ready(uart_io_in_bridge_io_in_req_ready),
    .io_in_req_valid(uart_io_in_bridge_io_in_req_valid),
    .io_in_req_bits_addr(uart_io_in_bridge_io_in_req_bits_addr),
    .io_in_req_bits_cmd(uart_io_in_bridge_io_in_req_bits_cmd),
    .io_in_req_bits_wmask(uart_io_in_bridge_io_in_req_bits_wmask),
    .io_in_req_bits_wdata(uart_io_in_bridge_io_in_req_bits_wdata),
    .io_in_resp_ready(uart_io_in_bridge_io_in_resp_ready),
    .io_in_resp_valid(uart_io_in_bridge_io_in_resp_valid),
    .io_in_resp_bits_rdata(uart_io_in_bridge_io_in_resp_bits_rdata),
    .io_out_aw_ready(uart_io_in_bridge_io_out_aw_ready),
    .io_out_aw_valid(uart_io_in_bridge_io_out_aw_valid),
    .io_out_aw_bits_addr(uart_io_in_bridge_io_out_aw_bits_addr),
    .io_out_w_ready(uart_io_in_bridge_io_out_w_ready),
    .io_out_w_valid(uart_io_in_bridge_io_out_w_valid),
    .io_out_w_bits_data(uart_io_in_bridge_io_out_w_bits_data),
    .io_out_w_bits_strb(uart_io_in_bridge_io_out_w_bits_strb),
    .io_out_b_ready(uart_io_in_bridge_io_out_b_ready),
    .io_out_b_valid(uart_io_in_bridge_io_out_b_valid),
    .io_out_ar_ready(uart_io_in_bridge_io_out_ar_ready),
    .io_out_ar_valid(uart_io_in_bridge_io_out_ar_valid),
    .io_out_ar_bits_addr(uart_io_in_bridge_io_out_ar_bits_addr),
    .io_out_r_ready(uart_io_in_bridge_io_out_r_ready),
    .io_out_r_valid(uart_io_in_bridge_io_out_r_valid),
    .io_out_r_bits_data(uart_io_in_bridge_io_out_r_bits_data)
  );
  SimpleBus2AXI4Converter_1 flash_io_in_bridge ( // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
    .clock(flash_io_in_bridge_clock),
    .reset(flash_io_in_bridge_reset),
    .io_in_req_ready(flash_io_in_bridge_io_in_req_ready),
    .io_in_req_valid(flash_io_in_bridge_io_in_req_valid),
    .io_in_req_bits_addr(flash_io_in_bridge_io_in_req_bits_addr),
    .io_in_req_bits_cmd(flash_io_in_bridge_io_in_req_bits_cmd),
    .io_in_req_bits_wmask(flash_io_in_bridge_io_in_req_bits_wmask),
    .io_in_req_bits_wdata(flash_io_in_bridge_io_in_req_bits_wdata),
    .io_in_resp_ready(flash_io_in_bridge_io_in_resp_ready),
    .io_in_resp_valid(flash_io_in_bridge_io_in_resp_valid),
    .io_in_resp_bits_rdata(flash_io_in_bridge_io_in_resp_bits_rdata),
    .io_out_aw_ready(flash_io_in_bridge_io_out_aw_ready),
    .io_out_aw_valid(flash_io_in_bridge_io_out_aw_valid),
    .io_out_aw_bits_addr(flash_io_in_bridge_io_out_aw_bits_addr),
    .io_out_w_ready(flash_io_in_bridge_io_out_w_ready),
    .io_out_w_valid(flash_io_in_bridge_io_out_w_valid),
    .io_out_w_bits_data(flash_io_in_bridge_io_out_w_bits_data),
    .io_out_w_bits_strb(flash_io_in_bridge_io_out_w_bits_strb),
    .io_out_b_ready(flash_io_in_bridge_io_out_b_ready),
    .io_out_b_valid(flash_io_in_bridge_io_out_b_valid),
    .io_out_ar_ready(flash_io_in_bridge_io_out_ar_ready),
    .io_out_ar_valid(flash_io_in_bridge_io_out_ar_valid),
    .io_out_ar_bits_addr(flash_io_in_bridge_io_out_ar_bits_addr),
    .io_out_r_ready(flash_io_in_bridge_io_out_r_ready),
    .io_out_r_valid(flash_io_in_bridge_io_out_r_valid),
    .io_out_r_bits_data(flash_io_in_bridge_io_out_r_bits_data)
  );
  SimpleBus2AXI4Converter_1 meipGen_io_in_bridge ( // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
    .clock(meipGen_io_in_bridge_clock),
    .reset(meipGen_io_in_bridge_reset),
    .io_in_req_ready(meipGen_io_in_bridge_io_in_req_ready),
    .io_in_req_valid(meipGen_io_in_bridge_io_in_req_valid),
    .io_in_req_bits_addr(meipGen_io_in_bridge_io_in_req_bits_addr),
    .io_in_req_bits_cmd(meipGen_io_in_bridge_io_in_req_bits_cmd),
    .io_in_req_bits_wmask(meipGen_io_in_bridge_io_in_req_bits_wmask),
    .io_in_req_bits_wdata(meipGen_io_in_bridge_io_in_req_bits_wdata),
    .io_in_resp_ready(meipGen_io_in_bridge_io_in_resp_ready),
    .io_in_resp_valid(meipGen_io_in_bridge_io_in_resp_valid),
    .io_in_resp_bits_rdata(meipGen_io_in_bridge_io_in_resp_bits_rdata),
    .io_out_aw_ready(meipGen_io_in_bridge_io_out_aw_ready),
    .io_out_aw_valid(meipGen_io_in_bridge_io_out_aw_valid),
    .io_out_aw_bits_addr(meipGen_io_in_bridge_io_out_aw_bits_addr),
    .io_out_w_ready(meipGen_io_in_bridge_io_out_w_ready),
    .io_out_w_valid(meipGen_io_in_bridge_io_out_w_valid),
    .io_out_w_bits_data(meipGen_io_in_bridge_io_out_w_bits_data),
    .io_out_w_bits_strb(meipGen_io_in_bridge_io_out_w_bits_strb),
    .io_out_b_ready(meipGen_io_in_bridge_io_out_b_ready),
    .io_out_b_valid(meipGen_io_in_bridge_io_out_b_valid),
    .io_out_ar_ready(meipGen_io_in_bridge_io_out_ar_ready),
    .io_out_ar_valid(meipGen_io_in_bridge_io_out_ar_valid),
    .io_out_ar_bits_addr(meipGen_io_in_bridge_io_out_ar_bits_addr),
    .io_out_r_ready(meipGen_io_in_bridge_io_out_r_ready),
    .io_out_r_valid(meipGen_io_in_bridge_io_out_r_valid),
    .io_out_r_bits_data(meipGen_io_in_bridge_io_out_r_bits_data)
  );
  SimpleBus2AXI4Converter_1 dma_io_in_bridge ( // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
    .clock(dma_io_in_bridge_clock),
    .reset(dma_io_in_bridge_reset),
    .io_in_req_ready(dma_io_in_bridge_io_in_req_ready),
    .io_in_req_valid(dma_io_in_bridge_io_in_req_valid),
    .io_in_req_bits_addr(dma_io_in_bridge_io_in_req_bits_addr),
    .io_in_req_bits_cmd(dma_io_in_bridge_io_in_req_bits_cmd),
    .io_in_req_bits_wmask(dma_io_in_bridge_io_in_req_bits_wmask),
    .io_in_req_bits_wdata(dma_io_in_bridge_io_in_req_bits_wdata),
    .io_in_resp_ready(dma_io_in_bridge_io_in_resp_ready),
    .io_in_resp_valid(dma_io_in_bridge_io_in_resp_valid),
    .io_in_resp_bits_rdata(dma_io_in_bridge_io_in_resp_bits_rdata),
    .io_out_aw_ready(dma_io_in_bridge_io_out_aw_ready),
    .io_out_aw_valid(dma_io_in_bridge_io_out_aw_valid),
    .io_out_aw_bits_addr(dma_io_in_bridge_io_out_aw_bits_addr),
    .io_out_w_ready(dma_io_in_bridge_io_out_w_ready),
    .io_out_w_valid(dma_io_in_bridge_io_out_w_valid),
    .io_out_w_bits_data(dma_io_in_bridge_io_out_w_bits_data),
    .io_out_w_bits_strb(dma_io_in_bridge_io_out_w_bits_strb),
    .io_out_b_ready(dma_io_in_bridge_io_out_b_ready),
    .io_out_b_valid(dma_io_in_bridge_io_out_b_valid),
    .io_out_ar_ready(dma_io_in_bridge_io_out_ar_ready),
    .io_out_ar_valid(dma_io_in_bridge_io_out_ar_valid),
    .io_out_ar_bits_addr(dma_io_in_bridge_io_out_ar_bits_addr),
    .io_out_r_ready(dma_io_in_bridge_io_out_r_ready),
    .io_out_r_valid(dma_io_in_bridge_io_out_r_valid),
    .io_out_r_bits_data(dma_io_in_bridge_io_out_r_bits_data)
  );
  assign io_rw_req_ready = xbar_io_in_req_ready; // @[src/main/scala/sim/SimMMIO.scala 46:14]
  assign io_rw_resp_valid = xbar_io_in_resp_valid; // @[src/main/scala/sim/SimMMIO.scala 46:14]
  assign io_rw_resp_bits_cmd = xbar_io_in_resp_bits_cmd; // @[src/main/scala/sim/SimMMIO.scala 46:14]
  assign io_rw_resp_bits_rdata = xbar_io_in_resp_bits_rdata; // @[src/main/scala/sim/SimMMIO.scala 46:14]
  assign io_meip = meipGen_io_extra_meip; // @[src/main/scala/sim/SimMMIO.scala 62:11]
  assign io_dma_aw_valid = dma_io_extra_dma_aw_valid; // @[src/main/scala/sim/SimMMIO.scala 61:10]
  assign io_dma_aw_bits_addr = dma_io_extra_dma_aw_bits_addr; // @[src/main/scala/sim/SimMMIO.scala 61:10]
  assign io_dma_aw_bits_len = dma_io_extra_dma_aw_bits_len; // @[src/main/scala/sim/SimMMIO.scala 61:10]
  assign io_dma_aw_bits_size = dma_io_extra_dma_aw_bits_size; // @[src/main/scala/sim/SimMMIO.scala 61:10]
  assign io_dma_w_valid = dma_io_extra_dma_w_valid; // @[src/main/scala/sim/SimMMIO.scala 61:10]
  assign io_dma_w_bits_data = dma_io_extra_dma_w_bits_data; // @[src/main/scala/sim/SimMMIO.scala 61:10]
  assign io_dma_w_bits_strb = dma_io_extra_dma_w_bits_strb; // @[src/main/scala/sim/SimMMIO.scala 61:10]
  assign io_dma_b_ready = dma_io_extra_dma_b_ready; // @[src/main/scala/sim/SimMMIO.scala 61:10]
  assign io_dma_ar_valid = dma_io_extra_dma_ar_valid; // @[src/main/scala/sim/SimMMIO.scala 61:10]
  assign io_dma_ar_bits_addr = dma_io_extra_dma_ar_bits_addr; // @[src/main/scala/sim/SimMMIO.scala 61:10]
  assign io_dma_r_ready = dma_io_extra_dma_r_ready; // @[src/main/scala/sim/SimMMIO.scala 61:10]
  assign io_uart_out_valid = uart_io_extra_out_valid; // @[src/main/scala/sim/SimMMIO.scala 63:21]
  assign io_uart_out_ch = uart_io_extra_out_ch; // @[src/main/scala/sim/SimMMIO.scala 63:21]
  assign io_uart_in_valid = uart_io_extra_in_valid; // @[src/main/scala/sim/SimMMIO.scala 63:21]
  assign xbar_clock = clock;
  assign xbar_reset = reset;
  assign xbar_io_in_req_valid = io_rw_req_valid; // @[src/main/scala/sim/SimMMIO.scala 46:14]
  assign xbar_io_in_req_bits_addr = io_rw_req_bits_addr; // @[src/main/scala/sim/SimMMIO.scala 46:14]
  assign xbar_io_in_req_bits_size = io_rw_req_bits_size; // @[src/main/scala/sim/SimMMIO.scala 46:14]
  assign xbar_io_in_req_bits_cmd = io_rw_req_bits_cmd; // @[src/main/scala/sim/SimMMIO.scala 46:14]
  assign xbar_io_in_req_bits_wmask = io_rw_req_bits_wmask; // @[src/main/scala/sim/SimMMIO.scala 46:14]
  assign xbar_io_in_req_bits_wdata = io_rw_req_bits_wdata; // @[src/main/scala/sim/SimMMIO.scala 46:14]
  assign xbar_io_in_resp_ready = io_rw_resp_ready; // @[src/main/scala/sim/SimMMIO.scala 46:14]
  assign xbar_io_out_0_req_ready = uart_io_in_bridge_io_in_req_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign xbar_io_out_0_resp_valid = uart_io_in_bridge_io_in_resp_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign xbar_io_out_0_resp_bits_rdata = uart_io_in_bridge_io_in_resp_bits_rdata; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign xbar_io_out_1_req_ready = flash_io_in_bridge_io_in_req_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign xbar_io_out_1_resp_valid = flash_io_in_bridge_io_in_resp_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign xbar_io_out_1_resp_bits_rdata = flash_io_in_bridge_io_in_resp_bits_rdata; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign xbar_io_out_2_req_ready = meipGen_io_in_bridge_io_in_req_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign xbar_io_out_2_resp_valid = meipGen_io_in_bridge_io_in_resp_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign xbar_io_out_2_resp_bits_rdata = meipGen_io_in_bridge_io_in_resp_bits_rdata; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign xbar_io_out_3_req_ready = dma_io_in_bridge_io_in_req_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign xbar_io_out_3_resp_valid = dma_io_in_bridge_io_in_resp_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign xbar_io_out_3_resp_bits_rdata = dma_io_in_bridge_io_in_resp_bits_rdata; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign xbar_DISPLAY_ENABLE = _WIRE_4;
  assign uart_clock = clock;
  assign uart_reset = reset;
  assign uart_io_in_aw_valid = uart_io_in_bridge_io_out_aw_valid; // @[src/main/scala/sim/SimMMIO.scala 54:14]
  assign uart_io_in_aw_bits_addr = uart_io_in_bridge_io_out_aw_bits_addr; // @[src/main/scala/sim/SimMMIO.scala 54:14]
  assign uart_io_in_w_valid = uart_io_in_bridge_io_out_w_valid; // @[src/main/scala/sim/SimMMIO.scala 54:14]
  assign uart_io_in_w_bits_data = uart_io_in_bridge_io_out_w_bits_data; // @[src/main/scala/sim/SimMMIO.scala 54:14]
  assign uart_io_in_w_bits_strb = uart_io_in_bridge_io_out_w_bits_strb; // @[src/main/scala/sim/SimMMIO.scala 54:14]
  assign uart_io_in_b_ready = uart_io_in_bridge_io_out_b_ready; // @[src/main/scala/sim/SimMMIO.scala 54:14]
  assign uart_io_in_ar_valid = uart_io_in_bridge_io_out_ar_valid; // @[src/main/scala/sim/SimMMIO.scala 54:14]
  assign uart_io_in_ar_bits_addr = uart_io_in_bridge_io_out_ar_bits_addr; // @[src/main/scala/sim/SimMMIO.scala 54:14]
  assign uart_io_in_r_ready = uart_io_in_bridge_io_out_r_ready; // @[src/main/scala/sim/SimMMIO.scala 54:14]
  assign uart_io_extra_in_ch = io_uart_in_ch; // @[src/main/scala/sim/SimMMIO.scala 63:21]
  assign flash_clock = clock;
  assign flash_reset = reset;
  assign flash_io_in_aw_valid = flash_io_in_bridge_io_out_aw_valid; // @[src/main/scala/sim/SimMMIO.scala 57:15]
  assign flash_io_in_w_valid = flash_io_in_bridge_io_out_w_valid; // @[src/main/scala/sim/SimMMIO.scala 57:15]
  assign flash_io_in_b_ready = flash_io_in_bridge_io_out_b_ready; // @[src/main/scala/sim/SimMMIO.scala 57:15]
  assign flash_io_in_ar_valid = flash_io_in_bridge_io_out_ar_valid; // @[src/main/scala/sim/SimMMIO.scala 57:15]
  assign flash_io_in_ar_bits_addr = flash_io_in_bridge_io_out_ar_bits_addr; // @[src/main/scala/sim/SimMMIO.scala 57:15]
  assign flash_io_in_r_ready = flash_io_in_bridge_io_out_r_ready; // @[src/main/scala/sim/SimMMIO.scala 57:15]
  assign meipGen_clock = clock;
  assign meipGen_reset = reset;
  assign meipGen_io_in_aw_valid = meipGen_io_in_bridge_io_out_aw_valid; // @[src/main/scala/sim/SimMMIO.scala 59:17]
  assign meipGen_io_in_aw_bits_addr = meipGen_io_in_bridge_io_out_aw_bits_addr; // @[src/main/scala/sim/SimMMIO.scala 59:17]
  assign meipGen_io_in_w_valid = meipGen_io_in_bridge_io_out_w_valid; // @[src/main/scala/sim/SimMMIO.scala 59:17]
  assign meipGen_io_in_w_bits_data = meipGen_io_in_bridge_io_out_w_bits_data; // @[src/main/scala/sim/SimMMIO.scala 59:17]
  assign meipGen_io_in_w_bits_strb = meipGen_io_in_bridge_io_out_w_bits_strb; // @[src/main/scala/sim/SimMMIO.scala 59:17]
  assign meipGen_io_in_b_ready = meipGen_io_in_bridge_io_out_b_ready; // @[src/main/scala/sim/SimMMIO.scala 59:17]
  assign meipGen_io_in_ar_valid = meipGen_io_in_bridge_io_out_ar_valid; // @[src/main/scala/sim/SimMMIO.scala 59:17]
  assign meipGen_io_in_r_ready = meipGen_io_in_bridge_io_out_r_ready; // @[src/main/scala/sim/SimMMIO.scala 59:17]
  assign dma_clock = clock;
  assign dma_reset = reset;
  assign dma_io_in_aw_valid = dma_io_in_bridge_io_out_aw_valid; // @[src/main/scala/sim/SimMMIO.scala 60:13]
  assign dma_io_in_aw_bits_addr = dma_io_in_bridge_io_out_aw_bits_addr; // @[src/main/scala/sim/SimMMIO.scala 60:13]
  assign dma_io_in_w_valid = dma_io_in_bridge_io_out_w_valid; // @[src/main/scala/sim/SimMMIO.scala 60:13]
  assign dma_io_in_w_bits_data = dma_io_in_bridge_io_out_w_bits_data; // @[src/main/scala/sim/SimMMIO.scala 60:13]
  assign dma_io_in_w_bits_strb = dma_io_in_bridge_io_out_w_bits_strb; // @[src/main/scala/sim/SimMMIO.scala 60:13]
  assign dma_io_in_b_ready = dma_io_in_bridge_io_out_b_ready; // @[src/main/scala/sim/SimMMIO.scala 60:13]
  assign dma_io_in_ar_valid = dma_io_in_bridge_io_out_ar_valid; // @[src/main/scala/sim/SimMMIO.scala 60:13]
  assign dma_io_in_ar_bits_addr = dma_io_in_bridge_io_out_ar_bits_addr; // @[src/main/scala/sim/SimMMIO.scala 60:13]
  assign dma_io_in_r_ready = dma_io_in_bridge_io_out_r_ready; // @[src/main/scala/sim/SimMMIO.scala 60:13]
  assign dma_io_extra_dma_aw_ready = io_dma_aw_ready; // @[src/main/scala/sim/SimMMIO.scala 61:10]
  assign dma_io_extra_dma_w_ready = io_dma_w_ready; // @[src/main/scala/sim/SimMMIO.scala 61:10]
  assign dma_io_extra_dma_b_valid = io_dma_b_valid; // @[src/main/scala/sim/SimMMIO.scala 61:10]
  assign dma_io_extra_dma_ar_ready = io_dma_ar_ready; // @[src/main/scala/sim/SimMMIO.scala 61:10]
  assign dma_io_extra_dma_r_valid = io_dma_r_valid; // @[src/main/scala/sim/SimMMIO.scala 61:10]
  assign dma_io_extra_dma_r_bits_data = io_dma_r_bits_data; // @[src/main/scala/sim/SimMMIO.scala 61:10]
  assign uart_io_in_bridge_clock = clock;
  assign uart_io_in_bridge_reset = reset;
  assign uart_io_in_bridge_io_in_req_valid = xbar_io_out_0_req_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign uart_io_in_bridge_io_in_req_bits_addr = xbar_io_out_0_req_bits_addr; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign uart_io_in_bridge_io_in_req_bits_cmd = xbar_io_out_0_req_bits_cmd; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign uart_io_in_bridge_io_in_req_bits_wmask = xbar_io_out_0_req_bits_wmask; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign uart_io_in_bridge_io_in_req_bits_wdata = xbar_io_out_0_req_bits_wdata; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign uart_io_in_bridge_io_in_resp_ready = xbar_io_out_0_resp_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign uart_io_in_bridge_io_out_aw_ready = uart_io_in_aw_ready; // @[src/main/scala/sim/SimMMIO.scala 54:14]
  assign uart_io_in_bridge_io_out_w_ready = uart_io_in_w_ready; // @[src/main/scala/sim/SimMMIO.scala 54:14]
  assign uart_io_in_bridge_io_out_b_valid = uart_io_in_b_valid; // @[src/main/scala/sim/SimMMIO.scala 54:14]
  assign uart_io_in_bridge_io_out_ar_ready = uart_io_in_ar_ready; // @[src/main/scala/sim/SimMMIO.scala 54:14]
  assign uart_io_in_bridge_io_out_r_valid = uart_io_in_r_valid; // @[src/main/scala/sim/SimMMIO.scala 54:14]
  assign uart_io_in_bridge_io_out_r_bits_data = uart_io_in_r_bits_data; // @[src/main/scala/sim/SimMMIO.scala 54:14]
  assign flash_io_in_bridge_clock = clock;
  assign flash_io_in_bridge_reset = reset;
  assign flash_io_in_bridge_io_in_req_valid = xbar_io_out_1_req_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign flash_io_in_bridge_io_in_req_bits_addr = xbar_io_out_1_req_bits_addr; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign flash_io_in_bridge_io_in_req_bits_cmd = xbar_io_out_1_req_bits_cmd; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign flash_io_in_bridge_io_in_req_bits_wmask = xbar_io_out_1_req_bits_wmask; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign flash_io_in_bridge_io_in_req_bits_wdata = xbar_io_out_1_req_bits_wdata; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign flash_io_in_bridge_io_in_resp_ready = xbar_io_out_1_resp_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign flash_io_in_bridge_io_out_aw_ready = flash_io_in_aw_ready; // @[src/main/scala/sim/SimMMIO.scala 57:15]
  assign flash_io_in_bridge_io_out_w_ready = flash_io_in_w_ready; // @[src/main/scala/sim/SimMMIO.scala 57:15]
  assign flash_io_in_bridge_io_out_b_valid = flash_io_in_b_valid; // @[src/main/scala/sim/SimMMIO.scala 57:15]
  assign flash_io_in_bridge_io_out_ar_ready = flash_io_in_ar_ready; // @[src/main/scala/sim/SimMMIO.scala 57:15]
  assign flash_io_in_bridge_io_out_r_valid = flash_io_in_r_valid; // @[src/main/scala/sim/SimMMIO.scala 57:15]
  assign flash_io_in_bridge_io_out_r_bits_data = flash_io_in_r_bits_data; // @[src/main/scala/sim/SimMMIO.scala 57:15]
  assign meipGen_io_in_bridge_clock = clock;
  assign meipGen_io_in_bridge_reset = reset;
  assign meipGen_io_in_bridge_io_in_req_valid = xbar_io_out_2_req_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign meipGen_io_in_bridge_io_in_req_bits_addr = xbar_io_out_2_req_bits_addr; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign meipGen_io_in_bridge_io_in_req_bits_cmd = xbar_io_out_2_req_bits_cmd; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign meipGen_io_in_bridge_io_in_req_bits_wmask = xbar_io_out_2_req_bits_wmask; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign meipGen_io_in_bridge_io_in_req_bits_wdata = xbar_io_out_2_req_bits_wdata; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign meipGen_io_in_bridge_io_in_resp_ready = xbar_io_out_2_resp_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign meipGen_io_in_bridge_io_out_aw_ready = meipGen_io_in_aw_ready; // @[src/main/scala/sim/SimMMIO.scala 59:17]
  assign meipGen_io_in_bridge_io_out_w_ready = meipGen_io_in_w_ready; // @[src/main/scala/sim/SimMMIO.scala 59:17]
  assign meipGen_io_in_bridge_io_out_b_valid = meipGen_io_in_b_valid; // @[src/main/scala/sim/SimMMIO.scala 59:17]
  assign meipGen_io_in_bridge_io_out_ar_ready = meipGen_io_in_ar_ready; // @[src/main/scala/sim/SimMMIO.scala 59:17]
  assign meipGen_io_in_bridge_io_out_r_valid = meipGen_io_in_r_valid; // @[src/main/scala/sim/SimMMIO.scala 59:17]
  assign meipGen_io_in_bridge_io_out_r_bits_data = meipGen_io_in_r_bits_data; // @[src/main/scala/sim/SimMMIO.scala 59:17]
  assign dma_io_in_bridge_clock = clock;
  assign dma_io_in_bridge_reset = reset;
  assign dma_io_in_bridge_io_in_req_valid = xbar_io_out_3_req_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign dma_io_in_bridge_io_in_req_bits_addr = xbar_io_out_3_req_bits_addr; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign dma_io_in_bridge_io_in_req_bits_cmd = xbar_io_out_3_req_bits_cmd; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign dma_io_in_bridge_io_in_req_bits_wmask = xbar_io_out_3_req_bits_wmask; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign dma_io_in_bridge_io_in_req_bits_wdata = xbar_io_out_3_req_bits_wdata; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign dma_io_in_bridge_io_in_resp_ready = xbar_io_out_3_resp_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign dma_io_in_bridge_io_out_aw_ready = dma_io_in_aw_ready; // @[src/main/scala/sim/SimMMIO.scala 60:13]
  assign dma_io_in_bridge_io_out_w_ready = dma_io_in_w_ready; // @[src/main/scala/sim/SimMMIO.scala 60:13]
  assign dma_io_in_bridge_io_out_b_valid = dma_io_in_b_valid; // @[src/main/scala/sim/SimMMIO.scala 60:13]
  assign dma_io_in_bridge_io_out_ar_ready = dma_io_in_ar_ready; // @[src/main/scala/sim/SimMMIO.scala 60:13]
  assign dma_io_in_bridge_io_out_r_valid = dma_io_in_r_valid; // @[src/main/scala/sim/SimMMIO.scala 60:13]
  assign dma_io_in_bridge_io_out_r_bits_data = dma_io_in_r_bits_data; // @[src/main/scala/sim/SimMMIO.scala 60:13]
endmodule
module SimTop(
  input         clock,
  input         reset,
  input  [63:0] io_logCtrl_log_begin, // @[src/main/scala/sim/NutShellSim.scala 33:14]
  input  [63:0] io_logCtrl_log_end, // @[src/main/scala/sim/NutShellSim.scala 33:14]
  input  [63:0] io_logCtrl_log_level, // @[src/main/scala/sim/NutShellSim.scala 33:14]
  input         io_perfInfo_clean, // @[src/main/scala/sim/NutShellSim.scala 33:14]
  input         io_perfInfo_dump, // @[src/main/scala/sim/NutShellSim.scala 33:14]
  output        io_uart_out_valid, // @[src/main/scala/sim/NutShellSim.scala 33:14]
  output [7:0]  io_uart_out_ch, // @[src/main/scala/sim/NutShellSim.scala 33:14]
  output        io_uart_in_valid, // @[src/main/scala/sim/NutShellSim.scala 33:14]
  input  [7:0]  io_uart_in_ch, // @[src/main/scala/sim/NutShellSim.scala 33:14]
  output        difftest_step // @[difftest/src/main/scala/Difftest.scala 310:27]
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  wire  soc_clock; // @[src/main/scala/sim/NutShellSim.scala 40:19]
  wire  soc_reset; // @[src/main/scala/sim/NutShellSim.scala 40:19]
  wire  soc_io_mem_aw_ready; // @[src/main/scala/sim/NutShellSim.scala 40:19]
  wire  soc_io_mem_aw_valid; // @[src/main/scala/sim/NutShellSim.scala 40:19]
  wire [31:0] soc_io_mem_aw_bits_addr; // @[src/main/scala/sim/NutShellSim.scala 40:19]
  wire [7:0] soc_io_mem_aw_bits_len; // @[src/main/scala/sim/NutShellSim.scala 40:19]
  wire [2:0] soc_io_mem_aw_bits_size; // @[src/main/scala/sim/NutShellSim.scala 40:19]
  wire [1:0] soc_io_mem_aw_bits_burst; // @[src/main/scala/sim/NutShellSim.scala 40:19]
  wire  soc_io_mem_w_ready; // @[src/main/scala/sim/NutShellSim.scala 40:19]
  wire  soc_io_mem_w_valid; // @[src/main/scala/sim/NutShellSim.scala 40:19]
  wire [63:0] soc_io_mem_w_bits_data; // @[src/main/scala/sim/NutShellSim.scala 40:19]
  wire  soc_io_mem_w_bits_last; // @[src/main/scala/sim/NutShellSim.scala 40:19]
  wire  soc_io_mem_b_valid; // @[src/main/scala/sim/NutShellSim.scala 40:19]
  wire  soc_io_mem_ar_ready; // @[src/main/scala/sim/NutShellSim.scala 40:19]
  wire  soc_io_mem_ar_valid; // @[src/main/scala/sim/NutShellSim.scala 40:19]
  wire [31:0] soc_io_mem_ar_bits_addr; // @[src/main/scala/sim/NutShellSim.scala 40:19]
  wire [7:0] soc_io_mem_ar_bits_len; // @[src/main/scala/sim/NutShellSim.scala 40:19]
  wire  soc_io_mem_r_valid; // @[src/main/scala/sim/NutShellSim.scala 40:19]
  wire [63:0] soc_io_mem_r_bits_data; // @[src/main/scala/sim/NutShellSim.scala 40:19]
  wire  soc_io_mem_r_bits_last; // @[src/main/scala/sim/NutShellSim.scala 40:19]
  wire  soc_io_mmio_req_ready; // @[src/main/scala/sim/NutShellSim.scala 40:19]
  wire  soc_io_mmio_req_valid; // @[src/main/scala/sim/NutShellSim.scala 40:19]
  wire [31:0] soc_io_mmio_req_bits_addr; // @[src/main/scala/sim/NutShellSim.scala 40:19]
  wire [2:0] soc_io_mmio_req_bits_size; // @[src/main/scala/sim/NutShellSim.scala 40:19]
  wire [3:0] soc_io_mmio_req_bits_cmd; // @[src/main/scala/sim/NutShellSim.scala 40:19]
  wire [7:0] soc_io_mmio_req_bits_wmask; // @[src/main/scala/sim/NutShellSim.scala 40:19]
  wire [63:0] soc_io_mmio_req_bits_wdata; // @[src/main/scala/sim/NutShellSim.scala 40:19]
  wire  soc_io_mmio_resp_ready; // @[src/main/scala/sim/NutShellSim.scala 40:19]
  wire  soc_io_mmio_resp_valid; // @[src/main/scala/sim/NutShellSim.scala 40:19]
  wire [3:0] soc_io_mmio_resp_bits_cmd; // @[src/main/scala/sim/NutShellSim.scala 40:19]
  wire [63:0] soc_io_mmio_resp_bits_rdata; // @[src/main/scala/sim/NutShellSim.scala 40:19]
  wire  soc_io_frontend_aw_ready; // @[src/main/scala/sim/NutShellSim.scala 40:19]
  wire  soc_io_frontend_aw_valid; // @[src/main/scala/sim/NutShellSim.scala 40:19]
  wire [31:0] soc_io_frontend_aw_bits_addr; // @[src/main/scala/sim/NutShellSim.scala 40:19]
  wire [7:0] soc_io_frontend_aw_bits_len; // @[src/main/scala/sim/NutShellSim.scala 40:19]
  wire [2:0] soc_io_frontend_aw_bits_size; // @[src/main/scala/sim/NutShellSim.scala 40:19]
  wire  soc_io_frontend_w_ready; // @[src/main/scala/sim/NutShellSim.scala 40:19]
  wire  soc_io_frontend_w_valid; // @[src/main/scala/sim/NutShellSim.scala 40:19]
  wire [63:0] soc_io_frontend_w_bits_data; // @[src/main/scala/sim/NutShellSim.scala 40:19]
  wire [7:0] soc_io_frontend_w_bits_strb; // @[src/main/scala/sim/NutShellSim.scala 40:19]
  wire  soc_io_frontend_b_ready; // @[src/main/scala/sim/NutShellSim.scala 40:19]
  wire  soc_io_frontend_b_valid; // @[src/main/scala/sim/NutShellSim.scala 40:19]
  wire  soc_io_frontend_ar_ready; // @[src/main/scala/sim/NutShellSim.scala 40:19]
  wire  soc_io_frontend_ar_valid; // @[src/main/scala/sim/NutShellSim.scala 40:19]
  wire [31:0] soc_io_frontend_ar_bits_addr; // @[src/main/scala/sim/NutShellSim.scala 40:19]
  wire  soc_io_frontend_r_ready; // @[src/main/scala/sim/NutShellSim.scala 40:19]
  wire  soc_io_frontend_r_valid; // @[src/main/scala/sim/NutShellSim.scala 40:19]
  wire [63:0] soc_io_frontend_r_bits_data; // @[src/main/scala/sim/NutShellSim.scala 40:19]
  wire  soc_io_meip; // @[src/main/scala/sim/NutShellSim.scala 40:19]
  wire  soc__WIRE_4; // @[src/main/scala/sim/NutShellSim.scala 40:19]
  wire  mem_clock; // @[src/main/scala/sim/NutShellSim.scala 41:19]
  wire  mem_reset; // @[src/main/scala/sim/NutShellSim.scala 41:19]
  wire  mem_io_in_aw_ready; // @[src/main/scala/sim/NutShellSim.scala 41:19]
  wire  mem_io_in_aw_valid; // @[src/main/scala/sim/NutShellSim.scala 41:19]
  wire [31:0] mem_io_in_aw_bits_addr; // @[src/main/scala/sim/NutShellSim.scala 41:19]
  wire  mem_io_in_w_ready; // @[src/main/scala/sim/NutShellSim.scala 41:19]
  wire  mem_io_in_w_valid; // @[src/main/scala/sim/NutShellSim.scala 41:19]
  wire [63:0] mem_io_in_w_bits_data; // @[src/main/scala/sim/NutShellSim.scala 41:19]
  wire  mem_io_in_w_bits_last; // @[src/main/scala/sim/NutShellSim.scala 41:19]
  wire  mem_io_in_b_valid; // @[src/main/scala/sim/NutShellSim.scala 41:19]
  wire  mem_io_in_ar_ready; // @[src/main/scala/sim/NutShellSim.scala 41:19]
  wire  mem_io_in_ar_valid; // @[src/main/scala/sim/NutShellSim.scala 41:19]
  wire [31:0] mem_io_in_ar_bits_addr; // @[src/main/scala/sim/NutShellSim.scala 41:19]
  wire [7:0] mem_io_in_ar_bits_len; // @[src/main/scala/sim/NutShellSim.scala 41:19]
  wire [2:0] mem_io_in_ar_bits_size; // @[src/main/scala/sim/NutShellSim.scala 41:19]
  wire [1:0] mem_io_in_ar_bits_burst; // @[src/main/scala/sim/NutShellSim.scala 41:19]
  wire  mem_io_in_r_valid; // @[src/main/scala/sim/NutShellSim.scala 41:19]
  wire [63:0] mem_io_in_r_bits_data; // @[src/main/scala/sim/NutShellSim.scala 41:19]
  wire  mem_io_in_r_bits_last; // @[src/main/scala/sim/NutShellSim.scala 41:19]
  wire  memdelay_io_in_aw_ready; // @[src/main/scala/sim/NutShellSim.scala 44:24]
  wire  memdelay_io_in_aw_valid; // @[src/main/scala/sim/NutShellSim.scala 44:24]
  wire [31:0] memdelay_io_in_aw_bits_addr; // @[src/main/scala/sim/NutShellSim.scala 44:24]
  wire [7:0] memdelay_io_in_aw_bits_len; // @[src/main/scala/sim/NutShellSim.scala 44:24]
  wire [2:0] memdelay_io_in_aw_bits_size; // @[src/main/scala/sim/NutShellSim.scala 44:24]
  wire [1:0] memdelay_io_in_aw_bits_burst; // @[src/main/scala/sim/NutShellSim.scala 44:24]
  wire  memdelay_io_in_w_ready; // @[src/main/scala/sim/NutShellSim.scala 44:24]
  wire  memdelay_io_in_w_valid; // @[src/main/scala/sim/NutShellSim.scala 44:24]
  wire [63:0] memdelay_io_in_w_bits_data; // @[src/main/scala/sim/NutShellSim.scala 44:24]
  wire  memdelay_io_in_w_bits_last; // @[src/main/scala/sim/NutShellSim.scala 44:24]
  wire  memdelay_io_in_b_valid; // @[src/main/scala/sim/NutShellSim.scala 44:24]
  wire  memdelay_io_in_ar_ready; // @[src/main/scala/sim/NutShellSim.scala 44:24]
  wire  memdelay_io_in_ar_valid; // @[src/main/scala/sim/NutShellSim.scala 44:24]
  wire [31:0] memdelay_io_in_ar_bits_addr; // @[src/main/scala/sim/NutShellSim.scala 44:24]
  wire [7:0] memdelay_io_in_ar_bits_len; // @[src/main/scala/sim/NutShellSim.scala 44:24]
  wire  memdelay_io_in_r_valid; // @[src/main/scala/sim/NutShellSim.scala 44:24]
  wire [63:0] memdelay_io_in_r_bits_data; // @[src/main/scala/sim/NutShellSim.scala 44:24]
  wire  memdelay_io_in_r_bits_last; // @[src/main/scala/sim/NutShellSim.scala 44:24]
  wire  memdelay_io_out_aw_ready; // @[src/main/scala/sim/NutShellSim.scala 44:24]
  wire  memdelay_io_out_aw_valid; // @[src/main/scala/sim/NutShellSim.scala 44:24]
  wire [31:0] memdelay_io_out_aw_bits_addr; // @[src/main/scala/sim/NutShellSim.scala 44:24]
  wire  memdelay_io_out_w_ready; // @[src/main/scala/sim/NutShellSim.scala 44:24]
  wire  memdelay_io_out_w_valid; // @[src/main/scala/sim/NutShellSim.scala 44:24]
  wire [63:0] memdelay_io_out_w_bits_data; // @[src/main/scala/sim/NutShellSim.scala 44:24]
  wire  memdelay_io_out_w_bits_last; // @[src/main/scala/sim/NutShellSim.scala 44:24]
  wire  memdelay_io_out_b_valid; // @[src/main/scala/sim/NutShellSim.scala 44:24]
  wire  memdelay_io_out_ar_valid; // @[src/main/scala/sim/NutShellSim.scala 44:24]
  wire [31:0] memdelay_io_out_ar_bits_addr; // @[src/main/scala/sim/NutShellSim.scala 44:24]
  wire [7:0] memdelay_io_out_ar_bits_len; // @[src/main/scala/sim/NutShellSim.scala 44:24]
  wire [2:0] memdelay_io_out_ar_bits_size; // @[src/main/scala/sim/NutShellSim.scala 44:24]
  wire [1:0] memdelay_io_out_ar_bits_burst; // @[src/main/scala/sim/NutShellSim.scala 44:24]
  wire  memdelay_io_out_r_valid; // @[src/main/scala/sim/NutShellSim.scala 44:24]
  wire [63:0] memdelay_io_out_r_bits_data; // @[src/main/scala/sim/NutShellSim.scala 44:24]
  wire  memdelay_io_out_r_bits_last; // @[src/main/scala/sim/NutShellSim.scala 44:24]
  wire  mmio_clock; // @[src/main/scala/sim/NutShellSim.scala 45:20]
  wire  mmio_reset; // @[src/main/scala/sim/NutShellSim.scala 45:20]
  wire  mmio_io_rw_req_ready; // @[src/main/scala/sim/NutShellSim.scala 45:20]
  wire  mmio_io_rw_req_valid; // @[src/main/scala/sim/NutShellSim.scala 45:20]
  wire [31:0] mmio_io_rw_req_bits_addr; // @[src/main/scala/sim/NutShellSim.scala 45:20]
  wire [2:0] mmio_io_rw_req_bits_size; // @[src/main/scala/sim/NutShellSim.scala 45:20]
  wire [3:0] mmio_io_rw_req_bits_cmd; // @[src/main/scala/sim/NutShellSim.scala 45:20]
  wire [7:0] mmio_io_rw_req_bits_wmask; // @[src/main/scala/sim/NutShellSim.scala 45:20]
  wire [63:0] mmio_io_rw_req_bits_wdata; // @[src/main/scala/sim/NutShellSim.scala 45:20]
  wire  mmio_io_rw_resp_ready; // @[src/main/scala/sim/NutShellSim.scala 45:20]
  wire  mmio_io_rw_resp_valid; // @[src/main/scala/sim/NutShellSim.scala 45:20]
  wire [3:0] mmio_io_rw_resp_bits_cmd; // @[src/main/scala/sim/NutShellSim.scala 45:20]
  wire [63:0] mmio_io_rw_resp_bits_rdata; // @[src/main/scala/sim/NutShellSim.scala 45:20]
  wire  mmio_io_meip; // @[src/main/scala/sim/NutShellSim.scala 45:20]
  wire  mmio_io_dma_aw_ready; // @[src/main/scala/sim/NutShellSim.scala 45:20]
  wire  mmio_io_dma_aw_valid; // @[src/main/scala/sim/NutShellSim.scala 45:20]
  wire [31:0] mmio_io_dma_aw_bits_addr; // @[src/main/scala/sim/NutShellSim.scala 45:20]
  wire [7:0] mmio_io_dma_aw_bits_len; // @[src/main/scala/sim/NutShellSim.scala 45:20]
  wire [2:0] mmio_io_dma_aw_bits_size; // @[src/main/scala/sim/NutShellSim.scala 45:20]
  wire  mmio_io_dma_w_ready; // @[src/main/scala/sim/NutShellSim.scala 45:20]
  wire  mmio_io_dma_w_valid; // @[src/main/scala/sim/NutShellSim.scala 45:20]
  wire [63:0] mmio_io_dma_w_bits_data; // @[src/main/scala/sim/NutShellSim.scala 45:20]
  wire [7:0] mmio_io_dma_w_bits_strb; // @[src/main/scala/sim/NutShellSim.scala 45:20]
  wire  mmio_io_dma_b_ready; // @[src/main/scala/sim/NutShellSim.scala 45:20]
  wire  mmio_io_dma_b_valid; // @[src/main/scala/sim/NutShellSim.scala 45:20]
  wire  mmio_io_dma_ar_ready; // @[src/main/scala/sim/NutShellSim.scala 45:20]
  wire  mmio_io_dma_ar_valid; // @[src/main/scala/sim/NutShellSim.scala 45:20]
  wire [31:0] mmio_io_dma_ar_bits_addr; // @[src/main/scala/sim/NutShellSim.scala 45:20]
  wire  mmio_io_dma_r_ready; // @[src/main/scala/sim/NutShellSim.scala 45:20]
  wire  mmio_io_dma_r_valid; // @[src/main/scala/sim/NutShellSim.scala 45:20]
  wire [63:0] mmio_io_dma_r_bits_data; // @[src/main/scala/sim/NutShellSim.scala 45:20]
  wire  mmio_io_uart_out_valid; // @[src/main/scala/sim/NutShellSim.scala 45:20]
  wire [7:0] mmio_io_uart_out_ch; // @[src/main/scala/sim/NutShellSim.scala 45:20]
  wire  mmio_io_uart_in_valid; // @[src/main/scala/sim/NutShellSim.scala 45:20]
  wire [7:0] mmio_io_uart_in_ch; // @[src/main/scala/sim/NutShellSim.scala 45:20]
  wire  mmio__WIRE_4; // @[src/main/scala/sim/NutShellSim.scala 45:20]
  reg [63:0] c; // @[src/main/scala/utils/GTimer.scala 24:20]
  wire [63:0] _c_T_1 = c + 64'h1; // @[src/main/scala/utils/GTimer.scala 25:12]
  reg [63:0] c_1; // @[src/main/scala/utils/GTimer.scala 24:20]
  wire [63:0] _c_T_3 = c_1 + 64'h1; // @[src/main/scala/utils/GTimer.scala 25:12]
  wire  DISPLAY_ENABLE = c >= io_logCtrl_log_begin & c_1 < io_logCtrl_log_end; // @[src/main/scala/sim/NutShellSim.scala 62:58]
  wire  _WIRE = DISPLAY_ENABLE; // @[src/main/scala/sim/NutShellSim.scala 62:58]
  NutShell soc ( // @[src/main/scala/sim/NutShellSim.scala 40:19]
    .clock(soc_clock),
    .reset(soc_reset),
    .io_mem_aw_ready(soc_io_mem_aw_ready),
    .io_mem_aw_valid(soc_io_mem_aw_valid),
    .io_mem_aw_bits_addr(soc_io_mem_aw_bits_addr),
    .io_mem_aw_bits_len(soc_io_mem_aw_bits_len),
    .io_mem_aw_bits_size(soc_io_mem_aw_bits_size),
    .io_mem_aw_bits_burst(soc_io_mem_aw_bits_burst),
    .io_mem_w_ready(soc_io_mem_w_ready),
    .io_mem_w_valid(soc_io_mem_w_valid),
    .io_mem_w_bits_data(soc_io_mem_w_bits_data),
    .io_mem_w_bits_last(soc_io_mem_w_bits_last),
    .io_mem_b_valid(soc_io_mem_b_valid),
    .io_mem_ar_ready(soc_io_mem_ar_ready),
    .io_mem_ar_valid(soc_io_mem_ar_valid),
    .io_mem_ar_bits_addr(soc_io_mem_ar_bits_addr),
    .io_mem_ar_bits_len(soc_io_mem_ar_bits_len),
    .io_mem_r_valid(soc_io_mem_r_valid),
    .io_mem_r_bits_data(soc_io_mem_r_bits_data),
    .io_mem_r_bits_last(soc_io_mem_r_bits_last),
    .io_mmio_req_ready(soc_io_mmio_req_ready),
    .io_mmio_req_valid(soc_io_mmio_req_valid),
    .io_mmio_req_bits_addr(soc_io_mmio_req_bits_addr),
    .io_mmio_req_bits_size(soc_io_mmio_req_bits_size),
    .io_mmio_req_bits_cmd(soc_io_mmio_req_bits_cmd),
    .io_mmio_req_bits_wmask(soc_io_mmio_req_bits_wmask),
    .io_mmio_req_bits_wdata(soc_io_mmio_req_bits_wdata),
    .io_mmio_resp_ready(soc_io_mmio_resp_ready),
    .io_mmio_resp_valid(soc_io_mmio_resp_valid),
    .io_mmio_resp_bits_cmd(soc_io_mmio_resp_bits_cmd),
    .io_mmio_resp_bits_rdata(soc_io_mmio_resp_bits_rdata),
    .io_frontend_aw_ready(soc_io_frontend_aw_ready),
    .io_frontend_aw_valid(soc_io_frontend_aw_valid),
    .io_frontend_aw_bits_addr(soc_io_frontend_aw_bits_addr),
    .io_frontend_aw_bits_len(soc_io_frontend_aw_bits_len),
    .io_frontend_aw_bits_size(soc_io_frontend_aw_bits_size),
    .io_frontend_w_ready(soc_io_frontend_w_ready),
    .io_frontend_w_valid(soc_io_frontend_w_valid),
    .io_frontend_w_bits_data(soc_io_frontend_w_bits_data),
    .io_frontend_w_bits_strb(soc_io_frontend_w_bits_strb),
    .io_frontend_b_ready(soc_io_frontend_b_ready),
    .io_frontend_b_valid(soc_io_frontend_b_valid),
    .io_frontend_ar_ready(soc_io_frontend_ar_ready),
    .io_frontend_ar_valid(soc_io_frontend_ar_valid),
    .io_frontend_ar_bits_addr(soc_io_frontend_ar_bits_addr),
    .io_frontend_r_ready(soc_io_frontend_r_ready),
    .io_frontend_r_valid(soc_io_frontend_r_valid),
    .io_frontend_r_bits_data(soc_io_frontend_r_bits_data),
    .io_meip(soc_io_meip),
    ._WIRE_4(soc__WIRE_4)
  );
  AXI4RAM mem ( // @[src/main/scala/sim/NutShellSim.scala 41:19]
    .clock(mem_clock),
    .reset(mem_reset),
    .io_in_aw_ready(mem_io_in_aw_ready),
    .io_in_aw_valid(mem_io_in_aw_valid),
    .io_in_aw_bits_addr(mem_io_in_aw_bits_addr),
    .io_in_w_ready(mem_io_in_w_ready),
    .io_in_w_valid(mem_io_in_w_valid),
    .io_in_w_bits_data(mem_io_in_w_bits_data),
    .io_in_w_bits_last(mem_io_in_w_bits_last),
    .io_in_b_valid(mem_io_in_b_valid),
    .io_in_ar_ready(mem_io_in_ar_ready),
    .io_in_ar_valid(mem_io_in_ar_valid),
    .io_in_ar_bits_addr(mem_io_in_ar_bits_addr),
    .io_in_ar_bits_len(mem_io_in_ar_bits_len),
    .io_in_ar_bits_size(mem_io_in_ar_bits_size),
    .io_in_ar_bits_burst(mem_io_in_ar_bits_burst),
    .io_in_r_valid(mem_io_in_r_valid),
    .io_in_r_bits_data(mem_io_in_r_bits_data),
    .io_in_r_bits_last(mem_io_in_r_bits_last)
  );
  AXI4Delayer memdelay ( // @[src/main/scala/sim/NutShellSim.scala 44:24]
    .io_in_aw_ready(memdelay_io_in_aw_ready),
    .io_in_aw_valid(memdelay_io_in_aw_valid),
    .io_in_aw_bits_addr(memdelay_io_in_aw_bits_addr),
    .io_in_aw_bits_len(memdelay_io_in_aw_bits_len),
    .io_in_aw_bits_size(memdelay_io_in_aw_bits_size),
    .io_in_aw_bits_burst(memdelay_io_in_aw_bits_burst),
    .io_in_w_ready(memdelay_io_in_w_ready),
    .io_in_w_valid(memdelay_io_in_w_valid),
    .io_in_w_bits_data(memdelay_io_in_w_bits_data),
    .io_in_w_bits_last(memdelay_io_in_w_bits_last),
    .io_in_b_valid(memdelay_io_in_b_valid),
    .io_in_ar_ready(memdelay_io_in_ar_ready),
    .io_in_ar_valid(memdelay_io_in_ar_valid),
    .io_in_ar_bits_addr(memdelay_io_in_ar_bits_addr),
    .io_in_ar_bits_len(memdelay_io_in_ar_bits_len),
    .io_in_r_valid(memdelay_io_in_r_valid),
    .io_in_r_bits_data(memdelay_io_in_r_bits_data),
    .io_in_r_bits_last(memdelay_io_in_r_bits_last),
    .io_out_aw_ready(memdelay_io_out_aw_ready),
    .io_out_aw_valid(memdelay_io_out_aw_valid),
    .io_out_aw_bits_addr(memdelay_io_out_aw_bits_addr),
    .io_out_w_ready(memdelay_io_out_w_ready),
    .io_out_w_valid(memdelay_io_out_w_valid),
    .io_out_w_bits_data(memdelay_io_out_w_bits_data),
    .io_out_w_bits_last(memdelay_io_out_w_bits_last),
    .io_out_b_valid(memdelay_io_out_b_valid),
    .io_out_ar_valid(memdelay_io_out_ar_valid),
    .io_out_ar_bits_addr(memdelay_io_out_ar_bits_addr),
    .io_out_ar_bits_len(memdelay_io_out_ar_bits_len),
    .io_out_ar_bits_size(memdelay_io_out_ar_bits_size),
    .io_out_ar_bits_burst(memdelay_io_out_ar_bits_burst),
    .io_out_r_valid(memdelay_io_out_r_valid),
    .io_out_r_bits_data(memdelay_io_out_r_bits_data),
    .io_out_r_bits_last(memdelay_io_out_r_bits_last)
  );
  SimMMIO mmio ( // @[src/main/scala/sim/NutShellSim.scala 45:20]
    .clock(mmio_clock),
    .reset(mmio_reset),
    .io_rw_req_ready(mmio_io_rw_req_ready),
    .io_rw_req_valid(mmio_io_rw_req_valid),
    .io_rw_req_bits_addr(mmio_io_rw_req_bits_addr),
    .io_rw_req_bits_size(mmio_io_rw_req_bits_size),
    .io_rw_req_bits_cmd(mmio_io_rw_req_bits_cmd),
    .io_rw_req_bits_wmask(mmio_io_rw_req_bits_wmask),
    .io_rw_req_bits_wdata(mmio_io_rw_req_bits_wdata),
    .io_rw_resp_ready(mmio_io_rw_resp_ready),
    .io_rw_resp_valid(mmio_io_rw_resp_valid),
    .io_rw_resp_bits_cmd(mmio_io_rw_resp_bits_cmd),
    .io_rw_resp_bits_rdata(mmio_io_rw_resp_bits_rdata),
    .io_meip(mmio_io_meip),
    .io_dma_aw_ready(mmio_io_dma_aw_ready),
    .io_dma_aw_valid(mmio_io_dma_aw_valid),
    .io_dma_aw_bits_addr(mmio_io_dma_aw_bits_addr),
    .io_dma_aw_bits_len(mmio_io_dma_aw_bits_len),
    .io_dma_aw_bits_size(mmio_io_dma_aw_bits_size),
    .io_dma_w_ready(mmio_io_dma_w_ready),
    .io_dma_w_valid(mmio_io_dma_w_valid),
    .io_dma_w_bits_data(mmio_io_dma_w_bits_data),
    .io_dma_w_bits_strb(mmio_io_dma_w_bits_strb),
    .io_dma_b_ready(mmio_io_dma_b_ready),
    .io_dma_b_valid(mmio_io_dma_b_valid),
    .io_dma_ar_ready(mmio_io_dma_ar_ready),
    .io_dma_ar_valid(mmio_io_dma_ar_valid),
    .io_dma_ar_bits_addr(mmio_io_dma_ar_bits_addr),
    .io_dma_r_ready(mmio_io_dma_r_ready),
    .io_dma_r_valid(mmio_io_dma_r_valid),
    .io_dma_r_bits_data(mmio_io_dma_r_bits_data),
    .io_uart_out_valid(mmio_io_uart_out_valid),
    .io_uart_out_ch(mmio_io_uart_out_ch),
    .io_uart_in_valid(mmio_io_uart_in_valid),
    .io_uart_in_ch(mmio_io_uart_in_ch),
    ._WIRE_4(mmio__WIRE_4)
  );
  assign io_uart_out_valid = mmio_io_uart_out_valid; // @[src/main/scala/sim/NutShellSim.scala 68:11]
  assign io_uart_out_ch = mmio_io_uart_out_ch; // @[src/main/scala/sim/NutShellSim.scala 68:11]
  assign io_uart_in_valid = mmio_io_uart_in_valid; // @[src/main/scala/sim/NutShellSim.scala 68:11]
  assign difftest_step = 1'h1; // @[difftest/src/main/scala/Difftest.scala 311:19]
  assign soc_clock = clock;
  assign soc_reset = reset;
  assign soc_io_mem_aw_ready = memdelay_io_in_aw_ready; // @[src/main/scala/sim/NutShellSim.scala 49:18]
  assign soc_io_mem_w_ready = memdelay_io_in_w_ready; // @[src/main/scala/sim/NutShellSim.scala 49:18]
  assign soc_io_mem_b_valid = memdelay_io_in_b_valid; // @[src/main/scala/sim/NutShellSim.scala 49:18]
  assign soc_io_mem_ar_ready = memdelay_io_in_ar_ready; // @[src/main/scala/sim/NutShellSim.scala 49:18]
  assign soc_io_mem_r_valid = memdelay_io_in_r_valid; // @[src/main/scala/sim/NutShellSim.scala 49:18]
  assign soc_io_mem_r_bits_data = memdelay_io_in_r_bits_data; // @[src/main/scala/sim/NutShellSim.scala 49:18]
  assign soc_io_mem_r_bits_last = memdelay_io_in_r_bits_last; // @[src/main/scala/sim/NutShellSim.scala 49:18]
  assign soc_io_mmio_req_ready = mmio_io_rw_req_ready; // @[src/main/scala/sim/NutShellSim.scala 52:14]
  assign soc_io_mmio_resp_valid = mmio_io_rw_resp_valid; // @[src/main/scala/sim/NutShellSim.scala 52:14]
  assign soc_io_mmio_resp_bits_cmd = mmio_io_rw_resp_bits_cmd; // @[src/main/scala/sim/NutShellSim.scala 52:14]
  assign soc_io_mmio_resp_bits_rdata = mmio_io_rw_resp_bits_rdata; // @[src/main/scala/sim/NutShellSim.scala 52:14]
  assign soc_io_frontend_aw_valid = mmio_io_dma_aw_valid; // @[src/main/scala/sim/NutShellSim.scala 47:19]
  assign soc_io_frontend_aw_bits_addr = mmio_io_dma_aw_bits_addr; // @[src/main/scala/sim/NutShellSim.scala 47:19]
  assign soc_io_frontend_aw_bits_len = mmio_io_dma_aw_bits_len; // @[src/main/scala/sim/NutShellSim.scala 47:19]
  assign soc_io_frontend_aw_bits_size = mmio_io_dma_aw_bits_size; // @[src/main/scala/sim/NutShellSim.scala 47:19]
  assign soc_io_frontend_w_valid = mmio_io_dma_w_valid; // @[src/main/scala/sim/NutShellSim.scala 47:19]
  assign soc_io_frontend_w_bits_data = mmio_io_dma_w_bits_data; // @[src/main/scala/sim/NutShellSim.scala 47:19]
  assign soc_io_frontend_w_bits_strb = mmio_io_dma_w_bits_strb; // @[src/main/scala/sim/NutShellSim.scala 47:19]
  assign soc_io_frontend_b_ready = mmio_io_dma_b_ready; // @[src/main/scala/sim/NutShellSim.scala 47:19]
  assign soc_io_frontend_ar_valid = mmio_io_dma_ar_valid; // @[src/main/scala/sim/NutShellSim.scala 47:19]
  assign soc_io_frontend_ar_bits_addr = mmio_io_dma_ar_bits_addr; // @[src/main/scala/sim/NutShellSim.scala 47:19]
  assign soc_io_frontend_r_ready = mmio_io_dma_r_ready; // @[src/main/scala/sim/NutShellSim.scala 47:19]
  assign soc_io_meip = mmio_io_meip; // @[src/main/scala/sim/NutShellSim.scala 54:15]
  assign soc__WIRE_4 = c >= io_logCtrl_log_begin & c_1 < io_logCtrl_log_end; // @[src/main/scala/sim/NutShellSim.scala 62:58]
  assign mem_clock = clock;
  assign mem_reset = reset;
  assign mem_io_in_aw_valid = memdelay_io_out_aw_valid; // @[src/main/scala/sim/NutShellSim.scala 50:13]
  assign mem_io_in_aw_bits_addr = memdelay_io_out_aw_bits_addr; // @[src/main/scala/sim/NutShellSim.scala 50:13]
  assign mem_io_in_w_valid = memdelay_io_out_w_valid; // @[src/main/scala/sim/NutShellSim.scala 50:13]
  assign mem_io_in_w_bits_data = memdelay_io_out_w_bits_data; // @[src/main/scala/sim/NutShellSim.scala 50:13]
  assign mem_io_in_w_bits_last = memdelay_io_out_w_bits_last; // @[src/main/scala/sim/NutShellSim.scala 50:13]
  assign mem_io_in_ar_valid = memdelay_io_out_ar_valid; // @[src/main/scala/sim/NutShellSim.scala 50:13]
  assign mem_io_in_ar_bits_addr = memdelay_io_out_ar_bits_addr; // @[src/main/scala/sim/NutShellSim.scala 50:13]
  assign mem_io_in_ar_bits_len = memdelay_io_out_ar_bits_len; // @[src/main/scala/sim/NutShellSim.scala 50:13]
  assign mem_io_in_ar_bits_size = memdelay_io_out_ar_bits_size; // @[src/main/scala/sim/NutShellSim.scala 50:13]
  assign mem_io_in_ar_bits_burst = memdelay_io_out_ar_bits_burst; // @[src/main/scala/sim/NutShellSim.scala 50:13]
  assign memdelay_io_in_aw_valid = soc_io_mem_aw_valid; // @[src/main/scala/sim/NutShellSim.scala 49:18]
  assign memdelay_io_in_aw_bits_addr = soc_io_mem_aw_bits_addr; // @[src/main/scala/sim/NutShellSim.scala 49:18]
  assign memdelay_io_in_aw_bits_len = soc_io_mem_aw_bits_len; // @[src/main/scala/sim/NutShellSim.scala 49:18]
  assign memdelay_io_in_aw_bits_size = soc_io_mem_aw_bits_size; // @[src/main/scala/sim/NutShellSim.scala 49:18]
  assign memdelay_io_in_aw_bits_burst = soc_io_mem_aw_bits_burst; // @[src/main/scala/sim/NutShellSim.scala 49:18]
  assign memdelay_io_in_w_valid = soc_io_mem_w_valid; // @[src/main/scala/sim/NutShellSim.scala 49:18]
  assign memdelay_io_in_w_bits_data = soc_io_mem_w_bits_data; // @[src/main/scala/sim/NutShellSim.scala 49:18]
  assign memdelay_io_in_w_bits_last = soc_io_mem_w_bits_last; // @[src/main/scala/sim/NutShellSim.scala 49:18]
  assign memdelay_io_in_ar_valid = soc_io_mem_ar_valid; // @[src/main/scala/sim/NutShellSim.scala 49:18]
  assign memdelay_io_in_ar_bits_addr = soc_io_mem_ar_bits_addr; // @[src/main/scala/sim/NutShellSim.scala 49:18]
  assign memdelay_io_in_ar_bits_len = soc_io_mem_ar_bits_len; // @[src/main/scala/sim/NutShellSim.scala 49:18]
  assign memdelay_io_out_aw_ready = mem_io_in_aw_ready; // @[src/main/scala/sim/NutShellSim.scala 50:13]
  assign memdelay_io_out_w_ready = mem_io_in_w_ready; // @[src/main/scala/sim/NutShellSim.scala 50:13]
  assign memdelay_io_out_b_valid = mem_io_in_b_valid; // @[src/main/scala/sim/NutShellSim.scala 50:13]
  assign memdelay_io_out_r_valid = mem_io_in_r_valid; // @[src/main/scala/sim/NutShellSim.scala 50:13]
  assign memdelay_io_out_r_bits_data = mem_io_in_r_bits_data; // @[src/main/scala/sim/NutShellSim.scala 50:13]
  assign memdelay_io_out_r_bits_last = mem_io_in_r_bits_last; // @[src/main/scala/sim/NutShellSim.scala 50:13]
  assign mmio_clock = clock;
  assign mmio_reset = reset;
  assign mmio_io_rw_req_valid = soc_io_mmio_req_valid; // @[src/main/scala/sim/NutShellSim.scala 52:14]
  assign mmio_io_rw_req_bits_addr = soc_io_mmio_req_bits_addr; // @[src/main/scala/sim/NutShellSim.scala 52:14]
  assign mmio_io_rw_req_bits_size = soc_io_mmio_req_bits_size; // @[src/main/scala/sim/NutShellSim.scala 52:14]
  assign mmio_io_rw_req_bits_cmd = soc_io_mmio_req_bits_cmd; // @[src/main/scala/sim/NutShellSim.scala 52:14]
  assign mmio_io_rw_req_bits_wmask = soc_io_mmio_req_bits_wmask; // @[src/main/scala/sim/NutShellSim.scala 52:14]
  assign mmio_io_rw_req_bits_wdata = soc_io_mmio_req_bits_wdata; // @[src/main/scala/sim/NutShellSim.scala 52:14]
  assign mmio_io_rw_resp_ready = soc_io_mmio_resp_ready; // @[src/main/scala/sim/NutShellSim.scala 52:14]
  assign mmio_io_dma_aw_ready = soc_io_frontend_aw_ready; // @[src/main/scala/sim/NutShellSim.scala 47:19]
  assign mmio_io_dma_w_ready = soc_io_frontend_w_ready; // @[src/main/scala/sim/NutShellSim.scala 47:19]
  assign mmio_io_dma_b_valid = soc_io_frontend_b_valid; // @[src/main/scala/sim/NutShellSim.scala 47:19]
  assign mmio_io_dma_ar_ready = soc_io_frontend_ar_ready; // @[src/main/scala/sim/NutShellSim.scala 47:19]
  assign mmio_io_dma_r_valid = soc_io_frontend_r_valid; // @[src/main/scala/sim/NutShellSim.scala 47:19]
  assign mmio_io_dma_r_bits_data = soc_io_frontend_r_bits_data; // @[src/main/scala/sim/NutShellSim.scala 47:19]
  assign mmio_io_uart_in_ch = io_uart_in_ch; // @[src/main/scala/sim/NutShellSim.scala 68:11]
  assign mmio__WIRE_4 = c >= io_logCtrl_log_begin & c_1 < io_logCtrl_log_end; // @[src/main/scala/sim/NutShellSim.scala 62:58]
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/utils/GTimer.scala 24:20]
      c <= 64'h0; // @[src/main/scala/utils/GTimer.scala 24:20]
    end else begin
      c <= _c_T_1; // @[src/main/scala/utils/GTimer.scala 25:7]
    end
    if (reset) begin // @[src/main/scala/utils/GTimer.scala 24:20]
      c_1 <= 64'h0; // @[src/main/scala/utils/GTimer.scala 24:20]
    end else begin
      c_1 <= _c_T_3; // @[src/main/scala/utils/GTimer.scala 25:7]
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_logCtrl_log_begin <= io_logCtrl_log_end)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at NutShellSim.scala:61 assert(log_begin <= log_end)\n"); // @[src/main/scala/sim/NutShellSim.scala 61:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(io_logCtrl_log_begin <= io_logCtrl_log_end) & ~reset) begin
          $fatal; // @[src/main/scala/sim/NutShellSim.scala 61:9]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  c = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  c_1 = _RAND_1[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
