module TransExcep(
    input           clock,
    input           intr,
    input [63:0]    cause,
    input [63:0]    pc
);

endmodule