
module DifftestMemInitializer();
       
endmodule
