module InstFinish (
    input           clock,
    input           is_mmio,
    input           valid,
    input [63:0]    pc,
    input [31:0]    inst,
    input [11:0]    rcsr_id
);

endmodule