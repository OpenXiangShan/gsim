module Fetch(
  input         clock,
  input         reset,
  output [31:0] io_instRead_addr, // @[playground/src/noop/fetch.scala 60:16]
  input  [63:0] io_instRead_inst, // @[playground/src/noop/fetch.scala 60:16]
  output        io_instRead_arvalid, // @[playground/src/noop/fetch.scala 60:16]
  input         io_instRead_rvalid, // @[playground/src/noop/fetch.scala 60:16]
  output [63:0] io_va2pa_vaddr, // @[playground/src/noop/fetch.scala 60:16]
  output        io_va2pa_vvalid, // @[playground/src/noop/fetch.scala 60:16]
  input  [31:0] io_va2pa_paddr, // @[playground/src/noop/fetch.scala 60:16]
  input         io_va2pa_pvalid, // @[playground/src/noop/fetch.scala 60:16]
  input  [63:0] io_va2pa_tlb_excep_cause, // @[playground/src/noop/fetch.scala 60:16]
  input  [63:0] io_va2pa_tlb_excep_tval, // @[playground/src/noop/fetch.scala 60:16]
  input         io_va2pa_tlb_excep_en, // @[playground/src/noop/fetch.scala 60:16]
  input  [63:0] io_reg2if_seq_pc, // @[playground/src/noop/fetch.scala 60:16]
  input         io_reg2if_valid, // @[playground/src/noop/fetch.scala 60:16]
  input  [63:0] io_wb2if_seq_pc, // @[playground/src/noop/fetch.scala 60:16]
  input         io_wb2if_valid, // @[playground/src/noop/fetch.scala 60:16]
  input         io_recov, // @[playground/src/noop/fetch.scala 60:16]
  input         io_intr_in_en, // @[playground/src/noop/fetch.scala 60:16]
  input  [63:0] io_intr_in_cause, // @[playground/src/noop/fetch.scala 60:16]
  input  [63:0] io_branchFail_seq_pc, // @[playground/src/noop/fetch.scala 60:16]
  input         io_branchFail_valid, // @[playground/src/noop/fetch.scala 60:16]
  output [31:0] io_if2id_inst, // @[playground/src/noop/fetch.scala 60:16]
  output [63:0] io_if2id_pc, // @[playground/src/noop/fetch.scala 60:16]
  output [63:0] io_if2id_excep_cause, // @[playground/src/noop/fetch.scala 60:16]
  output [63:0] io_if2id_excep_tval, // @[playground/src/noop/fetch.scala 60:16]
  output        io_if2id_excep_en, // @[playground/src/noop/fetch.scala 60:16]
  output [63:0] io_if2id_excep_pc, // @[playground/src/noop/fetch.scala 60:16]
  input         io_if2id_drop, // @[playground/src/noop/fetch.scala 60:16]
  input         io_if2id_stall, // @[playground/src/noop/fetch.scala 60:16]
  output        io_if2id_recov, // @[playground/src/noop/fetch.scala 60:16]
  output        io_if2id_valid, // @[playground/src/noop/fetch.scala 60:16]
  input         io_if2id_ready // @[playground/src/noop/fetch.scala 60:16]
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [63:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [63:0] _RAND_21;
  reg [63:0] _RAND_22;
  reg [63:0] _RAND_23;
  reg [63:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [63:0] _RAND_26;
  reg [63:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [63:0] _RAND_29;
  reg [63:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [127:0] _RAND_32;
  reg [63:0] _RAND_33;
  reg [63:0] _RAND_34;
  reg [63:0] _RAND_35;
  reg [63:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
`endif // RANDOMIZE_REG_INIT
  reg [63:0] pc; // @[playground/src/noop/fetch.scala 61:21]
  reg  drop1_r; // @[playground/src/noop/fetch.scala 63:26]
  reg  drop2_r; // @[playground/src/noop/fetch.scala 64:26]
  reg  drop3_r; // @[playground/src/noop/fetch.scala 65:26]
  reg  stall1_r; // @[playground/src/noop/fetch.scala 66:27]
  reg  stall2_r; // @[playground/src/noop/fetch.scala 67:27]
  reg  stall3_r; // @[playground/src/noop/fetch.scala 68:27]
  reg  recov3_r; // @[playground/src/noop/fetch.scala 71:27]
  wire  drop3_in = drop3_r | io_if2id_drop; // @[playground/src/noop/fetch.scala 83:28]
  wire  drop2_in = drop2_r | drop3_in; // @[playground/src/noop/fetch.scala 84:28]
  wire  drop1_in = drop1_r | drop2_in; // @[playground/src/noop/fetch.scala 85:28]
  wire  _stall3_in_T = ~io_if2id_drop; // @[playground/src/noop/fetch.scala 86:34]
  wire  stall3_in = stall3_r & ~io_if2id_drop | io_if2id_stall; // @[playground/src/noop/fetch.scala 86:50]
  wire  _stall2_in_T = ~drop3_in; // @[playground/src/noop/fetch.scala 87:34]
  wire  stall2_in = stall2_r & ~drop3_in | stall3_in; // @[playground/src/noop/fetch.scala 87:45]
  wire  _stall1_in_T = ~drop2_in; // @[playground/src/noop/fetch.scala 88:34]
  wire  stall1_in = stall1_r & ~drop2_in | stall2_in; // @[playground/src/noop/fetch.scala 88:45]
  reg  state; // @[playground/src/noop/fetch.scala 91:24]
  wire  _T = ~state; // @[playground/src/noop/fetch.scala 92:18]
  wire  _GEN_0 = stall1_in | state; // @[playground/src/noop/fetch.scala 94:28 95:23 91:24]
  reg [63:0] pc1_r; // @[playground/src/noop/fetch.scala 105:24]
  reg [63:0] excep1_r_cause; // @[playground/src/noop/fetch.scala 107:30]
  reg  excep1_r_en; // @[playground/src/noop/fetch.scala 107:30]
  reg  valid1_r; // @[playground/src/noop/fetch.scala 108:30]
  wire  hs_in = _T & ~drop1_in; // @[playground/src/noop/fetch.scala 109:39]
  wire [63:0] _cur_pc_T_1 = pc + 64'h8; // @[playground/src/noop/fetch.scala 114:40]
  reg  valid2_r; // @[playground/src/noop/fetch.scala 156:30]
  reg [1:0] buf_bitmap; // @[playground/src/noop/fetch.scala 212:34]
  wire  _T_14 = buf_bitmap == 2'h3; // @[playground/src/noop/fetch.scala 228:25]
  reg  excep_buf_en; // @[playground/src/noop/fetch.scala 213:34]
  reg  excep2_r_en; // @[playground/src/noop/fetch.scala 157:30]
  reg  reset_ic; // @[playground/src/noop/fetch.scala 217:30]
  wire  _T_19 = valid2_r & io_instRead_rvalid & ~reset_ic; // @[playground/src/noop/fetch.scala 233:51]
  wire  _GEN_76 = excep2_r_en & valid2_r | _T_19; // @[playground/src/noop/fetch.scala 229:44 231:17]
  wire  _GEN_88 = buf_bitmap == 2'h3 | excep_buf_en ? 1'h0 : _GEN_76; // @[playground/src/noop/fetch.scala 228:49 222:9]
  wire  hs2 = _stall2_in_T & _GEN_88; // @[playground/src/noop/fetch.scala 227:20 222:9]
  reg  reset_tlb; // @[playground/src/noop/fetch.scala 161:30]
  wire  _tlb_inp_valid_T_1 = io_va2pa_pvalid | io_va2pa_tlb_excep_en; // @[playground/src/noop/fetch.scala 166:58]
  wire  tlb_inp_valid = ~reset_tlb & (io_va2pa_pvalid | io_va2pa_tlb_excep_en); // @[playground/src/noop/fetch.scala 166:38]
  wire  _GEN_16 = (tlb_inp_valid | excep1_r_en) & valid1_r; // @[playground/src/noop/fetch.scala 172:49 173:17 168:9]
  wire  _GEN_17 = valid2_r & ~hs2 ? 1'h0 : _GEN_16; // @[playground/src/noop/fetch.scala 170:31 171:17]
  wire  hs1 = _stall1_in_T & _GEN_17; // @[playground/src/noop/fetch.scala 169:20 168:9]
  wire [63:0] cur_pc = hs1 ? _cur_pc_T_1 : pc; // @[src/main/scala/chisel3/util/Mux.scala 47:70]
  wire [63:0] _next_pc_T = io_branchFail_valid ? io_branchFail_seq_pc : cur_pc; // @[src/main/scala/chisel3/util/Mux.scala 47:70]
  wire  _GEN_10 = hs_in & io_intr_in_en; // @[playground/src/noop/fetch.scala 126:16 72:13]
  wire  _GEN_12 = hs1 ? 1'h0 : valid1_r; // @[playground/src/noop/fetch.scala 141:24 142:22 108:30]
  wire  _GEN_13 = hs_in | _GEN_12; // @[playground/src/noop/fetch.scala 139:20 140:22]
  wire  _GEN_14 = _stall1_in_T & _GEN_13; // @[playground/src/noop/fetch.scala 138:20 145:18]
  reg [63:0] pc2_r; // @[playground/src/noop/fetch.scala 154:30]
  reg [31:0] paddr2_r; // @[playground/src/noop/fetch.scala 155:30]
  reg [63:0] excep2_r_cause; // @[playground/src/noop/fetch.scala 157:30]
  reg [63:0] excep2_r_tval; // @[playground/src/noop/fetch.scala 157:30]
  reg [63:0] excep2_r_pc; // @[playground/src/noop/fetch.scala 157:30]
  wire  _GEN_19 = hs2 ? 1'h0 : valid2_r; // @[playground/src/noop/fetch.scala 181:24 182:22 156:30]
  wire  _GEN_20 = hs1 | _GEN_19; // @[playground/src/noop/fetch.scala 177:18 178:29]
  wire [63:0] _GEN_23 = io_va2pa_tlb_excep_en ? pc1_r : 64'h0; // @[playground/src/noop/fetch.scala 188:42 189:28 195:25]
  wire  _GEN_24 = io_va2pa_tlb_excep_en | excep1_r_en; // @[playground/src/noop/fetch.scala 188:42 190:28 195:25]
  wire [63:0] _GEN_25 = io_va2pa_tlb_excep_en ? io_va2pa_tlb_excep_tval : 64'h0; // @[playground/src/noop/fetch.scala 188:42 191:28 195:25]
  wire [63:0] _GEN_26 = io_va2pa_tlb_excep_en ? io_va2pa_tlb_excep_cause : excep1_r_cause; // @[playground/src/noop/fetch.scala 188:42 192:28 195:25]
  wire  _GEN_35 = io_va2pa_pvalid ? 1'h0 : io_va2pa_tlb_excep_en; // @[playground/src/noop/fetch.scala 185:36 72:33]
  wire  _GEN_43 = ~hs1 ? 1'h0 : _GEN_35; // @[playground/src/noop/fetch.scala 184:19 72:33]
  wire  _GEN_46 = _stall2_in_T & _GEN_20; // @[playground/src/noop/fetch.scala 176:20 198:18]
  wire  _GEN_54 = _stall2_in_T & _GEN_43; // @[playground/src/noop/fetch.scala 176:20 72:33]
  wire  cur_excep_en = hs1 ? _GEN_24 : excep2_r_en; // @[playground/src/noop/fetch.scala 202:27]
  reg [63:0] pc3_r; // @[playground/src/noop/fetch.scala 205:34]
  reg  valid3_r; // @[playground/src/noop/fetch.scala 206:34]
  reg [63:0] excep3_r_cause; // @[playground/src/noop/fetch.scala 207:34]
  reg [63:0] excep3_r_tval; // @[playground/src/noop/fetch.scala 207:34]
  reg  excep3_r_en; // @[playground/src/noop/fetch.scala 207:34]
  reg [63:0] excep3_r_pc; // @[playground/src/noop/fetch.scala 207:34]
  reg [63:0] next_pc_r; // @[playground/src/noop/fetch.scala 208:34]
  reg  wait_jmp_pc; // @[playground/src/noop/fetch.scala 209:34]
  reg [127:0] inst_buf; // @[playground/src/noop/fetch.scala 210:34]
  reg [63:0] buf_start_pc; // @[playground/src/noop/fetch.scala 211:34]
  reg [63:0] excep_buf_cause; // @[playground/src/noop/fetch.scala 213:34]
  reg [63:0] excep_buf_tval; // @[playground/src/noop/fetch.scala 213:34]
  reg [63:0] excep_buf_pc; // @[playground/src/noop/fetch.scala 213:34]
  reg [31:0] inst_r; // @[playground/src/noop/fetch.scala 214:34]
  reg  update_excep_pc; // @[playground/src/noop/fetch.scala 218:34]
  wire [63:0] buf_offset = next_pc_r - buf_start_pc; // @[playground/src/noop/fetch.scala 223:33]
  wire  hs_out = io_if2id_ready & io_if2id_valid; // @[playground/src/noop/fetch.scala 224:33]
  wire [127:0] _next_inst_buf_T_1 = {io_instRead_inst,inst_buf[63:0]}; // @[playground/src/noop/fetch.scala 236:37]
  wire [127:0] _next_inst_buf_T_2 = {64'h0,io_instRead_inst}; // @[playground/src/noop/fetch.scala 239:37]
  wire [63:0] _buf_start_pc_T_1 = {pc2_r[63:3],3'h0}; // @[playground/src/noop/fetch.scala 241:36]
  wire [63:0] _GEN_58 = wait_jmp_pc ? pc2_r : next_pc_r; // @[playground/src/noop/fetch.scala 242:34 243:33 208:34]
  wire  _GEN_59 = wait_jmp_pc ? 1'h0 : wait_jmp_pc; // @[playground/src/noop/fetch.scala 242:34 244:33 209:34]
  wire [127:0] _GEN_60 = buf_bitmap[0] ? _next_inst_buf_T_1 : _next_inst_buf_T_2; // @[playground/src/noop/fetch.scala 235:32 236:31 239:31]
  wire [1:0] _GEN_61 = buf_bitmap[0] ? 2'h3 : 2'h1; // @[playground/src/noop/fetch.scala 235:32 237:33 240:33]
  wire [63:0] _GEN_62 = buf_bitmap[0] ? buf_start_pc : _buf_start_pc_T_1; // @[playground/src/noop/fetch.scala 235:32 211:34 241:30]
  wire [63:0] _GEN_63 = buf_bitmap[0] ? next_pc_r : _GEN_58; // @[playground/src/noop/fetch.scala 235:32 208:34]
  wire  _GEN_64 = buf_bitmap[0] ? wait_jmp_pc : _GEN_59; // @[playground/src/noop/fetch.scala 235:32 209:34]
  wire [127:0] _GEN_66 = valid2_r & io_instRead_rvalid & ~reset_ic ? _GEN_60 : inst_buf; // @[playground/src/noop/fetch.scala 225:19 233:64]
  wire [1:0] _GEN_67 = valid2_r & io_instRead_rvalid & ~reset_ic ? _GEN_61 : buf_bitmap; // @[playground/src/noop/fetch.scala 226:21 233:64]
  wire [63:0] _GEN_68 = valid2_r & io_instRead_rvalid & ~reset_ic ? _GEN_62 : buf_start_pc; // @[playground/src/noop/fetch.scala 211:34 233:64]
  wire [63:0] _GEN_69 = valid2_r & io_instRead_rvalid & ~reset_ic ? _GEN_63 : next_pc_r; // @[playground/src/noop/fetch.scala 208:34 233:64]
  wire  _GEN_70 = valid2_r & io_instRead_rvalid & ~reset_ic ? _GEN_64 : wait_jmp_pc; // @[playground/src/noop/fetch.scala 209:34 233:64]
  wire  _GEN_73 = excep2_r_en & valid2_r ? excep2_r_en : excep_buf_en; // @[playground/src/noop/fetch.scala 229:44 230:23 213:34]
  wire [127:0] _GEN_78 = excep2_r_en & valid2_r ? inst_buf : _GEN_66; // @[playground/src/noop/fetch.scala 225:19 229:44]
  wire [1:0] _GEN_79 = excep2_r_en & valid2_r ? buf_bitmap : _GEN_67; // @[playground/src/noop/fetch.scala 226:21 229:44]
  wire [63:0] _GEN_80 = excep2_r_en & valid2_r ? buf_start_pc : _GEN_68; // @[playground/src/noop/fetch.scala 211:34 229:44]
  wire [63:0] _GEN_81 = excep2_r_en & valid2_r ? next_pc_r : _GEN_69; // @[playground/src/noop/fetch.scala 208:34 229:44]
  wire  _GEN_82 = excep2_r_en & valid2_r ? wait_jmp_pc : _GEN_70; // @[playground/src/noop/fetch.scala 209:34 229:44]
  wire  _GEN_85 = buf_bitmap == 2'h3 | excep_buf_en ? excep_buf_en : _GEN_73; // @[playground/src/noop/fetch.scala 213:34 228:49]
  wire [127:0] _GEN_90 = buf_bitmap == 2'h3 | excep_buf_en ? inst_buf : _GEN_78; // @[playground/src/noop/fetch.scala 225:19 228:49]
  wire [1:0] _GEN_91 = buf_bitmap == 2'h3 | excep_buf_en ? buf_bitmap : _GEN_79; // @[playground/src/noop/fetch.scala 226:21 228:49]
  wire [63:0] _GEN_92 = buf_bitmap == 2'h3 | excep_buf_en ? buf_start_pc : _GEN_80; // @[playground/src/noop/fetch.scala 211:34 228:49]
  wire [63:0] _GEN_93 = buf_bitmap == 2'h3 | excep_buf_en ? next_pc_r : _GEN_81; // @[playground/src/noop/fetch.scala 208:34 228:49]
  wire  _GEN_94 = buf_bitmap == 2'h3 | excep_buf_en ? wait_jmp_pc : _GEN_82; // @[playground/src/noop/fetch.scala 209:34 228:49]
  wire  _GEN_97 = _stall2_in_T & _GEN_85; // @[playground/src/noop/fetch.scala 227:20 252:22]
  wire [127:0] next_inst_buf = _stall2_in_T ? _GEN_90 : inst_buf; // @[playground/src/noop/fetch.scala 225:19 227:20]
  wire [1:0] next_buf_bitmap = _stall2_in_T ? _GEN_91 : buf_bitmap; // @[playground/src/noop/fetch.scala 227:20 226:21]
  wire [63:0] _GEN_104 = _stall2_in_T ? _GEN_92 : buf_start_pc; // @[playground/src/noop/fetch.scala 227:20 211:34]
  wire [63:0] _GEN_105 = _stall2_in_T ? _GEN_93 : next_pc_r; // @[playground/src/noop/fetch.scala 227:20 208:34]
  wire  _GEN_106 = _stall2_in_T ? _GEN_94 : 1'h1; // @[playground/src/noop/fetch.scala 227:20 254:21]
  wire [1:0] _GEN_107 = _stall2_in_T ? next_buf_bitmap : 2'h0; // @[playground/src/noop/fetch.scala 227:20 248:20 251:20]
  wire [127:0] _GEN_108 = _stall2_in_T ? next_inst_buf : inst_buf; // @[playground/src/noop/fetch.scala 227:20 249:18 210:34]
  wire [5:0] _top_inst32_T_1 = {buf_offset[2:0],3'h0}; // @[playground/src/noop/fetch.scala 258:37]
  wire [127:0] top_inst32 = inst_buf >> _top_inst32_T_1; // @[playground/src/noop/fetch.scala 258:31]
  wire  _top_inst_T_1 = top_inst32[1:0] == 2'h3; // @[playground/src/noop/fetch.scala 262:41]
  wire [31:0] _top_inst_T_3 = {16'h0,top_inst32[15:0]}; // @[playground/src/noop/fetch.scala 262:65]
  wire [127:0] _top_inst_T_4 = top_inst32[1:0] == 2'h3 ? top_inst32 : {{96'd0}, _top_inst_T_3}; // @[playground/src/noop/fetch.scala 262:24]
  wire  _T_22 = buf_bitmap == 2'h1; // @[playground/src/noop/fetch.scala 263:27]
  wire  _T_23 = buf_offset == 64'h6; // @[playground/src/noop/fetch.scala 264:25]
  wire  _T_27 = buf_offset <= 64'h4; // @[playground/src/noop/fetch.scala 267:31]
  wire [127:0] _GEN_111 = buf_offset <= 64'h4 ? _top_inst_T_4 : 128'h0; // @[playground/src/noop/fetch.scala 267:38 269:22 259:37]
  wire  _GEN_112 = buf_offset == 64'h6 & top_inst32[1:0] != 2'h3 | _T_27; // @[playground/src/noop/fetch.scala 264:60 265:24]
  wire [127:0] _GEN_113 = buf_offset == 64'h6 & top_inst32[1:0] != 2'h3 ? {{96'd0}, _top_inst_T_3} : _GEN_111; // @[playground/src/noop/fetch.scala 264:60 266:22]
  wire  _GEN_114 = buf_bitmap == 2'h1 & _GEN_112; // @[playground/src/noop/fetch.scala 259:16 263:35]
  wire [127:0] _GEN_115 = buf_bitmap == 2'h1 ? _GEN_113 : 128'h0; // @[playground/src/noop/fetch.scala 263:35 259:37]
  wire  inst_valid = _T_14 | _GEN_114; // @[playground/src/noop/fetch.scala 260:29 261:20]
  wire [127:0] _GEN_117 = _T_14 ? _top_inst_T_4 : _GEN_115; // @[playground/src/noop/fetch.scala 260:29 262:18]
  wire  fetch_page_fault_excep = excep_buf_cause == 64'hc; // @[playground/src/noop/fetch.scala 272:50]
  wire  cross_page_excep = fetch_page_fault_excep & _T_22 & _T_23 & _top_inst_T_1; // @[playground/src/noop/fetch.scala 273:95]
  wire [63:0] _excep3_r_T_tval = inst_valid ? 64'h0 : excep_buf_tval; // @[playground/src/noop/fetch.scala 277:31]
  wire [63:0] _excep3_r_T_pc = inst_valid ? 64'h0 : excep_buf_pc; // @[playground/src/noop/fetch.scala 277:31]
  wire [31:0] top_inst = _GEN_117[31:0]; // @[playground/src/noop/fetch.scala 257:24]
  wire [63:0] _excep3_r_tval_T_1 = next_pc_r + 64'h2; // @[playground/src/noop/fetch.scala 282:59]
  wire [63:0] _excep3_r_tval_T_2 = fetch_page_fault_excep ? next_pc_r : excep_buf_tval; // @[src/main/scala/chisel3/util/Mux.scala 47:70]
  wire [63:0] _excep3_r_tval_T_3 = cross_page_excep ? _excep3_r_tval_T_1 : _excep3_r_tval_T_2; // @[src/main/scala/chisel3/util/Mux.scala 47:70]
  wire [2:0] _next_pc_w_T_2 = top_inst[1:0] == 2'h3 ? 3'h4 : 3'h2; // @[playground/src/noop/fetch.scala 288:44]
  wire [63:0] _GEN_11 = {{61'd0}, _next_pc_w_T_2}; // @[playground/src/noop/fetch.scala 288:39]
  wire [63:0] next_pc_w = next_pc_r + _GEN_11; // @[playground/src/noop/fetch.scala 288:39]
  wire [63:0] _T_34 = next_pc_w - buf_start_pc; // @[playground/src/noop/fetch.scala 290:29]
  wire [63:0] _buf_start_pc_T_3 = buf_start_pc + 64'h8; // @[playground/src/noop/fetch.scala 291:46]
  wire [127:0] _inst_buf_T_1 = {64'h0,next_inst_buf[127:64]}; // @[playground/src/noop/fetch.scala 292:32]
  wire [1:0] _buf_bitmap_T_1 = {1'h0,next_buf_bitmap[1]}; // @[playground/src/noop/fetch.scala 293:34]
  wire  _T_38 = ~inst_valid; // @[playground/src/noop/fetch.scala 295:18]
  wire  _GEN_125 = hs_out ? 1'h0 : valid3_r; // @[playground/src/noop/fetch.scala 301:27 302:22 206:34]
  wire  _GEN_126 = (inst_valid | excep_buf_en) & (~valid3_r | hs_out) | _GEN_125; // @[playground/src/noop/fetch.scala 275:68 276:25]
  wire  _GEN_139 = (inst_valid | excep_buf_en) & (~valid3_r | hs_out) & _T_38; // @[playground/src/noop/fetch.scala 275:68 72:53]
  wire  _GEN_141 = _stall3_in_T & _GEN_126; // @[playground/src/noop/fetch.scala 274:25 305:18]
  wire  _GEN_154 = _stall3_in_T & _GEN_139; // @[playground/src/noop/fetch.scala 274:25 72:53]
  assign io_instRead_addr = hs1 ? io_va2pa_paddr : paddr2_r; // @[playground/src/noop/fetch.scala 201:28]
  assign io_instRead_arvalid = (hs1 | valid2_r) & _stall3_in_T & ~cur_excep_en; // @[playground/src/noop/fetch.scala 203:64]
  assign io_va2pa_vaddr = hs1 ? _cur_pc_T_1 : pc; // @[src/main/scala/chisel3/util/Mux.scala 47:70]
  assign io_va2pa_vvalid = hs_in & ~io_intr_in_en; // @[playground/src/noop/fetch.scala 150:30]
  assign io_if2id_inst = inst_r; // @[playground/src/noop/fetch.scala 308:25]
  assign io_if2id_pc = pc3_r; // @[playground/src/noop/fetch.scala 309:25]
  assign io_if2id_excep_cause = excep3_r_cause; // @[playground/src/noop/fetch.scala 310:25]
  assign io_if2id_excep_tval = excep3_r_tval; // @[playground/src/noop/fetch.scala 310:25]
  assign io_if2id_excep_en = excep3_r_en; // @[playground/src/noop/fetch.scala 310:25]
  assign io_if2id_excep_pc = excep3_r_pc; // @[playground/src/noop/fetch.scala 310:25]
  assign io_if2id_recov = recov3_r; // @[playground/src/noop/fetch.scala 312:25]
  assign io_if2id_valid = valid3_r; // @[playground/src/noop/fetch.scala 311:25]
  always @(posedge clock) begin
    if (reset) begin // @[playground/src/noop/fetch.scala 61:21]
      pc <= 64'h80000000; // @[playground/src/noop/fetch.scala 61:21]
    end else if (io_reg2if_valid) begin // @[src/main/scala/chisel3/util/Mux.scala 47:70]
      pc <= io_reg2if_seq_pc;
    end else if (io_wb2if_valid) begin // @[src/main/scala/chisel3/util/Mux.scala 47:70]
      pc <= io_wb2if_seq_pc;
    end else if (io_intr_in_en) begin // @[src/main/scala/chisel3/util/Mux.scala 47:70]
      pc <= cur_pc;
    end else begin
      pc <= _next_pc_T;
    end
    if (reset) begin // @[playground/src/noop/fetch.scala 63:26]
      drop1_r <= 1'h0; // @[playground/src/noop/fetch.scala 63:26]
    end else begin
      drop1_r <= _GEN_10;
    end
    if (reset) begin // @[playground/src/noop/fetch.scala 64:26]
      drop2_r <= 1'h0; // @[playground/src/noop/fetch.scala 64:26]
    end else begin
      drop2_r <= _GEN_54;
    end
    if (reset) begin // @[playground/src/noop/fetch.scala 65:26]
      drop3_r <= 1'h0; // @[playground/src/noop/fetch.scala 65:26]
    end else begin
      drop3_r <= _GEN_154;
    end
    if (reset) begin // @[playground/src/noop/fetch.scala 66:27]
      stall1_r <= 1'h0; // @[playground/src/noop/fetch.scala 66:27]
    end else begin
      stall1_r <= _GEN_10;
    end
    if (reset) begin // @[playground/src/noop/fetch.scala 67:27]
      stall2_r <= 1'h0; // @[playground/src/noop/fetch.scala 67:27]
    end else begin
      stall2_r <= _GEN_54;
    end
    if (reset) begin // @[playground/src/noop/fetch.scala 68:27]
      stall3_r <= 1'h0; // @[playground/src/noop/fetch.scala 68:27]
    end else begin
      stall3_r <= _GEN_154;
    end
    if (reset) begin // @[playground/src/noop/fetch.scala 71:27]
      recov3_r <= 1'h0; // @[playground/src/noop/fetch.scala 71:27]
    end else if (_stall3_in_T) begin // @[playground/src/noop/fetch.scala 274:25]
      if ((inst_valid | excep_buf_en) & (~valid3_r | hs_out)) begin // @[playground/src/noop/fetch.scala 275:68]
        recov3_r <= _T_38;
      end
    end
    if (reset) begin // @[playground/src/noop/fetch.scala 91:24]
      state <= 1'h0; // @[playground/src/noop/fetch.scala 91:24]
    end else if (~state) begin // @[playground/src/noop/fetch.scala 92:18]
      state <= _GEN_0;
    end else if (state) begin // @[playground/src/noop/fetch.scala 92:18]
      if (drop1_in & ~stall1_in | io_recov) begin // @[playground/src/noop/fetch.scala 99:55]
        state <= 1'h0; // @[playground/src/noop/fetch.scala 100:23]
      end
    end
    if (reset) begin // @[playground/src/noop/fetch.scala 105:24]
      pc1_r <= 64'h0; // @[playground/src/noop/fetch.scala 105:24]
    end else if (hs1) begin // @[src/main/scala/chisel3/util/Mux.scala 47:70]
      pc1_r <= _cur_pc_T_1;
    end else begin
      pc1_r <= pc;
    end
    if (reset) begin // @[playground/src/noop/fetch.scala 107:30]
      excep1_r_cause <= 64'h0; // @[playground/src/noop/fetch.scala 107:30]
    end else if (hs_in) begin // @[playground/src/noop/fetch.scala 126:16]
      excep1_r_cause <= io_intr_in_cause; // @[playground/src/noop/fetch.scala 129:25]
    end
    if (reset) begin // @[playground/src/noop/fetch.scala 107:30]
      excep1_r_en <= 1'h0; // @[playground/src/noop/fetch.scala 107:30]
    end else if (hs_in) begin // @[playground/src/noop/fetch.scala 126:16]
      excep1_r_en <= io_intr_in_en; // @[playground/src/noop/fetch.scala 127:25]
    end
    if (reset) begin // @[playground/src/noop/fetch.scala 108:30]
      valid1_r <= 1'h0; // @[playground/src/noop/fetch.scala 108:30]
    end else begin
      valid1_r <= _GEN_14;
    end
    if (reset) begin // @[playground/src/noop/fetch.scala 156:30]
      valid2_r <= 1'h0; // @[playground/src/noop/fetch.scala 156:30]
    end else begin
      valid2_r <= _GEN_46;
    end
    if (reset) begin // @[playground/src/noop/fetch.scala 212:34]
      buf_bitmap <= 2'h0; // @[playground/src/noop/fetch.scala 212:34]
    end else if (_stall3_in_T) begin // @[playground/src/noop/fetch.scala 274:25]
      if ((inst_valid | excep_buf_en) & (~valid3_r | hs_out)) begin // @[playground/src/noop/fetch.scala 275:68]
        if (_T_34 >= 64'h8 & buf_bitmap != 2'h0) begin // @[playground/src/noop/fetch.scala 290:74]
          buf_bitmap <= _buf_bitmap_T_1; // @[playground/src/noop/fetch.scala 293:28]
        end else begin
          buf_bitmap <= _GEN_107;
        end
      end else begin
        buf_bitmap <= _GEN_107;
      end
    end else begin
      buf_bitmap <= _GEN_107;
    end
    if (reset) begin // @[playground/src/noop/fetch.scala 213:34]
      excep_buf_en <= 1'h0; // @[playground/src/noop/fetch.scala 213:34]
    end else if (_stall3_in_T) begin // @[playground/src/noop/fetch.scala 274:25]
      if ((inst_valid | excep_buf_en) & (~valid3_r | hs_out)) begin // @[playground/src/noop/fetch.scala 275:68]
        if (~inst_valid) begin // @[playground/src/noop/fetch.scala 295:30]
          excep_buf_en <= 1'h0; // @[playground/src/noop/fetch.scala 296:30]
        end else begin
          excep_buf_en <= _GEN_97;
        end
      end else begin
        excep_buf_en <= _GEN_97;
      end
    end else begin
      excep_buf_en <= _GEN_97;
    end
    if (reset) begin // @[playground/src/noop/fetch.scala 157:30]
      excep2_r_en <= 1'h0; // @[playground/src/noop/fetch.scala 157:30]
    end else if (_stall2_in_T) begin // @[playground/src/noop/fetch.scala 176:20]
      if (!(~hs1)) begin // @[playground/src/noop/fetch.scala 184:19]
        if (io_va2pa_pvalid) begin // @[playground/src/noop/fetch.scala 185:36]
          excep2_r_en <= 1'h0; // @[playground/src/noop/fetch.scala 187:28]
        end else begin
          excep2_r_en <= _GEN_24;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/fetch.scala 217:30]
      reset_ic <= 1'h0; // @[playground/src/noop/fetch.scala 217:30]
    end else if (_stall2_in_T) begin // @[playground/src/noop/fetch.scala 227:20]
      if (io_instRead_rvalid) begin // @[playground/src/noop/fetch.scala 219:29]
        reset_ic <= 1'h0; // @[playground/src/noop/fetch.scala 220:18]
      end
    end else begin
      reset_ic <= reset_ic | valid2_r & ~excep2_r_en & ~io_instRead_rvalid; // @[playground/src/noop/fetch.scala 253:18]
    end
    if (reset) begin // @[playground/src/noop/fetch.scala 161:30]
      reset_tlb <= 1'h0; // @[playground/src/noop/fetch.scala 161:30]
    end else if (_stall2_in_T) begin // @[playground/src/noop/fetch.scala 176:20]
      if (_tlb_inp_valid_T_1) begin // @[playground/src/noop/fetch.scala 162:51]
        reset_tlb <= 1'h0; // @[playground/src/noop/fetch.scala 163:21]
      end
    end else begin
      reset_tlb <= ~_tlb_inp_valid_T_1; // @[playground/src/noop/fetch.scala 199:19]
    end
    if (reset) begin // @[playground/src/noop/fetch.scala 154:30]
      pc2_r <= 64'h0; // @[playground/src/noop/fetch.scala 154:30]
    end else if (_stall2_in_T) begin // @[playground/src/noop/fetch.scala 176:20]
      if (hs1) begin // @[playground/src/noop/fetch.scala 177:18]
        pc2_r <= pc1_r; // @[playground/src/noop/fetch.scala 179:29]
      end
    end
    if (reset) begin // @[playground/src/noop/fetch.scala 155:30]
      paddr2_r <= 32'h0; // @[playground/src/noop/fetch.scala 155:30]
    end else if (_stall2_in_T) begin // @[playground/src/noop/fetch.scala 176:20]
      if (!(~hs1)) begin // @[playground/src/noop/fetch.scala 184:19]
        if (io_va2pa_pvalid) begin // @[playground/src/noop/fetch.scala 185:36]
          paddr2_r <= io_va2pa_paddr; // @[playground/src/noop/fetch.scala 186:25]
        end
      end
    end
    if (reset) begin // @[playground/src/noop/fetch.scala 157:30]
      excep2_r_cause <= 64'h0; // @[playground/src/noop/fetch.scala 157:30]
    end else if (_stall2_in_T) begin // @[playground/src/noop/fetch.scala 176:20]
      if (!(~hs1)) begin // @[playground/src/noop/fetch.scala 184:19]
        if (!(io_va2pa_pvalid)) begin // @[playground/src/noop/fetch.scala 185:36]
          excep2_r_cause <= _GEN_26;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/fetch.scala 157:30]
      excep2_r_tval <= 64'h0; // @[playground/src/noop/fetch.scala 157:30]
    end else if (_stall2_in_T) begin // @[playground/src/noop/fetch.scala 176:20]
      if (!(~hs1)) begin // @[playground/src/noop/fetch.scala 184:19]
        if (!(io_va2pa_pvalid)) begin // @[playground/src/noop/fetch.scala 185:36]
          excep2_r_tval <= _GEN_25;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/fetch.scala 157:30]
      excep2_r_pc <= 64'h0; // @[playground/src/noop/fetch.scala 157:30]
    end else if (_stall2_in_T) begin // @[playground/src/noop/fetch.scala 176:20]
      if (!(~hs1)) begin // @[playground/src/noop/fetch.scala 184:19]
        if (!(io_va2pa_pvalid)) begin // @[playground/src/noop/fetch.scala 185:36]
          excep2_r_pc <= _GEN_23;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/fetch.scala 205:34]
      pc3_r <= 64'h0; // @[playground/src/noop/fetch.scala 205:34]
    end else if (_stall3_in_T) begin // @[playground/src/noop/fetch.scala 274:25]
      if ((inst_valid | excep_buf_en) & (~valid3_r | hs_out)) begin // @[playground/src/noop/fetch.scala 275:68]
        pc3_r <= next_pc_r; // @[playground/src/noop/fetch.scala 287:25]
      end
    end
    if (reset) begin // @[playground/src/noop/fetch.scala 206:34]
      valid3_r <= 1'h0; // @[playground/src/noop/fetch.scala 206:34]
    end else begin
      valid3_r <= _GEN_141;
    end
    if (reset) begin // @[playground/src/noop/fetch.scala 207:34]
      excep3_r_cause <= 64'h0; // @[playground/src/noop/fetch.scala 207:34]
    end else if (_stall3_in_T) begin // @[playground/src/noop/fetch.scala 274:25]
      if ((inst_valid | excep_buf_en) & (~valid3_r | hs_out)) begin // @[playground/src/noop/fetch.scala 275:68]
        if (inst_valid) begin // @[playground/src/noop/fetch.scala 277:31]
          excep3_r_cause <= 64'h0;
        end else begin
          excep3_r_cause <= excep_buf_cause;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/fetch.scala 207:34]
      excep3_r_tval <= 64'h0; // @[playground/src/noop/fetch.scala 207:34]
    end else if (_stall3_in_T) begin // @[playground/src/noop/fetch.scala 274:25]
      if ((inst_valid | excep_buf_en) & (~valid3_r | hs_out)) begin // @[playground/src/noop/fetch.scala 275:68]
        if (update_excep_pc) begin // @[playground/src/noop/fetch.scala 279:34]
          excep3_r_tval <= _excep3_r_tval_T_3; // @[playground/src/noop/fetch.scala 281:31]
        end else begin
          excep3_r_tval <= _excep3_r_T_tval; // @[playground/src/noop/fetch.scala 277:25]
        end
      end
    end
    if (reset) begin // @[playground/src/noop/fetch.scala 207:34]
      excep3_r_en <= 1'h0; // @[playground/src/noop/fetch.scala 207:34]
    end else if (_stall3_in_T) begin // @[playground/src/noop/fetch.scala 274:25]
      if ((inst_valid | excep_buf_en) & (~valid3_r | hs_out)) begin // @[playground/src/noop/fetch.scala 275:68]
        if (inst_valid) begin // @[playground/src/noop/fetch.scala 277:31]
          excep3_r_en <= 1'h0;
        end else begin
          excep3_r_en <= excep_buf_en;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/fetch.scala 207:34]
      excep3_r_pc <= 64'h0; // @[playground/src/noop/fetch.scala 207:34]
    end else if (_stall3_in_T) begin // @[playground/src/noop/fetch.scala 274:25]
      if ((inst_valid | excep_buf_en) & (~valid3_r | hs_out)) begin // @[playground/src/noop/fetch.scala 275:68]
        if (update_excep_pc) begin // @[playground/src/noop/fetch.scala 279:34]
          excep3_r_pc <= next_pc_r; // @[playground/src/noop/fetch.scala 280:29]
        end else begin
          excep3_r_pc <= _excep3_r_T_pc; // @[playground/src/noop/fetch.scala 277:25]
        end
      end
    end
    if (reset) begin // @[playground/src/noop/fetch.scala 208:34]
      next_pc_r <= 64'h0; // @[playground/src/noop/fetch.scala 208:34]
    end else if (_stall3_in_T) begin // @[playground/src/noop/fetch.scala 274:25]
      if ((inst_valid | excep_buf_en) & (~valid3_r | hs_out)) begin // @[playground/src/noop/fetch.scala 275:68]
        next_pc_r <= next_pc_w; // @[playground/src/noop/fetch.scala 289:25]
      end else begin
        next_pc_r <= _GEN_105;
      end
    end else begin
      next_pc_r <= _GEN_105;
    end
    wait_jmp_pc <= reset | _GEN_106; // @[playground/src/noop/fetch.scala 209:{34,34}]
    if (reset) begin // @[playground/src/noop/fetch.scala 210:34]
      inst_buf <= 128'h0; // @[playground/src/noop/fetch.scala 210:34]
    end else if (_stall3_in_T) begin // @[playground/src/noop/fetch.scala 274:25]
      if ((inst_valid | excep_buf_en) & (~valid3_r | hs_out)) begin // @[playground/src/noop/fetch.scala 275:68]
        if (_T_34 >= 64'h8 & buf_bitmap != 2'h0) begin // @[playground/src/noop/fetch.scala 290:74]
          inst_buf <= _inst_buf_T_1; // @[playground/src/noop/fetch.scala 292:26]
        end else begin
          inst_buf <= _GEN_108;
        end
      end else begin
        inst_buf <= _GEN_108;
      end
    end else begin
      inst_buf <= _GEN_108;
    end
    if (reset) begin // @[playground/src/noop/fetch.scala 211:34]
      buf_start_pc <= 64'h0; // @[playground/src/noop/fetch.scala 211:34]
    end else if (_stall3_in_T) begin // @[playground/src/noop/fetch.scala 274:25]
      if ((inst_valid | excep_buf_en) & (~valid3_r | hs_out)) begin // @[playground/src/noop/fetch.scala 275:68]
        if (_T_34 >= 64'h8 & buf_bitmap != 2'h0) begin // @[playground/src/noop/fetch.scala 290:74]
          buf_start_pc <= _buf_start_pc_T_3; // @[playground/src/noop/fetch.scala 291:30]
        end else begin
          buf_start_pc <= _GEN_104;
        end
      end else begin
        buf_start_pc <= _GEN_104;
      end
    end else begin
      buf_start_pc <= _GEN_104;
    end
    if (reset) begin // @[playground/src/noop/fetch.scala 213:34]
      excep_buf_cause <= 64'h0; // @[playground/src/noop/fetch.scala 213:34]
    end else if (_stall2_in_T) begin // @[playground/src/noop/fetch.scala 227:20]
      if (!(buf_bitmap == 2'h3 | excep_buf_en)) begin // @[playground/src/noop/fetch.scala 228:49]
        if (excep2_r_en & valid2_r) begin // @[playground/src/noop/fetch.scala 229:44]
          excep_buf_cause <= excep2_r_cause; // @[playground/src/noop/fetch.scala 230:23]
        end
      end
    end
    if (reset) begin // @[playground/src/noop/fetch.scala 213:34]
      excep_buf_tval <= 64'h0; // @[playground/src/noop/fetch.scala 213:34]
    end else if (_stall2_in_T) begin // @[playground/src/noop/fetch.scala 227:20]
      if (!(buf_bitmap == 2'h3 | excep_buf_en)) begin // @[playground/src/noop/fetch.scala 228:49]
        if (excep2_r_en & valid2_r) begin // @[playground/src/noop/fetch.scala 229:44]
          excep_buf_tval <= excep2_r_tval; // @[playground/src/noop/fetch.scala 230:23]
        end
      end
    end
    if (reset) begin // @[playground/src/noop/fetch.scala 213:34]
      excep_buf_pc <= 64'h0; // @[playground/src/noop/fetch.scala 213:34]
    end else if (_stall2_in_T) begin // @[playground/src/noop/fetch.scala 227:20]
      if (!(buf_bitmap == 2'h3 | excep_buf_en)) begin // @[playground/src/noop/fetch.scala 228:49]
        if (excep2_r_en & valid2_r) begin // @[playground/src/noop/fetch.scala 229:44]
          excep_buf_pc <= excep2_r_pc; // @[playground/src/noop/fetch.scala 230:23]
        end
      end
    end
    if (reset) begin // @[playground/src/noop/fetch.scala 214:34]
      inst_r <= 32'h0; // @[playground/src/noop/fetch.scala 214:34]
    end else if (_stall3_in_T) begin // @[playground/src/noop/fetch.scala 274:25]
      if ((inst_valid | excep_buf_en) & (~valid3_r | hs_out)) begin // @[playground/src/noop/fetch.scala 275:68]
        if (inst_valid) begin // @[playground/src/noop/fetch.scala 278:31]
          inst_r <= top_inst;
        end else begin
          inst_r <= 32'h0;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/fetch.scala 218:34]
      update_excep_pc <= 1'h0; // @[playground/src/noop/fetch.scala 218:34]
    end else if (_stall2_in_T) begin // @[playground/src/noop/fetch.scala 227:20]
      if (!(buf_bitmap == 2'h3 | excep_buf_en)) begin // @[playground/src/noop/fetch.scala 228:49]
        if (excep2_r_en & valid2_r) begin // @[playground/src/noop/fetch.scala 229:44]
          update_excep_pc <= ~wait_jmp_pc; // @[playground/src/noop/fetch.scala 232:29]
        end
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  pc = _RAND_0[63:0];
  _RAND_1 = {1{`RANDOM}};
  drop1_r = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  drop2_r = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  drop3_r = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  stall1_r = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  stall2_r = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  stall3_r = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  recov3_r = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  state = _RAND_8[0:0];
  _RAND_9 = {2{`RANDOM}};
  pc1_r = _RAND_9[63:0];
  _RAND_10 = {2{`RANDOM}};
  excep1_r_cause = _RAND_10[63:0];
  _RAND_11 = {1{`RANDOM}};
  excep1_r_en = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  valid1_r = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  valid2_r = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  buf_bitmap = _RAND_14[1:0];
  _RAND_15 = {1{`RANDOM}};
  excep_buf_en = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  excep2_r_en = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  reset_ic = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  reset_tlb = _RAND_18[0:0];
  _RAND_19 = {2{`RANDOM}};
  pc2_r = _RAND_19[63:0];
  _RAND_20 = {1{`RANDOM}};
  paddr2_r = _RAND_20[31:0];
  _RAND_21 = {2{`RANDOM}};
  excep2_r_cause = _RAND_21[63:0];
  _RAND_22 = {2{`RANDOM}};
  excep2_r_tval = _RAND_22[63:0];
  _RAND_23 = {2{`RANDOM}};
  excep2_r_pc = _RAND_23[63:0];
  _RAND_24 = {2{`RANDOM}};
  pc3_r = _RAND_24[63:0];
  _RAND_25 = {1{`RANDOM}};
  valid3_r = _RAND_25[0:0];
  _RAND_26 = {2{`RANDOM}};
  excep3_r_cause = _RAND_26[63:0];
  _RAND_27 = {2{`RANDOM}};
  excep3_r_tval = _RAND_27[63:0];
  _RAND_28 = {1{`RANDOM}};
  excep3_r_en = _RAND_28[0:0];
  _RAND_29 = {2{`RANDOM}};
  excep3_r_pc = _RAND_29[63:0];
  _RAND_30 = {2{`RANDOM}};
  next_pc_r = _RAND_30[63:0];
  _RAND_31 = {1{`RANDOM}};
  wait_jmp_pc = _RAND_31[0:0];
  _RAND_32 = {4{`RANDOM}};
  inst_buf = _RAND_32[127:0];
  _RAND_33 = {2{`RANDOM}};
  buf_start_pc = _RAND_33[63:0];
  _RAND_34 = {2{`RANDOM}};
  excep_buf_cause = _RAND_34[63:0];
  _RAND_35 = {2{`RANDOM}};
  excep_buf_tval = _RAND_35[63:0];
  _RAND_36 = {2{`RANDOM}};
  excep_buf_pc = _RAND_36[63:0];
  _RAND_37 = {1{`RANDOM}};
  inst_r = _RAND_37[31:0];
  _RAND_38 = {1{`RANDOM}};
  update_excep_pc = _RAND_38[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Decode(
  input         clock,
  input         reset,
  input  [31:0] io_if2id_inst, // @[playground/src/noop/decode.scala 11:16]
  input  [63:0] io_if2id_pc, // @[playground/src/noop/decode.scala 11:16]
  input  [63:0] io_if2id_excep_cause, // @[playground/src/noop/decode.scala 11:16]
  input  [63:0] io_if2id_excep_tval, // @[playground/src/noop/decode.scala 11:16]
  input         io_if2id_excep_en, // @[playground/src/noop/decode.scala 11:16]
  input  [63:0] io_if2id_excep_pc, // @[playground/src/noop/decode.scala 11:16]
  output        io_if2id_drop, // @[playground/src/noop/decode.scala 11:16]
  output        io_if2id_stall, // @[playground/src/noop/decode.scala 11:16]
  input         io_if2id_recov, // @[playground/src/noop/decode.scala 11:16]
  input         io_if2id_valid, // @[playground/src/noop/decode.scala 11:16]
  output        io_if2id_ready, // @[playground/src/noop/decode.scala 11:16]
  output [31:0] io_id2df_inst, // @[playground/src/noop/decode.scala 11:16]
  output [63:0] io_id2df_pc, // @[playground/src/noop/decode.scala 11:16]
  output [63:0] io_id2df_excep_cause, // @[playground/src/noop/decode.scala 11:16]
  output [63:0] io_id2df_excep_tval, // @[playground/src/noop/decode.scala 11:16]
  output        io_id2df_excep_en, // @[playground/src/noop/decode.scala 11:16]
  output [63:0] io_id2df_excep_pc, // @[playground/src/noop/decode.scala 11:16]
  output [1:0]  io_id2df_excep_etype, // @[playground/src/noop/decode.scala 11:16]
  output [4:0]  io_id2df_ctrl_aluOp, // @[playground/src/noop/decode.scala 11:16]
  output        io_id2df_ctrl_aluWidth, // @[playground/src/noop/decode.scala 11:16]
  output [4:0]  io_id2df_ctrl_dcMode, // @[playground/src/noop/decode.scala 11:16]
  output        io_id2df_ctrl_writeRegEn, // @[playground/src/noop/decode.scala 11:16]
  output        io_id2df_ctrl_writeCSREn, // @[playground/src/noop/decode.scala 11:16]
  output [2:0]  io_id2df_ctrl_brType, // @[playground/src/noop/decode.scala 11:16]
  output [4:0]  io_id2df_rs1, // @[playground/src/noop/decode.scala 11:16]
  output        io_id2df_rrs1, // @[playground/src/noop/decode.scala 11:16]
  output [63:0] io_id2df_rs1_d, // @[playground/src/noop/decode.scala 11:16]
  output [11:0] io_id2df_rs2, // @[playground/src/noop/decode.scala 11:16]
  output        io_id2df_rrs2, // @[playground/src/noop/decode.scala 11:16]
  output [63:0] io_id2df_rs2_d, // @[playground/src/noop/decode.scala 11:16]
  output [4:0]  io_id2df_dst, // @[playground/src/noop/decode.scala 11:16]
  output [63:0] io_id2df_dst_d, // @[playground/src/noop/decode.scala 11:16]
  output [1:0]  io_id2df_jmp_type, // @[playground/src/noop/decode.scala 11:16]
  output [1:0]  io_id2df_special, // @[playground/src/noop/decode.scala 11:16]
  output [5:0]  io_id2df_swap, // @[playground/src/noop/decode.scala 11:16]
  output [1:0]  io_id2df_indi, // @[playground/src/noop/decode.scala 11:16]
  input         io_id2df_drop, // @[playground/src/noop/decode.scala 11:16]
  input         io_id2df_stall, // @[playground/src/noop/decode.scala 11:16]
  output        io_id2df_recov, // @[playground/src/noop/decode.scala 11:16]
  output        io_id2df_valid, // @[playground/src/noop/decode.scala 11:16]
  input         io_id2df_ready, // @[playground/src/noop/decode.scala 11:16]
  input  [1:0]  io_idState_priv // @[playground/src/noop/decode.scala 11:16]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [63:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [63:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [63:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
`endif // RANDOMIZE_REG_INIT
  reg  drop_r; // @[playground/src/noop/decode.scala 17:30]
  reg  stall_r; // @[playground/src/noop/decode.scala 18:30]
  wire  drop_in = drop_r | io_id2df_drop; // @[playground/src/noop/decode.scala 20:30]
  wire  _io_if2id_stall_T = ~io_id2df_drop; // @[playground/src/noop/decode.scala 22:36]
  reg [31:0] inst_r; // @[playground/src/noop/decode.scala 23:30]
  reg [63:0] pc_r; // @[playground/src/noop/decode.scala 24:30]
  reg [63:0] excep_r_cause; // @[playground/src/noop/decode.scala 25:30]
  reg [63:0] excep_r_tval; // @[playground/src/noop/decode.scala 25:30]
  reg  excep_r_en; // @[playground/src/noop/decode.scala 25:30]
  reg [63:0] excep_r_pc; // @[playground/src/noop/decode.scala 25:30]
  reg [1:0] excep_r_etype; // @[playground/src/noop/decode.scala 25:30]
  reg [4:0] ctrl_r_aluOp; // @[playground/src/noop/decode.scala 26:30]
  reg  ctrl_r_aluWidth; // @[playground/src/noop/decode.scala 26:30]
  reg [4:0] ctrl_r_dcMode; // @[playground/src/noop/decode.scala 26:30]
  reg  ctrl_r_writeRegEn; // @[playground/src/noop/decode.scala 26:30]
  reg  ctrl_r_writeCSREn; // @[playground/src/noop/decode.scala 26:30]
  reg [2:0] ctrl_r_brType; // @[playground/src/noop/decode.scala 26:30]
  reg [4:0] rs1_r; // @[playground/src/noop/decode.scala 27:30]
  reg  rrs1_r; // @[playground/src/noop/decode.scala 28:30]
  reg [63:0] rs1_d_r; // @[playground/src/noop/decode.scala 29:30]
  reg [11:0] rs2_r; // @[playground/src/noop/decode.scala 30:30]
  reg  rrs2_r; // @[playground/src/noop/decode.scala 31:30]
  reg [63:0] rs2_d_r; // @[playground/src/noop/decode.scala 32:30]
  reg [4:0] dst_r; // @[playground/src/noop/decode.scala 33:30]
  reg [63:0] dst_d_r; // @[playground/src/noop/decode.scala 34:30]
  reg [1:0] jmp_type_r; // @[playground/src/noop/decode.scala 35:30]
  reg [1:0] special_r; // @[playground/src/noop/decode.scala 36:30]
  reg [5:0] swap_r; // @[playground/src/noop/decode.scala 37:30]
  reg [1:0] indi_r; // @[playground/src/noop/decode.scala 38:30]
  reg  recov_r; // @[playground/src/noop/decode.scala 39:30]
  reg  valid_r; // @[playground/src/noop/decode.scala 40:30]
  wire  hs_out = io_id2df_ready & io_id2df_valid; // @[playground/src/noop/decode.scala 46:33]
  wire  hs_in = io_if2id_ready & io_if2id_valid; // @[playground/src/noop/decode.scala 47:33]
  wire [31:0] _instType_T = io_if2id_inst & 32'h7f; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _instType_T_1 = 32'h37 == _instType_T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _instType_T_3 = 32'h17 == _instType_T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _instType_T_5 = 32'h6f == _instType_T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire [31:0] _instType_T_6 = io_if2id_inst & 32'h707f; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _instType_T_7 = 32'h67 == _instType_T_6; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _instType_T_9 = 32'h63 == _instType_T_6; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _instType_T_11 = 32'h1063 == _instType_T_6; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _instType_T_13 = 32'h4063 == _instType_T_6; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _instType_T_15 = 32'h5063 == _instType_T_6; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _instType_T_17 = 32'h6063 == _instType_T_6; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _instType_T_19 = 32'h7063 == _instType_T_6; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _instType_T_21 = 32'h3 == _instType_T_6; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _instType_T_23 = 32'h1003 == _instType_T_6; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _instType_T_25 = 32'h2003 == _instType_T_6; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _instType_T_27 = 32'h3003 == _instType_T_6; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _instType_T_29 = 32'h4003 == _instType_T_6; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _instType_T_31 = 32'h5003 == _instType_T_6; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _instType_T_33 = 32'h6003 == _instType_T_6; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _instType_T_35 = 32'h23 == _instType_T_6; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _instType_T_37 = 32'h1023 == _instType_T_6; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _instType_T_39 = 32'h2023 == _instType_T_6; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _instType_T_41 = 32'h3023 == _instType_T_6; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _instType_T_43 = 32'h13 == _instType_T_6; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _instType_T_45 = 32'h2013 == _instType_T_6; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _instType_T_47 = 32'h3013 == _instType_T_6; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _instType_T_49 = 32'h4013 == _instType_T_6; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _instType_T_51 = 32'h6013 == _instType_T_6; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _instType_T_53 = 32'h7013 == _instType_T_6; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire [31:0] _instType_T_54 = io_if2id_inst & 32'hfc00707f; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _instType_T_55 = 32'h1013 == _instType_T_54; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _instType_T_57 = 32'h5013 == _instType_T_54; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _instType_T_59 = 32'h40005013 == _instType_T_54; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire [31:0] _instType_T_60 = io_if2id_inst & 32'hfe00707f; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _instType_T_61 = 32'h33 == _instType_T_60; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _instType_T_63 = 32'h40000033 == _instType_T_60; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _instType_T_65 = 32'h1033 == _instType_T_60; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _instType_T_67 = 32'h2033 == _instType_T_60; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _instType_T_69 = 32'h3033 == _instType_T_60; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _instType_T_71 = 32'h4033 == _instType_T_60; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _instType_T_73 = 32'h5033 == _instType_T_60; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _instType_T_75 = 32'h40005033 == _instType_T_60; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _instType_T_77 = 32'h6033 == _instType_T_60; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _instType_T_79 = 32'h7033 == _instType_T_60; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _instType_T_81 = 32'h2000033 == _instType_T_60; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _instType_T_83 = 32'h2001033 == _instType_T_60; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _instType_T_85 = 32'h2003033 == _instType_T_60; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _instType_T_87 = 32'h2002033 == _instType_T_60; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _instType_T_89 = 32'h2004033 == _instType_T_60; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _instType_T_91 = 32'h2005033 == _instType_T_60; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _instType_T_93 = 32'h2006033 == _instType_T_60; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _instType_T_95 = 32'h2007033 == _instType_T_60; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _instType_T_97 = 32'h200003b == _instType_T_60; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _instType_T_99 = 32'h200403b == _instType_T_60; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _instType_T_101 = 32'h200503b == _instType_T_60; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _instType_T_103 = 32'h200603b == _instType_T_60; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _instType_T_105 = 32'h200703b == _instType_T_60; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _instType_T_107 = 32'h1b == _instType_T_6; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _instType_T_109 = 32'h101b == _instType_T_60; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _instType_T_111 = 32'h501b == _instType_T_60; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _instType_T_113 = 32'h4000501b == _instType_T_60; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _instType_T_115 = 32'h3b == _instType_T_60; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _instType_T_117 = 32'h4000003b == _instType_T_60; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _instType_T_119 = 32'h103b == _instType_T_60; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _instType_T_121 = 32'h503b == _instType_T_60; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _instType_T_123 = 32'h4000503b == _instType_T_60; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _instType_T_125 = 32'h1073 == _instType_T_6; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _instType_T_127 = 32'h2073 == _instType_T_6; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _instType_T_129 = 32'h3073 == _instType_T_6; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _instType_T_131 = 32'h5073 == _instType_T_6; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _instType_T_133 = 32'h6073 == _instType_T_6; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _instType_T_135 = 32'h7073 == _instType_T_6; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire [31:0] _instType_T_136 = io_if2id_inst & 32'hf9f0707f; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _instType_T_137 = 32'h1000202f == _instType_T_136; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire [31:0] _instType_T_138 = io_if2id_inst & 32'hf800707f; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _instType_T_139 = 32'h1800202f == _instType_T_138; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _instType_T_141 = 32'h800202f == _instType_T_138; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _instType_T_143 = 32'h202f == _instType_T_138; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _instType_T_145 = 32'h2000202f == _instType_T_138; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _instType_T_147 = 32'h6000202f == _instType_T_138; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _instType_T_149 = 32'h4000202f == _instType_T_138; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _instType_T_151 = 32'h8000202f == _instType_T_138; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _instType_T_153 = 32'ha000202f == _instType_T_138; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _instType_T_155 = 32'hc000202f == _instType_T_138; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _instType_T_157 = 32'he000202f == _instType_T_138; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _instType_T_159 = 32'h1000302f == _instType_T_136; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _instType_T_161 = 32'h1800302f == _instType_T_138; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _instType_T_163 = 32'h800302f == _instType_T_138; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _instType_T_165 = 32'h302f == _instType_T_138; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _instType_T_167 = 32'h4000302f == _instType_T_138; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _instType_T_169 = 32'h2000302f == _instType_T_138; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _instType_T_171 = 32'h6000302f == _instType_T_138; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _instType_T_173 = 32'h8000302f == _instType_T_138; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _instType_T_175 = 32'ha000302f == _instType_T_138; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _instType_T_177 = 32'hc000302f == _instType_T_138; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _instType_T_179 = 32'he000302f == _instType_T_138; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire [31:0] _instType_T_180 = io_if2id_inst & 32'hf00fffff; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _instType_T_181 = 32'hf == _instType_T_180; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _instType_T_183 = 32'h100f == io_if2id_inst; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire [31:0] _instType_T_184 = io_if2id_inst & 32'hfe007fff; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _instType_T_185 = 32'h12000073 == _instType_T_184; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _instType_T_187 = 32'h10500073 == io_if2id_inst; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _instType_T_189 = 32'h6b == io_if2id_inst; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire [2:0] _instType_T_190 = _instType_T_189 ? 3'h0 : 3'h7; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _instType_T_191 = _instType_T_187 ? 3'h0 : _instType_T_190; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _instType_T_192 = _instType_T_185 ? 3'h0 : _instType_T_191; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _instType_T_193 = _instType_T_183 ? 3'h0 : _instType_T_192; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _instType_T_194 = _instType_T_181 ? 3'h0 : _instType_T_193; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _instType_T_195 = _instType_T_179 ? 3'h1 : _instType_T_194; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _instType_T_196 = _instType_T_177 ? 3'h1 : _instType_T_195; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _instType_T_197 = _instType_T_175 ? 3'h1 : _instType_T_196; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _instType_T_198 = _instType_T_173 ? 3'h1 : _instType_T_197; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _instType_T_199 = _instType_T_171 ? 3'h1 : _instType_T_198; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _instType_T_200 = _instType_T_169 ? 3'h1 : _instType_T_199; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _instType_T_201 = _instType_T_167 ? 3'h1 : _instType_T_200; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _instType_T_202 = _instType_T_165 ? 3'h1 : _instType_T_201; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _instType_T_203 = _instType_T_163 ? 3'h1 : _instType_T_202; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _instType_T_204 = _instType_T_161 ? 3'h1 : _instType_T_203; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _instType_T_205 = _instType_T_159 ? 3'h1 : _instType_T_204; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _instType_T_206 = _instType_T_157 ? 3'h1 : _instType_T_205; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _instType_T_207 = _instType_T_155 ? 3'h1 : _instType_T_206; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _instType_T_208 = _instType_T_153 ? 3'h1 : _instType_T_207; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _instType_T_209 = _instType_T_151 ? 3'h1 : _instType_T_208; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _instType_T_210 = _instType_T_149 ? 3'h1 : _instType_T_209; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _instType_T_211 = _instType_T_147 ? 3'h1 : _instType_T_210; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _instType_T_212 = _instType_T_145 ? 3'h1 : _instType_T_211; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _instType_T_213 = _instType_T_143 ? 3'h1 : _instType_T_212; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _instType_T_214 = _instType_T_141 ? 3'h1 : _instType_T_213; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _instType_T_215 = _instType_T_139 ? 3'h1 : _instType_T_214; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _instType_T_216 = _instType_T_137 ? 3'h1 : _instType_T_215; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _instType_T_217 = _instType_T_135 ? 3'h2 : _instType_T_216; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _instType_T_218 = _instType_T_133 ? 3'h2 : _instType_T_217; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _instType_T_219 = _instType_T_131 ? 3'h2 : _instType_T_218; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _instType_T_220 = _instType_T_129 ? 3'h2 : _instType_T_219; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _instType_T_221 = _instType_T_127 ? 3'h2 : _instType_T_220; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _instType_T_222 = _instType_T_125 ? 3'h2 : _instType_T_221; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _instType_T_223 = _instType_T_123 ? 3'h1 : _instType_T_222; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _instType_T_224 = _instType_T_121 ? 3'h1 : _instType_T_223; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _instType_T_225 = _instType_T_119 ? 3'h1 : _instType_T_224; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _instType_T_226 = _instType_T_117 ? 3'h1 : _instType_T_225; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _instType_T_227 = _instType_T_115 ? 3'h1 : _instType_T_226; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _instType_T_228 = _instType_T_113 ? 3'h2 : _instType_T_227; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _instType_T_229 = _instType_T_111 ? 3'h2 : _instType_T_228; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _instType_T_230 = _instType_T_109 ? 3'h2 : _instType_T_229; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _instType_T_231 = _instType_T_107 ? 3'h2 : _instType_T_230; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _instType_T_232 = _instType_T_105 ? 3'h1 : _instType_T_231; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _instType_T_233 = _instType_T_103 ? 3'h1 : _instType_T_232; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _instType_T_234 = _instType_T_101 ? 3'h1 : _instType_T_233; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _instType_T_235 = _instType_T_99 ? 3'h1 : _instType_T_234; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _instType_T_236 = _instType_T_97 ? 3'h1 : _instType_T_235; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _instType_T_237 = _instType_T_95 ? 3'h1 : _instType_T_236; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _instType_T_238 = _instType_T_93 ? 3'h1 : _instType_T_237; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _instType_T_239 = _instType_T_91 ? 3'h1 : _instType_T_238; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _instType_T_240 = _instType_T_89 ? 3'h1 : _instType_T_239; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _instType_T_241 = _instType_T_87 ? 3'h1 : _instType_T_240; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _instType_T_242 = _instType_T_85 ? 3'h1 : _instType_T_241; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _instType_T_243 = _instType_T_83 ? 3'h1 : _instType_T_242; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _instType_T_244 = _instType_T_81 ? 3'h1 : _instType_T_243; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _instType_T_245 = _instType_T_79 ? 3'h1 : _instType_T_244; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _instType_T_246 = _instType_T_77 ? 3'h1 : _instType_T_245; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _instType_T_247 = _instType_T_75 ? 3'h1 : _instType_T_246; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _instType_T_248 = _instType_T_73 ? 3'h1 : _instType_T_247; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _instType_T_249 = _instType_T_71 ? 3'h1 : _instType_T_248; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _instType_T_250 = _instType_T_69 ? 3'h1 : _instType_T_249; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _instType_T_251 = _instType_T_67 ? 3'h1 : _instType_T_250; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _instType_T_252 = _instType_T_65 ? 3'h1 : _instType_T_251; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _instType_T_253 = _instType_T_63 ? 3'h1 : _instType_T_252; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _instType_T_254 = _instType_T_61 ? 3'h1 : _instType_T_253; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _instType_T_255 = _instType_T_59 ? 3'h2 : _instType_T_254; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _instType_T_256 = _instType_T_57 ? 3'h2 : _instType_T_255; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _instType_T_257 = _instType_T_55 ? 3'h2 : _instType_T_256; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _instType_T_258 = _instType_T_53 ? 3'h2 : _instType_T_257; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _instType_T_259 = _instType_T_51 ? 3'h2 : _instType_T_258; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _instType_T_260 = _instType_T_49 ? 3'h2 : _instType_T_259; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _instType_T_261 = _instType_T_47 ? 3'h2 : _instType_T_260; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _instType_T_262 = _instType_T_45 ? 3'h2 : _instType_T_261; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _instType_T_263 = _instType_T_43 ? 3'h2 : _instType_T_262; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _instType_T_264 = _instType_T_41 ? 3'h3 : _instType_T_263; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _instType_T_265 = _instType_T_39 ? 3'h3 : _instType_T_264; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _instType_T_266 = _instType_T_37 ? 3'h3 : _instType_T_265; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _instType_T_267 = _instType_T_35 ? 3'h3 : _instType_T_266; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _instType_T_268 = _instType_T_33 ? 3'h2 : _instType_T_267; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _instType_T_269 = _instType_T_31 ? 3'h2 : _instType_T_268; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _instType_T_270 = _instType_T_29 ? 3'h2 : _instType_T_269; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _instType_T_271 = _instType_T_27 ? 3'h2 : _instType_T_270; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _instType_T_272 = _instType_T_25 ? 3'h2 : _instType_T_271; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _instType_T_273 = _instType_T_23 ? 3'h2 : _instType_T_272; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _instType_T_274 = _instType_T_21 ? 3'h2 : _instType_T_273; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _instType_T_275 = _instType_T_19 ? 3'h4 : _instType_T_274; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _instType_T_276 = _instType_T_17 ? 3'h4 : _instType_T_275; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _instType_T_277 = _instType_T_15 ? 3'h4 : _instType_T_276; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _instType_T_278 = _instType_T_13 ? 3'h4 : _instType_T_277; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _instType_T_279 = _instType_T_11 ? 3'h4 : _instType_T_278; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _instType_T_280 = _instType_T_9 ? 3'h4 : _instType_T_279; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _instType_T_281 = _instType_T_7 ? 3'h2 : _instType_T_280; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _instType_T_282 = _instType_T_5 ? 3'h6 : _instType_T_281; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _instType_T_283 = _instType_T_3 ? 3'h5 : _instType_T_282; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] instType_0 = _instType_T_1 ? 3'h5 : _instType_T_283; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_T_289 = _instType_T_179 ? 5'h1 : 5'h0; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_T_290 = _instType_T_177 ? 5'h1 : _instType_T_289; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_T_291 = _instType_T_175 ? 5'h1 : _instType_T_290; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_T_292 = _instType_T_173 ? 5'h1 : _instType_T_291; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_T_293 = _instType_T_171 ? 5'h1 : _instType_T_292; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_T_294 = _instType_T_169 ? 5'h1 : _instType_T_293; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_T_295 = _instType_T_167 ? 5'h1 : _instType_T_294; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_T_296 = _instType_T_165 ? 5'h1 : _instType_T_295; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_T_297 = _instType_T_163 ? 5'h1 : _instType_T_296; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_T_298 = _instType_T_161 ? 5'h1 : _instType_T_297; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_T_299 = _instType_T_159 ? 5'h1 : _instType_T_298; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_T_300 = _instType_T_157 ? 5'h1 : _instType_T_299; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_T_301 = _instType_T_155 ? 5'h1 : _instType_T_300; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_T_302 = _instType_T_153 ? 5'h1 : _instType_T_301; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_T_303 = _instType_T_151 ? 5'h1 : _instType_T_302; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_T_304 = _instType_T_149 ? 5'h1 : _instType_T_303; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_T_305 = _instType_T_147 ? 5'h1 : _instType_T_304; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_T_306 = _instType_T_145 ? 5'h1 : _instType_T_305; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_T_307 = _instType_T_143 ? 5'h1 : _instType_T_306; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_T_308 = _instType_T_141 ? 5'h1 : _instType_T_307; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_T_309 = _instType_T_139 ? 5'h1 : _instType_T_308; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_T_310 = _instType_T_137 ? 5'h1 : _instType_T_309; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_T_311 = _instType_T_135 ? 5'h15 : _instType_T_310; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_T_312 = _instType_T_133 ? 5'h5 : _instType_T_311; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_T_313 = _instType_T_131 ? 5'h1 : _instType_T_312; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_T_314 = _instType_T_129 ? 5'h15 : _instType_T_313; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_T_315 = _instType_T_127 ? 5'h5 : _instType_T_314; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_T_316 = _instType_T_125 ? 5'h1 : _instType_T_315; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_T_317 = _instType_T_123 ? 5'h9 : _instType_T_316; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_T_318 = _instType_T_121 ? 5'h8 : _instType_T_317; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_T_319 = _instType_T_119 ? 5'h7 : _instType_T_318; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_T_320 = _instType_T_117 ? 5'ha : _instType_T_319; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_T_321 = _instType_T_115 ? 5'h3 : _instType_T_320; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_T_322 = _instType_T_113 ? 5'h9 : _instType_T_321; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_T_323 = _instType_T_111 ? 5'h8 : _instType_T_322; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_T_324 = _instType_T_109 ? 5'h7 : _instType_T_323; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_T_325 = _instType_T_107 ? 5'h3 : _instType_T_324; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_T_326 = _instType_T_105 ? 5'h14 : _instType_T_325; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_T_327 = _instType_T_103 ? 5'h13 : _instType_T_326; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_T_328 = _instType_T_101 ? 5'h12 : _instType_T_327; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_T_329 = _instType_T_99 ? 5'h11 : _instType_T_328; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_T_330 = _instType_T_97 ? 5'hd : _instType_T_329; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_T_331 = _instType_T_95 ? 5'h14 : _instType_T_330; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_T_332 = _instType_T_93 ? 5'h13 : _instType_T_331; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_T_333 = _instType_T_91 ? 5'h12 : _instType_T_332; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_T_334 = _instType_T_89 ? 5'h11 : _instType_T_333; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_T_335 = _instType_T_87 ? 5'h10 : _instType_T_334; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_T_336 = _instType_T_85 ? 5'hf : _instType_T_335; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_T_337 = _instType_T_83 ? 5'he : _instType_T_336; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_T_338 = _instType_T_81 ? 5'hd : _instType_T_337; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_T_339 = _instType_T_79 ? 5'h6 : _instType_T_338; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_T_340 = _instType_T_77 ? 5'h5 : _instType_T_339; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_T_341 = _instType_T_75 ? 5'h9 : _instType_T_340; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_T_342 = _instType_T_73 ? 5'h8 : _instType_T_341; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_T_343 = _instType_T_71 ? 5'h4 : _instType_T_342; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_T_344 = _instType_T_69 ? 5'hc : _instType_T_343; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_T_345 = _instType_T_67 ? 5'hb : _instType_T_344; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_T_346 = _instType_T_65 ? 5'h7 : _instType_T_345; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_T_347 = _instType_T_63 ? 5'ha : _instType_T_346; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_T_348 = _instType_T_61 ? 5'h3 : _instType_T_347; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_T_349 = _instType_T_59 ? 5'h9 : _instType_T_348; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_T_350 = _instType_T_57 ? 5'h8 : _instType_T_349; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_T_351 = _instType_T_55 ? 5'h7 : _instType_T_350; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_T_352 = _instType_T_53 ? 5'h6 : _instType_T_351; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_T_353 = _instType_T_51 ? 5'h5 : _instType_T_352; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_T_354 = _instType_T_49 ? 5'h4 : _instType_T_353; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_T_355 = _instType_T_47 ? 5'hc : _instType_T_354; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_T_356 = _instType_T_45 ? 5'hb : _instType_T_355; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_T_357 = _instType_T_43 ? 5'h3 : _instType_T_356; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_T_358 = _instType_T_41 ? 5'h3 : _instType_T_357; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_T_359 = _instType_T_39 ? 5'h3 : _instType_T_358; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_T_360 = _instType_T_37 ? 5'h3 : _instType_T_359; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_T_361 = _instType_T_35 ? 5'h3 : _instType_T_360; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_T_362 = _instType_T_33 ? 5'h3 : _instType_T_361; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_T_363 = _instType_T_31 ? 5'h3 : _instType_T_362; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_T_364 = _instType_T_29 ? 5'h3 : _instType_T_363; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_T_365 = _instType_T_27 ? 5'h3 : _instType_T_364; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_T_366 = _instType_T_25 ? 5'h3 : _instType_T_365; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_T_367 = _instType_T_23 ? 5'h3 : _instType_T_366; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_T_368 = _instType_T_21 ? 5'h3 : _instType_T_367; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_T_369 = _instType_T_19 ? 5'h0 : _instType_T_368; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_T_370 = _instType_T_17 ? 5'h0 : _instType_T_369; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_T_371 = _instType_T_15 ? 5'h0 : _instType_T_370; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_T_372 = _instType_T_13 ? 5'h0 : _instType_T_371; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_T_373 = _instType_T_11 ? 5'h0 : _instType_T_372; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_T_374 = _instType_T_9 ? 5'h0 : _instType_T_373; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_T_375 = _instType_T_7 ? 5'h2 : _instType_T_374; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_T_376 = _instType_T_5 ? 5'h2 : _instType_T_375; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_T_377 = _instType_T_3 ? 5'h3 : _instType_T_376; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] instType_1 = _instType_T_1 ? 5'h1 : _instType_T_377; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_425 = _instType_T_95 ? 1'h0 : _instType_T_97 | (_instType_T_99 | (_instType_T_101 | (_instType_T_103
     | (_instType_T_105 | (_instType_T_107 | (_instType_T_109 | (_instType_T_111 | (_instType_T_113 | (_instType_T_115
     | (_instType_T_117 | (_instType_T_119 | (_instType_T_121 | _instType_T_123)))))))))))); // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_426 = _instType_T_93 ? 1'h0 : _instType_T_425; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_427 = _instType_T_91 ? 1'h0 : _instType_T_426; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_428 = _instType_T_89 ? 1'h0 : _instType_T_427; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_429 = _instType_T_87 ? 1'h0 : _instType_T_428; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_430 = _instType_T_85 ? 1'h0 : _instType_T_429; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_431 = _instType_T_83 ? 1'h0 : _instType_T_430; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_432 = _instType_T_81 ? 1'h0 : _instType_T_431; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_433 = _instType_T_79 ? 1'h0 : _instType_T_432; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_434 = _instType_T_77 ? 1'h0 : _instType_T_433; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_435 = _instType_T_75 ? 1'h0 : _instType_T_434; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_436 = _instType_T_73 ? 1'h0 : _instType_T_435; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_437 = _instType_T_71 ? 1'h0 : _instType_T_436; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_438 = _instType_T_69 ? 1'h0 : _instType_T_437; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_439 = _instType_T_67 ? 1'h0 : _instType_T_438; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_440 = _instType_T_65 ? 1'h0 : _instType_T_439; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_441 = _instType_T_63 ? 1'h0 : _instType_T_440; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_442 = _instType_T_61 ? 1'h0 : _instType_T_441; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_443 = _instType_T_59 ? 1'h0 : _instType_T_442; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_444 = _instType_T_57 ? 1'h0 : _instType_T_443; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_445 = _instType_T_55 ? 1'h0 : _instType_T_444; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_446 = _instType_T_53 ? 1'h0 : _instType_T_445; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_447 = _instType_T_51 ? 1'h0 : _instType_T_446; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_448 = _instType_T_49 ? 1'h0 : _instType_T_447; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_449 = _instType_T_47 ? 1'h0 : _instType_T_448; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_450 = _instType_T_45 ? 1'h0 : _instType_T_449; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_451 = _instType_T_43 ? 1'h0 : _instType_T_450; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_452 = _instType_T_41 ? 1'h0 : _instType_T_451; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_453 = _instType_T_39 ? 1'h0 : _instType_T_452; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_454 = _instType_T_37 ? 1'h0 : _instType_T_453; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_455 = _instType_T_35 ? 1'h0 : _instType_T_454; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_456 = _instType_T_33 ? 1'h0 : _instType_T_455; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_457 = _instType_T_31 ? 1'h0 : _instType_T_456; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_458 = _instType_T_29 ? 1'h0 : _instType_T_457; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_459 = _instType_T_27 ? 1'h0 : _instType_T_458; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_460 = _instType_T_25 ? 1'h0 : _instType_T_459; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_461 = _instType_T_23 ? 1'h0 : _instType_T_460; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_462 = _instType_T_21 ? 1'h0 : _instType_T_461; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_463 = _instType_T_19 ? 1'h0 : _instType_T_462; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_464 = _instType_T_17 ? 1'h0 : _instType_T_463; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_465 = _instType_T_15 ? 1'h0 : _instType_T_464; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_466 = _instType_T_13 ? 1'h0 : _instType_T_465; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_467 = _instType_T_11 ? 1'h0 : _instType_T_466; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_468 = _instType_T_9 ? 1'h0 : _instType_T_467; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_469 = _instType_T_7 ? 1'h0 : _instType_T_468; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_470 = _instType_T_5 ? 1'h0 : _instType_T_469; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_471 = _instType_T_3 ? 1'h0 : _instType_T_470; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  instType_2 = _instType_T_1 ? 1'h0 : _instType_T_471; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_T_477 = _instType_T_179 ? 5'hf : 5'h0; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_T_478 = _instType_T_177 ? 5'hf : _instType_T_477; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_T_479 = _instType_T_175 ? 5'hf : _instType_T_478; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_T_480 = _instType_T_173 ? 5'hf : _instType_T_479; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_T_481 = _instType_T_171 ? 5'hf : _instType_T_480; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_T_482 = _instType_T_169 ? 5'hf : _instType_T_481; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_T_483 = _instType_T_167 ? 5'hf : _instType_T_482; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_T_484 = _instType_T_165 ? 5'hf : _instType_T_483; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_T_485 = _instType_T_163 ? 5'hf : _instType_T_484; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_T_486 = _instType_T_161 ? 5'hb : _instType_T_485; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_T_487 = _instType_T_159 ? 5'h7 : _instType_T_486; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_T_488 = _instType_T_157 ? 5'he : _instType_T_487; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_T_489 = _instType_T_155 ? 5'he : _instType_T_488; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_T_490 = _instType_T_153 ? 5'he : _instType_T_489; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_T_491 = _instType_T_151 ? 5'he : _instType_T_490; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_T_492 = _instType_T_149 ? 5'he : _instType_T_491; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_T_493 = _instType_T_147 ? 5'he : _instType_T_492; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_T_494 = _instType_T_145 ? 5'he : _instType_T_493; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_T_495 = _instType_T_143 ? 5'he : _instType_T_494; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_T_496 = _instType_T_141 ? 5'he : _instType_T_495; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_T_497 = _instType_T_139 ? 5'ha : _instType_T_496; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_T_498 = _instType_T_137 ? 5'h6 : _instType_T_497; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_T_499 = _instType_T_135 ? 5'h0 : _instType_T_498; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_T_500 = _instType_T_133 ? 5'h0 : _instType_T_499; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_T_501 = _instType_T_131 ? 5'h0 : _instType_T_500; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_T_502 = _instType_T_129 ? 5'h0 : _instType_T_501; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_T_503 = _instType_T_127 ? 5'h0 : _instType_T_502; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_T_504 = _instType_T_125 ? 5'h0 : _instType_T_503; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_T_505 = _instType_T_123 ? 5'h0 : _instType_T_504; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_T_506 = _instType_T_121 ? 5'h0 : _instType_T_505; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_T_507 = _instType_T_119 ? 5'h0 : _instType_T_506; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_T_508 = _instType_T_117 ? 5'h0 : _instType_T_507; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_T_509 = _instType_T_115 ? 5'h0 : _instType_T_508; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_T_510 = _instType_T_113 ? 5'h0 : _instType_T_509; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_T_511 = _instType_T_111 ? 5'h0 : _instType_T_510; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_T_512 = _instType_T_109 ? 5'h0 : _instType_T_511; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_T_513 = _instType_T_107 ? 5'h0 : _instType_T_512; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_T_514 = _instType_T_105 ? 5'h0 : _instType_T_513; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_T_515 = _instType_T_103 ? 5'h0 : _instType_T_514; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_T_516 = _instType_T_101 ? 5'h0 : _instType_T_515; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_T_517 = _instType_T_99 ? 5'h0 : _instType_T_516; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_T_518 = _instType_T_97 ? 5'h0 : _instType_T_517; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_T_519 = _instType_T_95 ? 5'h0 : _instType_T_518; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_T_520 = _instType_T_93 ? 5'h0 : _instType_T_519; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_T_521 = _instType_T_91 ? 5'h0 : _instType_T_520; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_T_522 = _instType_T_89 ? 5'h0 : _instType_T_521; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_T_523 = _instType_T_87 ? 5'h0 : _instType_T_522; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_T_524 = _instType_T_85 ? 5'h0 : _instType_T_523; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_T_525 = _instType_T_83 ? 5'h0 : _instType_T_524; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_T_526 = _instType_T_81 ? 5'h0 : _instType_T_525; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_T_527 = _instType_T_79 ? 5'h0 : _instType_T_526; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_T_528 = _instType_T_77 ? 5'h0 : _instType_T_527; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_T_529 = _instType_T_75 ? 5'h0 : _instType_T_528; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_T_530 = _instType_T_73 ? 5'h0 : _instType_T_529; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_T_531 = _instType_T_71 ? 5'h0 : _instType_T_530; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_T_532 = _instType_T_69 ? 5'h0 : _instType_T_531; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_T_533 = _instType_T_67 ? 5'h0 : _instType_T_532; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_T_534 = _instType_T_65 ? 5'h0 : _instType_T_533; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_T_535 = _instType_T_63 ? 5'h0 : _instType_T_534; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_T_536 = _instType_T_61 ? 5'h0 : _instType_T_535; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_T_537 = _instType_T_59 ? 5'h0 : _instType_T_536; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_T_538 = _instType_T_57 ? 5'h0 : _instType_T_537; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_T_539 = _instType_T_55 ? 5'h0 : _instType_T_538; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_T_540 = _instType_T_53 ? 5'h0 : _instType_T_539; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_T_541 = _instType_T_51 ? 5'h0 : _instType_T_540; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_T_542 = _instType_T_49 ? 5'h0 : _instType_T_541; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_T_543 = _instType_T_47 ? 5'h0 : _instType_T_542; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_T_544 = _instType_T_45 ? 5'h0 : _instType_T_543; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_T_545 = _instType_T_43 ? 5'h0 : _instType_T_544; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_T_546 = _instType_T_41 ? 5'hb : _instType_T_545; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_T_547 = _instType_T_39 ? 5'ha : _instType_T_546; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_T_548 = _instType_T_37 ? 5'h9 : _instType_T_547; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_T_549 = _instType_T_35 ? 5'h8 : _instType_T_548; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_T_550 = _instType_T_33 ? 5'h16 : _instType_T_549; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_T_551 = _instType_T_31 ? 5'h15 : _instType_T_550; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_T_552 = _instType_T_29 ? 5'h14 : _instType_T_551; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_T_553 = _instType_T_27 ? 5'h7 : _instType_T_552; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_T_554 = _instType_T_25 ? 5'h6 : _instType_T_553; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_T_555 = _instType_T_23 ? 5'h5 : _instType_T_554; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_T_556 = _instType_T_21 ? 5'h4 : _instType_T_555; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_T_557 = _instType_T_19 ? 5'h0 : _instType_T_556; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_T_558 = _instType_T_17 ? 5'h0 : _instType_T_557; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_T_559 = _instType_T_15 ? 5'h0 : _instType_T_558; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_T_560 = _instType_T_13 ? 5'h0 : _instType_T_559; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_T_561 = _instType_T_11 ? 5'h0 : _instType_T_560; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_T_562 = _instType_T_9 ? 5'h0 : _instType_T_561; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_T_563 = _instType_T_7 ? 5'h0 : _instType_T_562; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_T_564 = _instType_T_5 ? 5'h0 : _instType_T_563; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_T_565 = _instType_T_3 ? 5'h0 : _instType_T_564; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] instType_3 = _instType_T_1 ? 5'h0 : _instType_T_565; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_601 = _instType_T_119 | (_instType_T_121 | (_instType_T_123 | (_instType_T_125 | (_instType_T_127 |
    (_instType_T_129 | (_instType_T_131 | (_instType_T_133 | (_instType_T_135 | (_instType_T_137 | (_instType_T_139 | (
    _instType_T_141 | (_instType_T_143 | (_instType_T_145 | (_instType_T_147 | (_instType_T_149 | (_instType_T_151 | (
    _instType_T_153 | (_instType_T_155 | (_instType_T_157 | (_instType_T_159 | (_instType_T_161 | (_instType_T_163 | (
    _instType_T_165 | (_instType_T_167 | (_instType_T_169 | (_instType_T_171 | (_instType_T_173 | (_instType_T_175 | (
    _instType_T_177 | _instType_T_179))))))))))))))))))))))))))))); // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_631 = _instType_T_59 | (_instType_T_61 | (_instType_T_63 | (_instType_T_65 | (_instType_T_67 | (
    _instType_T_69 | (_instType_T_71 | (_instType_T_73 | (_instType_T_75 | (_instType_T_77 | (_instType_T_79 | (
    _instType_T_81 | (_instType_T_83 | (_instType_T_85 | (_instType_T_87 | (_instType_T_89 | (_instType_T_91 | (
    _instType_T_93 | (_instType_T_95 | (_instType_T_97 | (_instType_T_99 | (_instType_T_101 | (_instType_T_103 | (
    _instType_T_105 | (_instType_T_107 | (_instType_T_109 | (_instType_T_111 | (_instType_T_113 | (_instType_T_115 | (
    _instType_T_117 | _instType_T_601))))))))))))))))))))))))))))); // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_640 = _instType_T_41 ? 1'h0 : _instType_T_43 | (_instType_T_45 | (_instType_T_47 | (_instType_T_49
     | (_instType_T_51 | (_instType_T_53 | (_instType_T_55 | (_instType_T_57 | _instType_T_631))))))); // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_641 = _instType_T_39 ? 1'h0 : _instType_T_640; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_642 = _instType_T_37 ? 1'h0 : _instType_T_641; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_643 = _instType_T_35 ? 1'h0 : _instType_T_642; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_651 = _instType_T_19 ? 1'h0 : _instType_T_21 | (_instType_T_23 | (_instType_T_25 | (_instType_T_27
     | (_instType_T_29 | (_instType_T_31 | (_instType_T_33 | _instType_T_643)))))); // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_652 = _instType_T_17 ? 1'h0 : _instType_T_651; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_653 = _instType_T_15 ? 1'h0 : _instType_T_652; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_654 = _instType_T_13 ? 1'h0 : _instType_T_653; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_655 = _instType_T_11 ? 1'h0 : _instType_T_654; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_656 = _instType_T_9 ? 1'h0 : _instType_T_655; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  instType_4 = _instType_T_1 | (_instType_T_3 | (_instType_T_5 | (_instType_T_7 | _instType_T_656))); // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_753 = _instType_T_3 ? 1'h0 : _instType_T_5 | (_instType_T_7 | (_instType_T_9 | (_instType_T_11 | (
    _instType_T_13 | (_instType_T_15 | (_instType_T_17 | _instType_T_19)))))); // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  instType_5 = _instType_T_1 ? 1'h0 : _instType_T_753; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_787 = _instType_T_123 ? 1'h0 : _instType_T_125 | (_instType_T_127 | (_instType_T_129 | (
    _instType_T_131 | (_instType_T_133 | _instType_T_135)))); // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_788 = _instType_T_121 ? 1'h0 : _instType_T_787; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_789 = _instType_T_119 ? 1'h0 : _instType_T_788; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_790 = _instType_T_117 ? 1'h0 : _instType_T_789; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_791 = _instType_T_115 ? 1'h0 : _instType_T_790; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_792 = _instType_T_113 ? 1'h0 : _instType_T_791; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_793 = _instType_T_111 ? 1'h0 : _instType_T_792; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_794 = _instType_T_109 ? 1'h0 : _instType_T_793; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_795 = _instType_T_107 ? 1'h0 : _instType_T_794; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_796 = _instType_T_105 ? 1'h0 : _instType_T_795; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_797 = _instType_T_103 ? 1'h0 : _instType_T_796; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_798 = _instType_T_101 ? 1'h0 : _instType_T_797; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_799 = _instType_T_99 ? 1'h0 : _instType_T_798; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_800 = _instType_T_97 ? 1'h0 : _instType_T_799; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_801 = _instType_T_95 ? 1'h0 : _instType_T_800; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_802 = _instType_T_93 ? 1'h0 : _instType_T_801; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_803 = _instType_T_91 ? 1'h0 : _instType_T_802; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_804 = _instType_T_89 ? 1'h0 : _instType_T_803; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_805 = _instType_T_87 ? 1'h0 : _instType_T_804; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_806 = _instType_T_85 ? 1'h0 : _instType_T_805; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_807 = _instType_T_83 ? 1'h0 : _instType_T_806; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_808 = _instType_T_81 ? 1'h0 : _instType_T_807; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_809 = _instType_T_79 ? 1'h0 : _instType_T_808; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_810 = _instType_T_77 ? 1'h0 : _instType_T_809; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_811 = _instType_T_75 ? 1'h0 : _instType_T_810; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_812 = _instType_T_73 ? 1'h0 : _instType_T_811; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_813 = _instType_T_71 ? 1'h0 : _instType_T_812; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_814 = _instType_T_69 ? 1'h0 : _instType_T_813; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_815 = _instType_T_67 ? 1'h0 : _instType_T_814; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_816 = _instType_T_65 ? 1'h0 : _instType_T_815; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_817 = _instType_T_63 ? 1'h0 : _instType_T_816; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_818 = _instType_T_61 ? 1'h0 : _instType_T_817; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_819 = _instType_T_59 ? 1'h0 : _instType_T_818; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_820 = _instType_T_57 ? 1'h0 : _instType_T_819; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_821 = _instType_T_55 ? 1'h0 : _instType_T_820; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_822 = _instType_T_53 ? 1'h0 : _instType_T_821; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_823 = _instType_T_51 ? 1'h0 : _instType_T_822; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_824 = _instType_T_49 ? 1'h0 : _instType_T_823; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_825 = _instType_T_47 ? 1'h0 : _instType_T_824; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_826 = _instType_T_45 ? 1'h0 : _instType_T_825; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_827 = _instType_T_43 ? 1'h0 : _instType_T_826; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_828 = _instType_T_41 ? 1'h0 : _instType_T_827; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_829 = _instType_T_39 ? 1'h0 : _instType_T_828; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_830 = _instType_T_37 ? 1'h0 : _instType_T_829; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_831 = _instType_T_35 ? 1'h0 : _instType_T_830; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_832 = _instType_T_33 ? 1'h0 : _instType_T_831; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_833 = _instType_T_31 ? 1'h0 : _instType_T_832; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_834 = _instType_T_29 ? 1'h0 : _instType_T_833; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_835 = _instType_T_27 ? 1'h0 : _instType_T_834; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_836 = _instType_T_25 ? 1'h0 : _instType_T_835; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_837 = _instType_T_23 ? 1'h0 : _instType_T_836; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_838 = _instType_T_21 ? 1'h0 : _instType_T_837; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_839 = _instType_T_19 ? 1'h0 : _instType_T_838; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_840 = _instType_T_17 ? 1'h0 : _instType_T_839; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_841 = _instType_T_15 ? 1'h0 : _instType_T_840; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_842 = _instType_T_13 ? 1'h0 : _instType_T_841; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_843 = _instType_T_11 ? 1'h0 : _instType_T_842; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_844 = _instType_T_9 ? 1'h0 : _instType_T_843; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_845 = _instType_T_7 ? 1'h0 : _instType_T_844; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_846 = _instType_T_5 ? 1'h0 : _instType_T_845; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_847 = _instType_T_3 ? 1'h0 : _instType_T_846; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  instType_6 = _instType_T_1 ? 1'h0 : _instType_T_847; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_972 = _instType_T_129 ? 1'h0 : _instType_T_131 | (_instType_T_133 | _instType_T_135); // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_973 = _instType_T_127 ? 1'h0 : _instType_T_972; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_974 = _instType_T_125 ? 1'h0 : _instType_T_973; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_975 = _instType_T_123 ? 1'h0 : _instType_T_974; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_976 = _instType_T_121 ? 1'h0 : _instType_T_975; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_977 = _instType_T_119 ? 1'h0 : _instType_T_976; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_978 = _instType_T_117 ? 1'h0 : _instType_T_977; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_979 = _instType_T_115 ? 1'h0 : _instType_T_978; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_980 = _instType_T_113 ? 1'h0 : _instType_T_979; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_981 = _instType_T_111 ? 1'h0 : _instType_T_980; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_982 = _instType_T_109 ? 1'h0 : _instType_T_981; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_983 = _instType_T_107 ? 1'h0 : _instType_T_982; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_984 = _instType_T_105 ? 1'h0 : _instType_T_983; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_985 = _instType_T_103 ? 1'h0 : _instType_T_984; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_986 = _instType_T_101 ? 1'h0 : _instType_T_985; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_987 = _instType_T_99 ? 1'h0 : _instType_T_986; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_988 = _instType_T_97 ? 1'h0 : _instType_T_987; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_989 = _instType_T_95 ? 1'h0 : _instType_T_988; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_990 = _instType_T_93 ? 1'h0 : _instType_T_989; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_991 = _instType_T_91 ? 1'h0 : _instType_T_990; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_992 = _instType_T_89 ? 1'h0 : _instType_T_991; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_993 = _instType_T_87 ? 1'h0 : _instType_T_992; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_994 = _instType_T_85 ? 1'h0 : _instType_T_993; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_995 = _instType_T_83 ? 1'h0 : _instType_T_994; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_996 = _instType_T_81 ? 1'h0 : _instType_T_995; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_997 = _instType_T_79 ? 1'h0 : _instType_T_996; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_998 = _instType_T_77 ? 1'h0 : _instType_T_997; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_999 = _instType_T_75 ? 1'h0 : _instType_T_998; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_1000 = _instType_T_73 ? 1'h0 : _instType_T_999; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_1001 = _instType_T_71 ? 1'h0 : _instType_T_1000; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_1002 = _instType_T_69 ? 1'h0 : _instType_T_1001; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_1003 = _instType_T_67 ? 1'h0 : _instType_T_1002; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_1004 = _instType_T_65 ? 1'h0 : _instType_T_1003; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_1005 = _instType_T_63 ? 1'h0 : _instType_T_1004; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_1006 = _instType_T_61 ? 1'h0 : _instType_T_1005; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_1007 = _instType_T_59 ? 1'h0 : _instType_T_1006; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_1008 = _instType_T_57 ? 1'h0 : _instType_T_1007; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_1009 = _instType_T_55 ? 1'h0 : _instType_T_1008; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_1010 = _instType_T_53 ? 1'h0 : _instType_T_1009; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_1011 = _instType_T_51 ? 1'h0 : _instType_T_1010; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_1012 = _instType_T_49 ? 1'h0 : _instType_T_1011; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_1013 = _instType_T_47 ? 1'h0 : _instType_T_1012; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_1014 = _instType_T_45 ? 1'h0 : _instType_T_1013; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_1015 = _instType_T_43 ? 1'h0 : _instType_T_1014; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_1016 = _instType_T_41 ? 1'h0 : _instType_T_1015; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_1017 = _instType_T_39 ? 1'h0 : _instType_T_1016; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_1018 = _instType_T_37 ? 1'h0 : _instType_T_1017; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_1019 = _instType_T_35 ? 1'h0 : _instType_T_1018; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_1020 = _instType_T_33 ? 1'h0 : _instType_T_1019; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_1021 = _instType_T_31 ? 1'h0 : _instType_T_1020; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_1022 = _instType_T_29 ? 1'h0 : _instType_T_1021; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_1023 = _instType_T_27 ? 1'h0 : _instType_T_1022; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_1024 = _instType_T_25 ? 1'h0 : _instType_T_1023; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_1025 = _instType_T_23 ? 1'h0 : _instType_T_1024; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_1026 = _instType_T_21 ? 1'h0 : _instType_T_1025; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_1027 = _instType_T_19 ? 1'h0 : _instType_T_1026; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_1028 = _instType_T_17 ? 1'h0 : _instType_T_1027; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_1029 = _instType_T_15 ? 1'h0 : _instType_T_1028; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_1030 = _instType_T_13 ? 1'h0 : _instType_T_1029; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_1031 = _instType_T_11 ? 1'h0 : _instType_T_1030; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_1032 = _instType_T_9 ? 1'h0 : _instType_T_1031; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_1033 = _instType_T_7 ? 1'h0 : _instType_T_1032; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_1034 = _instType_T_5 ? 1'h0 : _instType_T_1033; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_T_1035 = _instType_T_3 ? 1'h0 : _instType_T_1034; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  instType_8 = _instType_T_1 ? 1'h0 : _instType_T_1035; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [15:0] _instType_c_T_1 = io_if2id_inst[15:0] & 16'he003; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _instType_c_T_2 = 16'h0 == _instType_c_T_1; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _instType_c_T_4 = 16'h4000 == _instType_c_T_1; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _instType_c_T_6 = 16'h6000 == _instType_c_T_1; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _instType_c_T_8 = 16'hc000 == _instType_c_T_1; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _instType_c_T_10 = 16'he000 == _instType_c_T_1; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _instType_c_T_12 = 16'h1 == _instType_c_T_1; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _instType_c_T_14 = 16'h2001 == _instType_c_T_1; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _instType_c_T_16 = 16'h4001 == _instType_c_T_1; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire [15:0] _instType_c_T_17 = io_if2id_inst[15:0] & 16'hef83; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _instType_c_T_18 = 16'h6101 == _instType_c_T_17; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _instType_c_T_20 = 16'h6001 == _instType_c_T_1; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire [15:0] _instType_c_T_21 = io_if2id_inst[15:0] & 16'hec03; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _instType_c_T_22 = 16'h8001 == _instType_c_T_21; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _instType_c_T_24 = 16'h8401 == _instType_c_T_21; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _instType_c_T_26 = 16'h8801 == _instType_c_T_21; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire [15:0] _instType_c_T_27 = io_if2id_inst[15:0] & 16'hfc63; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _instType_c_T_28 = 16'h8c01 == _instType_c_T_27; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _instType_c_T_30 = 16'h8c21 == _instType_c_T_27; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _instType_c_T_32 = 16'h8c41 == _instType_c_T_27; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _instType_c_T_34 = 16'h8c61 == _instType_c_T_27; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _instType_c_T_36 = 16'h9c01 == _instType_c_T_27; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _instType_c_T_38 = 16'h9c21 == _instType_c_T_27; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _instType_c_T_40 = 16'ha001 == _instType_c_T_1; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _instType_c_T_42 = 16'hc001 == _instType_c_T_1; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _instType_c_T_44 = 16'he001 == _instType_c_T_1; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _instType_c_T_46 = 16'h2 == _instType_c_T_1; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _instType_c_T_48 = 16'h4002 == _instType_c_T_1; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _instType_c_T_50 = 16'h6002 == _instType_c_T_1; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire [15:0] _instType_c_T_51 = io_if2id_inst[15:0] & 16'hf07f; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _instType_c_T_52 = 16'h8002 == _instType_c_T_51; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire [15:0] _instType_c_T_53 = io_if2id_inst[15:0] & 16'hf003; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _instType_c_T_54 = 16'h8002 == _instType_c_T_53; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _instType_c_T_56 = 16'h9002 == _instType_c_T_51; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _instType_c_T_58 = 16'h9002 == _instType_c_T_53; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _instType_c_T_60 = 16'hc002 == _instType_c_T_1; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _instType_c_T_62 = 16'he002 == _instType_c_T_1; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire [3:0] _instType_c_T_63 = _instType_c_T_62 ? 4'h3 : 4'h0; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _instType_c_T_64 = _instType_c_T_60 ? 4'h3 : _instType_c_T_63; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _instType_c_T_65 = _instType_c_T_58 ? 4'h1 : _instType_c_T_64; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _instType_c_T_66 = _instType_c_T_56 ? 4'h1 : _instType_c_T_65; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _instType_c_T_67 = _instType_c_T_54 ? 4'h1 : _instType_c_T_66; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _instType_c_T_68 = _instType_c_T_52 ? 4'h1 : _instType_c_T_67; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _instType_c_T_69 = _instType_c_T_50 ? 4'h2 : _instType_c_T_68; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _instType_c_T_70 = _instType_c_T_48 ? 4'h2 : _instType_c_T_69; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _instType_c_T_71 = _instType_c_T_46 ? 4'h2 : _instType_c_T_70; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _instType_c_T_72 = _instType_c_T_44 ? 4'h7 : _instType_c_T_71; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _instType_c_T_73 = _instType_c_T_42 ? 4'h7 : _instType_c_T_72; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _instType_c_T_74 = _instType_c_T_40 ? 4'h8 : _instType_c_T_73; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _instType_c_T_75 = _instType_c_T_38 ? 4'h6 : _instType_c_T_74; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _instType_c_T_76 = _instType_c_T_36 ? 4'h6 : _instType_c_T_75; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _instType_c_T_77 = _instType_c_T_34 ? 4'h6 : _instType_c_T_76; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _instType_c_T_78 = _instType_c_T_32 ? 4'h6 : _instType_c_T_77; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _instType_c_T_79 = _instType_c_T_30 ? 4'h6 : _instType_c_T_78; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _instType_c_T_80 = _instType_c_T_28 ? 4'h6 : _instType_c_T_79; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _instType_c_T_81 = _instType_c_T_26 ? 4'h7 : _instType_c_T_80; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _instType_c_T_82 = _instType_c_T_24 ? 4'h7 : _instType_c_T_81; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _instType_c_T_83 = _instType_c_T_22 ? 4'h7 : _instType_c_T_82; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _instType_c_T_84 = _instType_c_T_20 ? 4'h2 : _instType_c_T_83; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _instType_c_T_85 = _instType_c_T_18 ? 4'h2 : _instType_c_T_84; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _instType_c_T_86 = _instType_c_T_16 ? 4'h2 : _instType_c_T_85; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _instType_c_T_87 = _instType_c_T_14 ? 4'h2 : _instType_c_T_86; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _instType_c_T_88 = _instType_c_T_12 ? 4'h2 : _instType_c_T_87; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _instType_c_T_89 = _instType_c_T_10 ? 4'h6 : _instType_c_T_88; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _instType_c_T_90 = _instType_c_T_8 ? 4'h6 : _instType_c_T_89; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _instType_c_T_91 = _instType_c_T_6 ? 4'h5 : _instType_c_T_90; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _instType_c_T_92 = _instType_c_T_4 ? 4'h5 : _instType_c_T_91; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] instType_c_0 = _instType_c_T_2 ? 4'h4 : _instType_c_T_92; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _instType_c_T_93 = _instType_c_T_62 ? 4'hd : 4'h0; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _instType_c_T_94 = _instType_c_T_60 ? 4'hc : _instType_c_T_93; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _instType_c_T_95 = _instType_c_T_58 ? 4'h0 : _instType_c_T_94; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _instType_c_T_96 = _instType_c_T_56 ? 4'h0 : _instType_c_T_95; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _instType_c_T_97 = _instType_c_T_54 ? 4'h0 : _instType_c_T_96; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _instType_c_T_98 = _instType_c_T_52 ? 4'h0 : _instType_c_T_97; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _instType_c_T_99 = _instType_c_T_50 ? 4'h7 : _instType_c_T_98; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _instType_c_T_100 = _instType_c_T_48 ? 4'h6 : _instType_c_T_99; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _instType_c_T_101 = _instType_c_T_46 ? 4'h4 : _instType_c_T_100; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _instType_c_T_102 = _instType_c_T_44 ? 4'hb : _instType_c_T_101; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _instType_c_T_103 = _instType_c_T_42 ? 4'hb : _instType_c_T_102; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _instType_c_T_104 = _instType_c_T_40 ? 4'ha : _instType_c_T_103; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _instType_c_T_105 = _instType_c_T_38 ? 4'h0 : _instType_c_T_104; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _instType_c_T_106 = _instType_c_T_36 ? 4'h0 : _instType_c_T_105; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _instType_c_T_107 = _instType_c_T_34 ? 4'h0 : _instType_c_T_106; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _instType_c_T_108 = _instType_c_T_32 ? 4'h0 : _instType_c_T_107; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _instType_c_T_109 = _instType_c_T_30 ? 4'h0 : _instType_c_T_108; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _instType_c_T_110 = _instType_c_T_28 ? 4'h0 : _instType_c_T_109; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _instType_c_T_111 = _instType_c_T_26 ? 4'h5 : _instType_c_T_110; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _instType_c_T_112 = _instType_c_T_24 ? 4'h4 : _instType_c_T_111; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _instType_c_T_113 = _instType_c_T_22 ? 4'h4 : _instType_c_T_112; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _instType_c_T_114 = _instType_c_T_20 ? 4'h9 : _instType_c_T_113; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _instType_c_T_115 = _instType_c_T_18 ? 4'h8 : _instType_c_T_114; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _instType_c_T_116 = _instType_c_T_16 ? 4'h5 : _instType_c_T_115; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _instType_c_T_117 = _instType_c_T_14 ? 4'h5 : _instType_c_T_116; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _instType_c_T_118 = _instType_c_T_12 ? 4'h5 : _instType_c_T_117; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _instType_c_T_119 = _instType_c_T_10 ? 4'h3 : _instType_c_T_118; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _instType_c_T_120 = _instType_c_T_8 ? 4'h2 : _instType_c_T_119; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _instType_c_T_121 = _instType_c_T_6 ? 4'h3 : _instType_c_T_120; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _instType_c_T_122 = _instType_c_T_4 ? 4'h2 : _instType_c_T_121; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] instType_c_1 = _instType_c_T_2 ? 4'h1 : _instType_c_T_122; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_c_T_123 = _instType_c_T_62 ? 5'h3 : 5'h0; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_c_T_124 = _instType_c_T_60 ? 5'h3 : _instType_c_T_123; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_c_T_125 = _instType_c_T_58 ? 5'h3 : _instType_c_T_124; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_c_T_126 = _instType_c_T_56 ? 5'h2 : _instType_c_T_125; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_c_T_127 = _instType_c_T_54 ? 5'h2 : _instType_c_T_126; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_c_T_128 = _instType_c_T_52 ? 5'h1 : _instType_c_T_127; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_c_T_129 = _instType_c_T_50 ? 5'h3 : _instType_c_T_128; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_c_T_130 = _instType_c_T_48 ? 5'h3 : _instType_c_T_129; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_c_T_131 = _instType_c_T_46 ? 5'h7 : _instType_c_T_130; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_c_T_132 = _instType_c_T_44 ? 5'h0 : _instType_c_T_131; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_c_T_133 = _instType_c_T_42 ? 5'h0 : _instType_c_T_132; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_c_T_134 = _instType_c_T_40 ? 5'h2 : _instType_c_T_133; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_c_T_135 = _instType_c_T_38 ? 5'h3 : _instType_c_T_134; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_c_T_136 = _instType_c_T_36 ? 5'ha : _instType_c_T_135; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_c_T_137 = _instType_c_T_34 ? 5'h6 : _instType_c_T_136; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_c_T_138 = _instType_c_T_32 ? 5'h5 : _instType_c_T_137; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_c_T_139 = _instType_c_T_30 ? 5'h4 : _instType_c_T_138; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_c_T_140 = _instType_c_T_28 ? 5'ha : _instType_c_T_139; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_c_T_141 = _instType_c_T_26 ? 5'h6 : _instType_c_T_140; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_c_T_142 = _instType_c_T_24 ? 5'h9 : _instType_c_T_141; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_c_T_143 = _instType_c_T_22 ? 5'h8 : _instType_c_T_142; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_c_T_144 = _instType_c_T_20 ? 5'h2 : _instType_c_T_143; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_c_T_145 = _instType_c_T_18 ? 5'h3 : _instType_c_T_144; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_c_T_146 = _instType_c_T_16 ? 5'h2 : _instType_c_T_145; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_c_T_147 = _instType_c_T_14 ? 5'h3 : _instType_c_T_146; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_c_T_148 = _instType_c_T_12 ? 5'h3 : _instType_c_T_147; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_c_T_149 = _instType_c_T_10 ? 5'h3 : _instType_c_T_148; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_c_T_150 = _instType_c_T_8 ? 5'h3 : _instType_c_T_149; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_c_T_151 = _instType_c_T_6 ? 5'h3 : _instType_c_T_150; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_c_T_152 = _instType_c_T_4 ? 5'h3 : _instType_c_T_151; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_c_T_167 = _instType_c_T_34 ? 1'h0 : _instType_c_T_36 | _instType_c_T_38; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_c_T_168 = _instType_c_T_32 ? 1'h0 : _instType_c_T_167; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_c_T_169 = _instType_c_T_30 ? 1'h0 : _instType_c_T_168; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_c_T_170 = _instType_c_T_28 ? 1'h0 : _instType_c_T_169; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_c_T_171 = _instType_c_T_26 ? 1'h0 : _instType_c_T_170; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_c_T_172 = _instType_c_T_24 ? 1'h0 : _instType_c_T_171; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_c_T_173 = _instType_c_T_22 ? 1'h0 : _instType_c_T_172; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_c_T_174 = _instType_c_T_20 ? 1'h0 : _instType_c_T_173; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_c_T_175 = _instType_c_T_18 ? 1'h0 : _instType_c_T_174; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_c_T_176 = _instType_c_T_16 ? 1'h0 : _instType_c_T_175; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_c_T_178 = _instType_c_T_12 ? 1'h0 : _instType_c_T_14 | _instType_c_T_176; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_c_T_179 = _instType_c_T_10 ? 1'h0 : _instType_c_T_178; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_c_T_180 = _instType_c_T_8 ? 1'h0 : _instType_c_T_179; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_c_T_181 = _instType_c_T_6 ? 1'h0 : _instType_c_T_180; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_c_T_182 = _instType_c_T_4 ? 1'h0 : _instType_c_T_181; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_c_T_183 = _instType_c_T_62 ? 5'hb : 5'h0; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_c_T_184 = _instType_c_T_60 ? 5'ha : _instType_c_T_183; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_c_T_185 = _instType_c_T_58 ? 5'h0 : _instType_c_T_184; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_c_T_186 = _instType_c_T_56 ? 5'h0 : _instType_c_T_185; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_c_T_187 = _instType_c_T_54 ? 5'h0 : _instType_c_T_186; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_c_T_188 = _instType_c_T_52 ? 5'h0 : _instType_c_T_187; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_c_T_189 = _instType_c_T_50 ? 5'h7 : _instType_c_T_188; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_c_T_190 = _instType_c_T_48 ? 5'h6 : _instType_c_T_189; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_c_T_191 = _instType_c_T_46 ? 5'h0 : _instType_c_T_190; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_c_T_192 = _instType_c_T_44 ? 5'h0 : _instType_c_T_191; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_c_T_193 = _instType_c_T_42 ? 5'h0 : _instType_c_T_192; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_c_T_194 = _instType_c_T_40 ? 5'h0 : _instType_c_T_193; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_c_T_195 = _instType_c_T_38 ? 5'h0 : _instType_c_T_194; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_c_T_196 = _instType_c_T_36 ? 5'h0 : _instType_c_T_195; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_c_T_197 = _instType_c_T_34 ? 5'h0 : _instType_c_T_196; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_c_T_198 = _instType_c_T_32 ? 5'h0 : _instType_c_T_197; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_c_T_199 = _instType_c_T_30 ? 5'h0 : _instType_c_T_198; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_c_T_200 = _instType_c_T_28 ? 5'h0 : _instType_c_T_199; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_c_T_201 = _instType_c_T_26 ? 5'h0 : _instType_c_T_200; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_c_T_202 = _instType_c_T_24 ? 5'h0 : _instType_c_T_201; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_c_T_203 = _instType_c_T_22 ? 5'h0 : _instType_c_T_202; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_c_T_204 = _instType_c_T_20 ? 5'h0 : _instType_c_T_203; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_c_T_205 = _instType_c_T_18 ? 5'h0 : _instType_c_T_204; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_c_T_206 = _instType_c_T_16 ? 5'h0 : _instType_c_T_205; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_c_T_207 = _instType_c_T_14 ? 5'h0 : _instType_c_T_206; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_c_T_208 = _instType_c_T_12 ? 5'h0 : _instType_c_T_207; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_c_T_209 = _instType_c_T_10 ? 5'hb : _instType_c_T_208; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_c_T_210 = _instType_c_T_8 ? 5'ha : _instType_c_T_209; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_c_T_211 = _instType_c_T_6 ? 5'h7 : _instType_c_T_210; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [4:0] _instType_c_T_212 = _instType_c_T_4 ? 5'h6 : _instType_c_T_211; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_c_T_218 = _instType_c_T_52 ? 1'h0 : _instType_c_T_54 | (_instType_c_T_56 | _instType_c_T_58); // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_c_T_222 = _instType_c_T_44 ? 1'h0 : _instType_c_T_46 | (_instType_c_T_48 | (_instType_c_T_50 |
    _instType_c_T_218)); // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_c_T_223 = _instType_c_T_42 ? 1'h0 : _instType_c_T_222; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_c_T_224 = _instType_c_T_40 ? 1'h0 : _instType_c_T_223; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_c_T_239 = _instType_c_T_10 ? 1'h0 : _instType_c_T_12 | (_instType_c_T_14 | (_instType_c_T_16 | (
    _instType_c_T_18 | (_instType_c_T_20 | (_instType_c_T_22 | (_instType_c_T_24 | (_instType_c_T_26 | (_instType_c_T_28
     | (_instType_c_T_30 | (_instType_c_T_32 | (_instType_c_T_34 | (_instType_c_T_36 | (_instType_c_T_38 |
    _instType_c_T_224))))))))))))); // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _instType_c_T_240 = _instType_c_T_8 ? 1'h0 : _instType_c_T_239; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  instType_c_5 = _instType_c_T_2 | (_instType_c_T_4 | (_instType_c_T_6 | _instType_c_T_240)); // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  is_compress = io_if2id_inst[1:0] != 2'h3; // @[playground/src/noop/decode.scala 56:36]
  wire [11:0] _imm_T_1 = io_if2id_inst[31:20]; // @[playground/src/noop/decode.scala 59:42]
  wire [11:0] _imm_T_5 = {io_if2id_inst[31:25],io_if2id_inst[11:7]}; // @[playground/src/noop/decode.scala 60:64]
  wire [12:0] _imm_T_11 = {io_if2id_inst[31],io_if2id_inst[7],io_if2id_inst[30:25],io_if2id_inst[11:8],1'h0}; // @[playground/src/noop/decode.scala 61:99]
  wire [31:0] _imm_T_14 = {io_if2id_inst[31:12],12'h0}; // @[playground/src/noop/decode.scala 62:59]
  wire [20:0] _imm_T_20 = {io_if2id_inst[31],io_if2id_inst[19:12],io_if2id_inst[20],io_if2id_inst[30:21],1'h0}; // @[playground/src/noop/decode.scala 63:101]
  wire [20:0] _GEN_0 = 3'h6 == instType_0 ? $signed(_imm_T_20) : $signed(21'sh0); // @[playground/src/noop/decode.scala 58:18 63:24 57:9]
  wire [31:0] _GEN_1 = 3'h5 == instType_0 ? $signed(_imm_T_14) : $signed({{11{_GEN_0[20]}},_GEN_0}); // @[playground/src/noop/decode.scala 58:18 62:24]
  wire [31:0] _GEN_2 = 3'h4 == instType_0 ? $signed({{19{_imm_T_11[12]}},_imm_T_11}) : $signed(_GEN_1); // @[playground/src/noop/decode.scala 58:18 61:24]
  wire [31:0] _GEN_3 = 3'h3 == instType_0 ? $signed({{20{_imm_T_5[11]}},_imm_T_5}) : $signed(_GEN_2); // @[playground/src/noop/decode.scala 58:18 60:24]
  wire [31:0] _GEN_4 = 3'h2 == instType_0 ? $signed({{20{_imm_T_1[11]}},_imm_T_1}) : $signed(_GEN_3); // @[playground/src/noop/decode.scala 58:18 59:24]
  wire  _T_7 = ~io_if2id_excep_en; // @[playground/src/noop/decode.scala 65:35]
  wire [11:0] _rs2_r_T_2 = instType_6 ? io_if2id_inst[31:20] : {{7'd0}, io_if2id_inst[24:20]}; // @[playground/src/noop/decode.scala 76:31]
  wire  _indi_r_T_4 = _instType_T_139 | _instType_T_161; // @[playground/src/noop/decode.scala 81:55]
  wire  _indi_r_T_9 = _instType_T_137 | _instType_T_159; // @[playground/src/noop/decode.scala 82:56]
  wire [1:0] _indi_r_T_10 = {_indi_r_T_4,_indi_r_T_9}; // @[playground/src/noop/decode.scala 81:31]
  wire  _T_11 = instType_0 == 3'h7 & _T_7; // @[playground/src/noop/decode.scala 85:32]
  wire  _GEN_5 = instType_0 == 3'h7 & _T_7 | io_if2id_excep_en; // @[playground/src/noop/decode.scala 68:25 85:54 86:29]
  wire [63:0] _GEN_6 = instType_0 == 3'h7 & _T_7 ? 64'h2 : io_if2id_excep_cause; // @[playground/src/noop/decode.scala 68:25 85:54 87:29]
  wire [63:0] _GEN_7 = instType_0 == 3'h7 & _T_7 ? {{32'd0}, io_if2id_inst} : io_if2id_excep_tval; // @[playground/src/noop/decode.scala 68:25 85:54 88:29]
  wire [63:0] _GEN_8 = instType_0 == 3'h7 & _T_7 ? io_if2id_pc : io_if2id_excep_pc; // @[playground/src/noop/decode.scala 68:25 85:54 89:29]
  wire  _GEN_11 = instType_0 == 3'h7 & _T_7 | io_if2id_recov; // @[playground/src/noop/decode.scala 85:54 43:57 84:25]
  wire  _T_12 = instType_0 == 3'h1; // @[playground/src/noop/decode.scala 93:20]
  wire [5:0] _GEN_13 = instType_0 == 3'h1 ? 6'h1a : 6'h1b; // @[playground/src/noop/decode.scala 93:30 96:21 83:25]
  wire [63:0] _rs2_d_r_T_1 = io_if2id_pc + 64'h4; // @[playground/src/noop/decode.scala 102:44]
  wire [63:0] imm = {{32{_GEN_4[31]}},_GEN_4}; // @[playground/src/noop/decode.scala 55:19]
  wire [63:0] _dst_d_r_T = {{32{_GEN_4[31]}},_GEN_4}; // @[playground/src/noop/decode.scala 103:36]
  wire [63:0] _GEN_14 = instType_6 ? {{59'd0}, io_if2id_inst[19:15]} : rs1_d_r; // @[playground/src/noop/decode.scala 104:35 105:29 29:30]
  wire  _GEN_15 = instType_6 ? ~instType_8 : 1'h1; // @[playground/src/noop/decode.scala 104:35 106:29 110:29]
  wire  _GEN_16 = instType_6 | _T_12; // @[playground/src/noop/decode.scala 104:35 107:29]
  wire  _GEN_17 = instType_6 | _T_11; // @[playground/src/noop/decode.scala 104:35 43:17]
  wire  _GEN_18 = instType_6 | _GEN_11; // @[playground/src/noop/decode.scala 104:35 43:57]
  wire [63:0] _GEN_19 = instType_6 ? rs2_d_r : _dst_d_r_T; // @[playground/src/noop/decode.scala 104:35 111:29 32:30]
  wire [1:0] _GEN_20 = instType_5 ? 2'h1 : 2'h0; // @[playground/src/noop/decode.scala 99:27 100:29 79:25]
  wire  _GEN_21 = instType_5 | _GEN_15; // @[playground/src/noop/decode.scala 99:27 101:29]
  wire [63:0] _GEN_22 = instType_5 ? _rs2_d_r_T_1 : _GEN_19; // @[playground/src/noop/decode.scala 99:27 102:29]
  wire [63:0] _GEN_23 = instType_5 ? _dst_d_r_T : dst_d_r; // @[playground/src/noop/decode.scala 99:27 103:29 34:30]
  wire [63:0] _GEN_24 = instType_5 ? rs1_d_r : _GEN_14; // @[playground/src/noop/decode.scala 99:27 29:30]
  wire  _GEN_25 = instType_5 ? _T_12 : _GEN_16; // @[playground/src/noop/decode.scala 99:27]
  wire  _GEN_26 = instType_5 ? _T_11 : _GEN_17; // @[playground/src/noop/decode.scala 99:27]
  wire  _GEN_27 = instType_5 ? _GEN_11 : _GEN_18; // @[playground/src/noop/decode.scala 99:27]
  wire [1:0] _GEN_28 = instType_0 == 3'h2 ? _GEN_20 : 2'h0; // @[playground/src/noop/decode.scala 79:25 98:30]
  wire  _GEN_29 = instType_0 == 3'h2 ? _GEN_21 : _T_12; // @[playground/src/noop/decode.scala 98:30]
  wire [63:0] _GEN_30 = instType_0 == 3'h2 ? _GEN_22 : rs2_d_r; // @[playground/src/noop/decode.scala 32:30 98:30]
  wire [63:0] _GEN_31 = instType_0 == 3'h2 ? _GEN_23 : dst_d_r; // @[playground/src/noop/decode.scala 34:30 98:30]
  wire [63:0] _GEN_32 = instType_0 == 3'h2 ? _GEN_24 : rs1_d_r; // @[playground/src/noop/decode.scala 29:30 98:30]
  wire  _GEN_33 = instType_0 == 3'h2 ? _GEN_25 : _T_12; // @[playground/src/noop/decode.scala 98:30]
  wire  _GEN_34 = instType_0 == 3'h2 ? _GEN_26 : _T_11; // @[playground/src/noop/decode.scala 98:30]
  wire  _GEN_35 = instType_0 == 3'h2 ? _GEN_27 : _GEN_11; // @[playground/src/noop/decode.scala 98:30]
  wire  _GEN_36 = instType_0 == 3'h3 | _GEN_29; // @[playground/src/noop/decode.scala 114:30 115:25]
  wire  _GEN_37 = instType_0 == 3'h3 | _GEN_33; // @[playground/src/noop/decode.scala 114:30 116:25]
  wire [5:0] _GEN_38 = instType_0 == 3'h3 ? 6'h1e : _GEN_13; // @[playground/src/noop/decode.scala 114:30 117:25]
  wire [63:0] _GEN_39 = instType_0 == 3'h3 ? _dst_d_r_T : _GEN_31; // @[playground/src/noop/decode.scala 114:30 118:25]
  wire [63:0] _dst_d_r_T_6 = $signed(io_if2id_pc) + $signed(imm); // @[playground/src/noop/decode.scala 123:61]
  wire  _GEN_40 = instType_0 == 3'h4 | _GEN_36; // @[playground/src/noop/decode.scala 120:30 121:25]
  wire  _GEN_41 = instType_0 == 3'h4 | _GEN_37; // @[playground/src/noop/decode.scala 120:30 122:25]
  wire [63:0] _GEN_42 = instType_0 == 3'h4 ? _dst_d_r_T_6 : _GEN_39; // @[playground/src/noop/decode.scala 120:30 123:25]
  wire [2:0] _GEN_43 = instType_0 == 3'h4 ? io_if2id_inst[14:12] : ctrl_r_brType; // @[playground/src/noop/decode.scala 120:30 124:27 26:30]
  wire [1:0] _GEN_44 = instType_0 == 3'h4 ? 2'h2 : _GEN_28; // @[playground/src/noop/decode.scala 120:30 125:25]
  wire [63:0] _GEN_45 = instType_0 == 3'h5 ? _dst_d_r_T : _GEN_32; // @[playground/src/noop/decode.scala 127:30 128:25]
  wire [63:0] _GEN_46 = instType_0 == 3'h5 ? io_if2id_pc : _GEN_30; // @[playground/src/noop/decode.scala 127:30 129:25]
  wire [63:0] _GEN_47 = instType_0 == 3'h6 ? _dst_d_r_T_6 : _GEN_45; // @[playground/src/noop/decode.scala 131:30 132:25]
  wire [63:0] _GEN_48 = instType_0 == 3'h6 ? _rs2_d_r_T_1 : _GEN_46; // @[playground/src/noop/decode.scala 131:30 133:25]
  wire [63:0] _GEN_49 = instType_0 == 3'h6 ? 64'h0 : _GEN_42; // @[playground/src/noop/decode.scala 131:30 134:25]
  wire [1:0] _GEN_50 = instType_0 == 3'h6 ? 2'h1 : _GEN_44; // @[playground/src/noop/decode.scala 131:30 135:24]
  wire  _excep_r_cause_T = io_idState_priv == 2'h3; // @[playground/src/noop/decode.scala 141:34]
  wire  _excep_r_cause_T_1 = io_idState_priv == 2'h1; // @[playground/src/noop/decode.scala 142:34]
  wire [3:0] _excep_r_cause_T_2 = _excep_r_cause_T_1 ? 4'h9 : 4'h8; // @[src/main/scala/chisel3/util/Mux.scala 47:70]
  wire [3:0] _excep_r_cause_T_3 = _excep_r_cause_T ? 4'hb : _excep_r_cause_T_2; // @[src/main/scala/chisel3/util/Mux.scala 47:70]
  wire [9:0] _rs2_r_T_4 = _excep_r_cause_T ? 10'h305 : 10'h105; // @[playground/src/noop/decode.scala 146:32]
  wire [63:0] _GEN_51 = 32'h73 == io_if2id_inst ? io_if2id_pc : _GEN_8; // @[playground/src/noop/decode.scala 137:38 138:25]
  wire  _GEN_52 = 32'h73 == io_if2id_inst | _GEN_5; // @[playground/src/noop/decode.scala 137:38 139:25]
  wire [63:0] _GEN_53 = 32'h73 == io_if2id_inst ? {{60'd0}, _excep_r_cause_T_3} : _GEN_6; // @[playground/src/noop/decode.scala 137:38 140:27]
  wire [63:0] _GEN_54 = 32'h73 == io_if2id_inst ? 64'h0 : _GEN_7; // @[playground/src/noop/decode.scala 137:38 144:27]
  wire [1:0] _GEN_55 = 32'h73 == io_if2id_inst ? 2'h3 : _GEN_50; // @[playground/src/noop/decode.scala 137:38 145:25]
  wire [11:0] _GEN_56 = 32'h73 == io_if2id_inst ? {{2'd0}, _rs2_r_T_4} : _rs2_r_T_2; // @[playground/src/noop/decode.scala 137:38 146:25 76:25]
  wire  _GEN_57 = 32'h73 == io_if2id_inst | _GEN_34; // @[playground/src/noop/decode.scala 137:38 43:17]
  wire  _GEN_58 = 32'h73 == io_if2id_inst | _GEN_35; // @[playground/src/noop/decode.scala 137:38 43:57]
  wire [63:0] _GEN_59 = 32'h10200073 == io_if2id_inst ? io_if2id_pc : _GEN_51; // @[playground/src/noop/decode.scala 149:37 150:25]
  wire  _GEN_60 = 32'h10200073 == io_if2id_inst | _GEN_52; // @[playground/src/noop/decode.scala 149:37 151:25]
  wire [1:0] _GEN_61 = 32'h10200073 == io_if2id_inst ? 2'h2 : 2'h0; // @[playground/src/noop/decode.scala 149:37 152:27]
  wire [63:0] _GEN_62 = 32'h10200073 == io_if2id_inst ? 64'h0 : _GEN_53; // @[playground/src/noop/decode.scala 149:37 153:27]
  wire [63:0] _GEN_63 = 32'h10200073 == io_if2id_inst ? 64'h0 : _GEN_54; // @[playground/src/noop/decode.scala 149:37 154:27]
  wire [1:0] _GEN_64 = 32'h10200073 == io_if2id_inst ? 2'h3 : _GEN_55; // @[playground/src/noop/decode.scala 149:37 155:25]
  wire [11:0] _GEN_65 = 32'h10200073 == io_if2id_inst ? 12'h141 : _GEN_56; // @[playground/src/noop/decode.scala 149:37 156:25]
  wire  _GEN_66 = 32'h10200073 == io_if2id_inst | _GEN_57; // @[playground/src/noop/decode.scala 149:37 43:17]
  wire  _GEN_67 = 32'h10200073 == io_if2id_inst | _GEN_58; // @[playground/src/noop/decode.scala 149:37 43:57]
  wire [63:0] _GEN_68 = 32'h30200073 == io_if2id_inst ? io_if2id_pc : _GEN_59; // @[playground/src/noop/decode.scala 159:37 160:25]
  wire  _GEN_69 = 32'h30200073 == io_if2id_inst | _GEN_60; // @[playground/src/noop/decode.scala 159:37 161:25]
  wire [1:0] _GEN_70 = 32'h30200073 == io_if2id_inst ? 2'h3 : _GEN_61; // @[playground/src/noop/decode.scala 159:37 162:27]
  wire [63:0] _GEN_71 = 32'h30200073 == io_if2id_inst ? 64'h0 : _GEN_62; // @[playground/src/noop/decode.scala 159:37 163:27]
  wire [63:0] _GEN_72 = 32'h30200073 == io_if2id_inst ? 64'h0 : _GEN_63; // @[playground/src/noop/decode.scala 159:37 164:27]
  wire [1:0] _GEN_73 = 32'h30200073 == io_if2id_inst ? 2'h3 : _GEN_64; // @[playground/src/noop/decode.scala 159:37 165:25]
  wire  _GEN_75 = 32'h30200073 == io_if2id_inst | _GEN_66; // @[playground/src/noop/decode.scala 159:37 43:17]
  wire  _GEN_76 = 32'h30200073 == io_if2id_inst | _GEN_67; // @[playground/src/noop/decode.scala 159:37 43:57]
  wire [1:0] _GEN_77 = _instType_T_183 ? 2'h1 : 2'h0; // @[playground/src/noop/decode.scala 169:40 170:23 80:25]
  wire  _GEN_78 = _instType_T_183 | _GEN_75; // @[playground/src/noop/decode.scala 169:40 43:17]
  wire  _GEN_79 = _instType_T_183 | _GEN_76; // @[playground/src/noop/decode.scala 169:40 43:57]
  wire [1:0] _GEN_80 = _instType_T_185 ? 2'h2 : _GEN_77; // @[playground/src/noop/decode.scala 173:43 174:23]
  wire  _GEN_81 = _instType_T_185 | _GEN_78; // @[playground/src/noop/decode.scala 173:43 43:17]
  wire  _GEN_82 = _instType_T_185 | _GEN_79; // @[playground/src/noop/decode.scala 173:43 43:57]
  wire  _GEN_105 = hs_in & ~is_compress & ~io_if2id_excep_en & _GEN_81; // @[playground/src/noop/decode.scala 19:33 65:54]
  wire [63:0] _GEN_106 = hs_in & ~is_compress & ~io_if2id_excep_en ? _GEN_48 : rs2_d_r; // @[playground/src/noop/decode.scala 32:30 65:54]
  wire [63:0] _GEN_107 = hs_in & ~is_compress & ~io_if2id_excep_en ? _GEN_49 : dst_d_r; // @[playground/src/noop/decode.scala 34:30 65:54]
  wire [63:0] _GEN_108 = hs_in & ~is_compress & ~io_if2id_excep_en ? _GEN_47 : rs1_d_r; // @[playground/src/noop/decode.scala 29:30 65:54]
  wire [2:0] _GEN_109 = hs_in & ~is_compress & ~io_if2id_excep_en ? _GEN_43 : ctrl_r_brType; // @[playground/src/noop/decode.scala 26:30 65:54]
  wire [63:0] _imm_c_T_5 = {54'h0,io_if2id_inst[10:7],io_if2id_inst[12:11],io_if2id_inst[5],io_if2id_inst[6],2'h0}; // @[playground/src/noop/decode.scala 185:106]
  wire [63:0] _imm_c_T_10 = {57'h0,io_if2id_inst[5],io_if2id_inst[12:10],io_if2id_inst[6],2'h0}; // @[playground/src/noop/decode.scala 186:92]
  wire [63:0] _imm_c_T_14 = {56'h0,io_if2id_inst[6:5],io_if2id_inst[12:10],3'h0}; // @[playground/src/noop/decode.scala 187:83]
  wire [63:0] _imm_c_T_18 = {58'h0,io_if2id_inst[12],io_if2id_inst[6:2]}; // @[playground/src/noop/decode.scala 188:70]
  wire [5:0] _imm_c_T_22 = {io_if2id_inst[12],io_if2id_inst[6:2]}; // @[playground/src/noop/decode.scala 189:59]
  wire [63:0] _imm_c_T_27 = {56'h0,io_if2id_inst[3:2],io_if2id_inst[12],io_if2id_inst[6:4],2'h0}; // @[playground/src/noop/decode.scala 190:93]
  wire [63:0] _imm_c_T_32 = {55'h0,io_if2id_inst[4:2],io_if2id_inst[12],io_if2id_inst[6:5],3'h0}; // @[playground/src/noop/decode.scala 191:93]
  wire [9:0] _imm_c_T_39 = {io_if2id_inst[12],io_if2id_inst[4:3],io_if2id_inst[5],io_if2id_inst[2],io_if2id_inst[6],4'h0
    }; // @[playground/src/noop/decode.scala 192:102]
  wire [17:0] _imm_c_T_43 = {io_if2id_inst[12],io_if2id_inst[6:2],12'h0}; // @[playground/src/noop/decode.scala 193:70]
  wire [11:0] _imm_c_T_53 = {io_if2id_inst[12],io_if2id_inst[8],io_if2id_inst[10:9],io_if2id_inst[6],io_if2id_inst[7],
    io_if2id_inst[2],io_if2id_inst[11],io_if2id_inst[5:3],1'h0}; // @[playground/src/noop/decode.scala 194:139]
  wire [8:0] _imm_c_T_60 = {io_if2id_inst[12],io_if2id_inst[6:5],io_if2id_inst[2],io_if2id_inst[11:10],io_if2id_inst[4:3
    ],1'h0}; // @[playground/src/noop/decode.scala 195:108]
  wire [63:0] _imm_c_T_64 = {56'h0,io_if2id_inst[8:7],io_if2id_inst[12:9],2'h0}; // @[playground/src/noop/decode.scala 196:82]
  wire [63:0] _imm_c_T_68 = {55'h0,io_if2id_inst[9:7],io_if2id_inst[12:10],3'h0}; // @[playground/src/noop/decode.scala 197:83]
  wire [63:0] _GEN_110 = 4'hd == instType_c_1 ? $signed(_imm_c_T_68) : $signed(64'sh0); // @[playground/src/noop/decode.scala 182:11 184:20 197:27]
  wire [63:0] _GEN_111 = 4'hc == instType_c_1 ? $signed(_imm_c_T_64) : $signed(_GEN_110); // @[playground/src/noop/decode.scala 184:20 196:27]
  wire [63:0] _GEN_112 = 4'hb == instType_c_1 ? $signed({{55{_imm_c_T_60[8]}},_imm_c_T_60}) : $signed(_GEN_111); // @[playground/src/noop/decode.scala 184:20 195:27]
  wire [63:0] _GEN_113 = 4'ha == instType_c_1 ? $signed({{52{_imm_c_T_53[11]}},_imm_c_T_53}) : $signed(_GEN_112); // @[playground/src/noop/decode.scala 184:20 194:27]
  wire [63:0] _GEN_114 = 4'h9 == instType_c_1 ? $signed({{46{_imm_c_T_43[17]}},_imm_c_T_43}) : $signed(_GEN_113); // @[playground/src/noop/decode.scala 184:20 193:27]
  wire [63:0] _GEN_115 = 4'h8 == instType_c_1 ? $signed({{54{_imm_c_T_39[9]}},_imm_c_T_39}) : $signed(_GEN_114); // @[playground/src/noop/decode.scala 184:20 192:27]
  wire [63:0] _GEN_116 = 4'h7 == instType_c_1 ? $signed(_imm_c_T_32) : $signed(_GEN_115); // @[playground/src/noop/decode.scala 184:20 191:27]
  wire [63:0] _GEN_117 = 4'h6 == instType_c_1 ? $signed(_imm_c_T_27) : $signed(_GEN_116); // @[playground/src/noop/decode.scala 184:20 190:27]
  wire [63:0] _GEN_118 = 4'h5 == instType_c_1 ? $signed({{58{_imm_c_T_22[5]}},_imm_c_T_22}) : $signed(_GEN_117); // @[playground/src/noop/decode.scala 184:20 189:27]
  wire [63:0] _GEN_119 = 4'h4 == instType_c_1 ? $signed(_imm_c_T_18) : $signed(_GEN_118); // @[playground/src/noop/decode.scala 184:20 188:27]
  wire [63:0] _GEN_120 = 4'h3 == instType_c_1 ? $signed(_imm_c_T_14) : $signed(_GEN_119); // @[playground/src/noop/decode.scala 184:20 187:27]
  wire [63:0] _GEN_121 = 4'h2 == instType_c_1 ? $signed(_imm_c_T_10) : $signed(_GEN_120); // @[playground/src/noop/decode.scala 184:20 186:27]
  wire [63:0] imm_c = 4'h1 == instType_c_1 ? $signed(_imm_c_T_5) : $signed(_GEN_121); // @[playground/src/noop/decode.scala 184:20 185:27]
  wire [30:0] _inst_r_T = {15'h0,io_if2id_inst[15:0]}; // @[playground/src/noop/decode.scala 200:23]
  wire  _GEN_123 = instType_c_0 == 4'h0 & _T_7 | io_if2id_excep_en; // @[playground/src/noop/decode.scala 202:25 218:58 219:29]
  wire  _GEN_128 = instType_c_0 == 4'h0 & _T_7 | _GEN_105; // @[playground/src/noop/decode.scala 218:58 43:17]
  wire  _GEN_129 = instType_c_0 == 4'h0 & _T_7 | io_if2id_recov; // @[playground/src/noop/decode.scala 217:25 218:58 43:57]
  wire  _T_47 = instType_c_0 == 4'h1; // @[playground/src/noop/decode.scala 226:22]
  wire [1:0] _GEN_130 = _instType_c_T_52 ? 2'h1 : 2'h0; // @[playground/src/noop/decode.scala 213:25 229:34 230:29]
  wire [63:0] _GEN_131 = _instType_c_T_52 ? 64'h0 : _GEN_107; // @[playground/src/noop/decode.scala 229:34 231:29]
  wire [63:0] _rs2_d_r_T_6 = io_if2id_pc + 64'h2; // @[playground/src/noop/decode.scala 236:44]
  wire [1:0] _GEN_132 = _instType_c_T_56 ? 2'h1 : _GEN_130; // @[playground/src/noop/decode.scala 233:36 234:29]
  wire  _GEN_133 = _instType_c_T_56 ? 1'h0 : 1'h1; // @[playground/src/noop/decode.scala 228:20 233:36 235:29]
  wire [63:0] _GEN_134 = _instType_c_T_56 ? _rs2_d_r_T_6 : _GEN_106; // @[playground/src/noop/decode.scala 233:36 236:29]
  wire [63:0] _GEN_135 = _instType_c_T_56 ? 64'h0 : _GEN_131; // @[playground/src/noop/decode.scala 233:36 237:29]
  wire [4:0] _GEN_136 = _instType_c_T_56 ? 5'h1 : io_if2id_inst[11:7]; // @[playground/src/noop/decode.scala 212:25 233:36 238:29]
  wire  _GEN_138 = instType_c_0 == 4'h1 & _GEN_133; // @[playground/src/noop/decode.scala 211:25 226:29]
  wire [1:0] _GEN_139 = instType_c_0 == 4'h1 ? _GEN_132 : 2'h0; // @[playground/src/noop/decode.scala 213:25 226:29]
  wire [63:0] _GEN_140 = instType_c_0 == 4'h1 ? _GEN_135 : _GEN_107; // @[playground/src/noop/decode.scala 226:29]
  wire [63:0] _GEN_141 = instType_c_0 == 4'h1 ? _GEN_134 : _GEN_106; // @[playground/src/noop/decode.scala 226:29]
  wire [4:0] _GEN_142 = instType_c_0 == 4'h1 ? _GEN_136 : io_if2id_inst[11:7]; // @[playground/src/noop/decode.scala 212:25 226:29]
  wire [63:0] _rs2_d_r_T_7 = 4'h1 == instType_c_1 ? $signed(_imm_c_T_5) : $signed(_GEN_121); // @[playground/src/noop/decode.scala 243:30]
  wire [4:0] _GEN_143 = _instType_c_T_48 | _instType_c_T_50 ? 5'h2 : io_if2id_inst[11:7]; // @[playground/src/noop/decode.scala 244:57 245:23 208:25]
  wire  _GEN_144 = instType_c_0 == 4'h2 | _T_47; // @[playground/src/noop/decode.scala 241:29 242:21]
  wire [63:0] _GEN_145 = instType_c_0 == 4'h2 ? _rs2_d_r_T_7 : _GEN_141; // @[playground/src/noop/decode.scala 241:29 243:21]
  wire [4:0] _GEN_146 = instType_c_0 == 4'h2 ? _GEN_143 : io_if2id_inst[11:7]; // @[playground/src/noop/decode.scala 208:25 241:29]
  wire  _GEN_147 = instType_c_0 == 4'h3 | _GEN_144; // @[playground/src/noop/decode.scala 248:30 249:21]
  wire [4:0] _GEN_148 = instType_c_0 == 4'h3 ? 5'h2 : _GEN_146; // @[playground/src/noop/decode.scala 248:30 250:21]
  wire  _GEN_149 = instType_c_0 == 4'h3 | _GEN_138; // @[playground/src/noop/decode.scala 248:30 251:21]
  wire [4:0] _GEN_150 = instType_c_0 == 4'h3 ? io_if2id_inst[6:2] : io_if2id_inst[6:2]; // @[playground/src/noop/decode.scala 248:30 252:21 210:25]
  wire [63:0] _GEN_151 = instType_c_0 == 4'h3 ? _rs2_d_r_T_7 : _GEN_140; // @[playground/src/noop/decode.scala 248:30 253:21]
  wire [5:0] _GEN_152 = instType_c_0 == 4'h3 ? 6'h1e : 6'h1b; // @[playground/src/noop/decode.scala 248:30 254:21 216:25]
  wire [3:0] _dst_r_T_4 = {1'h1,io_if2id_inst[4:2]}; // @[playground/src/noop/common.scala 675:12]
  wire  _GEN_153 = instType_c_0 == 4'h4 | _GEN_147; // @[playground/src/noop/decode.scala 256:30 257:21]
  wire [4:0] _GEN_154 = instType_c_0 == 4'h4 ? 5'h2 : _GEN_148; // @[playground/src/noop/decode.scala 256:30 258:21]
  wire [63:0] _GEN_155 = instType_c_0 == 4'h4 ? _rs2_d_r_T_7 : _GEN_145; // @[playground/src/noop/decode.scala 256:30 259:21]
  wire [4:0] _GEN_156 = instType_c_0 == 4'h4 ? {{1'd0}, _dst_r_T_4} : _GEN_142; // @[playground/src/noop/decode.scala 256:30 260:21]
  wire [3:0] _rs1_r_T_4 = {1'h1,io_if2id_inst[9:7]}; // @[playground/src/noop/common.scala 675:12]
  wire  _GEN_157 = instType_c_0 == 4'h5 | _GEN_153; // @[playground/src/noop/decode.scala 262:29 263:21]
  wire [4:0] _GEN_158 = instType_c_0 == 4'h5 ? {{1'd0}, _rs1_r_T_4} : _GEN_154; // @[playground/src/noop/decode.scala 262:29 264:21]
  wire [4:0] _GEN_160 = instType_c_0 == 4'h5 ? {{1'd0}, _dst_r_T_4} : _GEN_156; // @[playground/src/noop/decode.scala 262:29 266:21]
  wire [5:0] _GEN_161 = io_if2id_inst[1:0] == 2'h0 ? 6'h1e : _GEN_152; // @[playground/src/noop/decode.scala 275:38 276:25]
  wire  _GEN_162 = instType_c_0 == 4'h6 | _GEN_157; // @[playground/src/noop/decode.scala 268:29 269:21]
  wire  _GEN_164 = instType_c_0 == 4'h6 | _GEN_149; // @[playground/src/noop/decode.scala 268:29 271:21]
  wire [4:0] _GEN_165 = instType_c_0 == 4'h6 ? {{1'd0}, _dst_r_T_4} : _GEN_150; // @[playground/src/noop/decode.scala 268:29 272:21]
  wire [63:0] _GEN_166 = instType_c_0 == 4'h6 ? _rs2_d_r_T_7 : _GEN_151; // @[playground/src/noop/decode.scala 268:29 273:21]
  wire [63:0] _dst_d_r_T_13 = $signed(io_if2id_pc) + $signed(imm_c); // @[playground/src/noop/decode.scala 283:53]
  wire [2:0] _GEN_169 = _instType_c_T_42 ? 3'h0 : _GEN_109; // @[playground/src/noop/decode.scala 285:36 286:31]
  wire [63:0] _GEN_170 = _instType_c_T_42 ? 64'h0 : _rs2_d_r_T_7; // @[playground/src/noop/decode.scala 282:21 285:36 287:29]
  wire [1:0] _GEN_171 = _instType_c_T_42 ? 2'h2 : _GEN_139; // @[playground/src/noop/decode.scala 285:36 288:29]
  wire [2:0] _GEN_172 = _instType_c_T_44 ? 3'h1 : _GEN_169; // @[playground/src/noop/decode.scala 290:36 291:31]
  wire [1:0] _GEN_174 = _instType_c_T_44 ? 2'h2 : _GEN_171; // @[playground/src/noop/decode.scala 290:36 293:29]
  wire  _GEN_175 = instType_c_0 == 4'h7 | _GEN_162; // @[playground/src/noop/decode.scala 279:29 280:21]
  wire [1:0] _GEN_181 = instType_c_0 == 4'h7 ? _GEN_174 : _GEN_139; // @[playground/src/noop/decode.scala 279:29]
  wire  _GEN_233 = valid_r & ~hs_out ? 1'h0 : io_if2id_valid; // @[playground/src/noop/decode.scala 316:20 318:33]
  wire  _GEN_235 = hs_out ? 1'h0 : valid_r; // @[playground/src/noop/decode.scala 326:26 327:20 40:30]
  wire  _GEN_236 = hs_in | _GEN_235; // @[playground/src/noop/decode.scala 324:19 325:20]
  wire  _GEN_237 = _io_if2id_stall_T & _GEN_236; // @[playground/src/noop/decode.scala 323:25 331:17]
  assign io_if2id_drop = drop_r | io_id2df_drop; // @[playground/src/noop/decode.scala 20:30]
  assign io_if2id_stall = stall_r & ~io_id2df_drop | io_id2df_stall; // @[playground/src/noop/decode.scala 22:52]
  assign io_if2id_ready = ~drop_in & _GEN_233; // @[playground/src/noop/decode.scala 317:19 316:20]
  assign io_id2df_inst = inst_r; // @[playground/src/noop/decode.scala 333:25]
  assign io_id2df_pc = pc_r; // @[playground/src/noop/decode.scala 334:25]
  assign io_id2df_excep_cause = excep_r_cause; // @[playground/src/noop/decode.scala 335:25]
  assign io_id2df_excep_tval = excep_r_tval; // @[playground/src/noop/decode.scala 335:25]
  assign io_id2df_excep_en = excep_r_en; // @[playground/src/noop/decode.scala 335:25]
  assign io_id2df_excep_pc = excep_r_pc; // @[playground/src/noop/decode.scala 335:25]
  assign io_id2df_excep_etype = excep_r_etype; // @[playground/src/noop/decode.scala 335:25]
  assign io_id2df_ctrl_aluOp = ctrl_r_aluOp; // @[playground/src/noop/decode.scala 336:25]
  assign io_id2df_ctrl_aluWidth = ctrl_r_aluWidth; // @[playground/src/noop/decode.scala 336:25]
  assign io_id2df_ctrl_dcMode = ctrl_r_dcMode; // @[playground/src/noop/decode.scala 336:25]
  assign io_id2df_ctrl_writeRegEn = ctrl_r_writeRegEn; // @[playground/src/noop/decode.scala 336:25]
  assign io_id2df_ctrl_writeCSREn = ctrl_r_writeCSREn; // @[playground/src/noop/decode.scala 336:25]
  assign io_id2df_ctrl_brType = ctrl_r_brType; // @[playground/src/noop/decode.scala 336:25]
  assign io_id2df_rs1 = rs1_r; // @[playground/src/noop/decode.scala 337:25]
  assign io_id2df_rrs1 = rrs1_r; // @[playground/src/noop/decode.scala 338:25]
  assign io_id2df_rs1_d = rs1_d_r; // @[playground/src/noop/decode.scala 339:25]
  assign io_id2df_rs2 = rs2_r; // @[playground/src/noop/decode.scala 340:25]
  assign io_id2df_rrs2 = rrs2_r; // @[playground/src/noop/decode.scala 341:25]
  assign io_id2df_rs2_d = rs2_d_r; // @[playground/src/noop/decode.scala 342:25]
  assign io_id2df_dst = dst_r; // @[playground/src/noop/decode.scala 343:25]
  assign io_id2df_dst_d = dst_d_r; // @[playground/src/noop/decode.scala 344:25]
  assign io_id2df_jmp_type = jmp_type_r; // @[playground/src/noop/decode.scala 345:25]
  assign io_id2df_special = special_r; // @[playground/src/noop/decode.scala 346:25]
  assign io_id2df_swap = swap_r; // @[playground/src/noop/decode.scala 347:25]
  assign io_id2df_indi = indi_r; // @[playground/src/noop/decode.scala 348:25]
  assign io_id2df_recov = recov_r; // @[playground/src/noop/decode.scala 349:25]
  assign io_id2df_valid = valid_r; // @[playground/src/noop/decode.scala 350:25]
  always @(posedge clock) begin
    if (reset) begin // @[playground/src/noop/decode.scala 17:30]
      drop_r <= 1'h0; // @[playground/src/noop/decode.scala 17:30]
    end else if (hs_in & is_compress & _T_7) begin // @[playground/src/noop/decode.scala 199:53]
      drop_r <= _GEN_128;
    end else begin
      drop_r <= _GEN_105;
    end
    if (reset) begin // @[playground/src/noop/decode.scala 18:30]
      stall_r <= 1'h0; // @[playground/src/noop/decode.scala 18:30]
    end else if (hs_in & is_compress & _T_7) begin // @[playground/src/noop/decode.scala 199:53]
      stall_r <= _GEN_128;
    end else begin
      stall_r <= _GEN_105;
    end
    if (reset) begin // @[playground/src/noop/decode.scala 23:30]
      inst_r <= 32'h0; // @[playground/src/noop/decode.scala 23:30]
    end else if (hs_in & io_if2id_excep_en) begin // @[playground/src/noop/decode.scala 302:37]
      inst_r <= io_if2id_inst; // @[playground/src/noop/decode.scala 303:25]
    end else if (hs_in & is_compress & _T_7) begin // @[playground/src/noop/decode.scala 199:53]
      inst_r <= {{1'd0}, _inst_r_T}; // @[playground/src/noop/decode.scala 200:17]
    end else if (hs_in & ~is_compress & ~io_if2id_excep_en) begin // @[playground/src/noop/decode.scala 65:54]
      inst_r <= io_if2id_inst; // @[playground/src/noop/decode.scala 66:25]
    end
    if (reset) begin // @[playground/src/noop/decode.scala 24:30]
      pc_r <= 64'h0; // @[playground/src/noop/decode.scala 24:30]
    end else if (hs_in & io_if2id_excep_en) begin // @[playground/src/noop/decode.scala 302:37]
      pc_r <= io_if2id_pc; // @[playground/src/noop/decode.scala 304:25]
    end else if (hs_in & is_compress & _T_7) begin // @[playground/src/noop/decode.scala 199:53]
      pc_r <= io_if2id_pc; // @[playground/src/noop/decode.scala 201:17]
    end else if (hs_in & ~is_compress & ~io_if2id_excep_en) begin // @[playground/src/noop/decode.scala 65:54]
      pc_r <= io_if2id_pc; // @[playground/src/noop/decode.scala 67:25]
    end
    if (reset) begin // @[playground/src/noop/decode.scala 25:30]
      excep_r_cause <= 64'h0; // @[playground/src/noop/decode.scala 25:30]
    end else if (hs_in & io_if2id_excep_en) begin // @[playground/src/noop/decode.scala 302:37]
      excep_r_cause <= io_if2id_excep_cause; // @[playground/src/noop/decode.scala 305:25]
    end else if (hs_in & is_compress & _T_7) begin // @[playground/src/noop/decode.scala 199:53]
      if (instType_c_0 == 4'h0 & _T_7) begin // @[playground/src/noop/decode.scala 218:58]
        excep_r_cause <= 64'h2; // @[playground/src/noop/decode.scala 220:29]
      end else begin
        excep_r_cause <= io_if2id_excep_cause; // @[playground/src/noop/decode.scala 202:25]
      end
    end else if (hs_in & ~is_compress & ~io_if2id_excep_en) begin // @[playground/src/noop/decode.scala 65:54]
      excep_r_cause <= _GEN_71;
    end
    if (reset) begin // @[playground/src/noop/decode.scala 25:30]
      excep_r_tval <= 64'h0; // @[playground/src/noop/decode.scala 25:30]
    end else if (hs_in & io_if2id_excep_en) begin // @[playground/src/noop/decode.scala 302:37]
      excep_r_tval <= io_if2id_excep_tval; // @[playground/src/noop/decode.scala 305:25]
    end else if (hs_in & is_compress & _T_7) begin // @[playground/src/noop/decode.scala 199:53]
      if (instType_c_0 == 4'h0 & _T_7) begin // @[playground/src/noop/decode.scala 218:58]
        excep_r_tval <= {{33'd0}, _inst_r_T}; // @[playground/src/noop/decode.scala 221:29]
      end else begin
        excep_r_tval <= io_if2id_excep_tval; // @[playground/src/noop/decode.scala 202:25]
      end
    end else if (hs_in & ~is_compress & ~io_if2id_excep_en) begin // @[playground/src/noop/decode.scala 65:54]
      excep_r_tval <= _GEN_72;
    end
    if (reset) begin // @[playground/src/noop/decode.scala 25:30]
      excep_r_en <= 1'h0; // @[playground/src/noop/decode.scala 25:30]
    end else if (hs_in & io_if2id_excep_en) begin // @[playground/src/noop/decode.scala 302:37]
      excep_r_en <= io_if2id_excep_en; // @[playground/src/noop/decode.scala 305:25]
    end else if (hs_in & is_compress & _T_7) begin // @[playground/src/noop/decode.scala 199:53]
      excep_r_en <= _GEN_123;
    end else if (hs_in & ~is_compress & ~io_if2id_excep_en) begin // @[playground/src/noop/decode.scala 65:54]
      excep_r_en <= _GEN_69;
    end
    if (reset) begin // @[playground/src/noop/decode.scala 25:30]
      excep_r_pc <= 64'h0; // @[playground/src/noop/decode.scala 25:30]
    end else if (hs_in & io_if2id_excep_en) begin // @[playground/src/noop/decode.scala 302:37]
      excep_r_pc <= io_if2id_excep_pc; // @[playground/src/noop/decode.scala 305:25]
    end else if (hs_in & is_compress & _T_7) begin // @[playground/src/noop/decode.scala 199:53]
      if (instType_c_0 == 4'h0 & _T_7) begin // @[playground/src/noop/decode.scala 218:58]
        excep_r_pc <= io_if2id_pc; // @[playground/src/noop/decode.scala 222:29]
      end else begin
        excep_r_pc <= io_if2id_excep_pc; // @[playground/src/noop/decode.scala 202:25]
      end
    end else if (hs_in & ~is_compress & ~io_if2id_excep_en) begin // @[playground/src/noop/decode.scala 65:54]
      excep_r_pc <= _GEN_68;
    end
    if (reset) begin // @[playground/src/noop/decode.scala 25:30]
      excep_r_etype <= 2'h0; // @[playground/src/noop/decode.scala 25:30]
    end else if (hs_in & io_if2id_excep_en) begin // @[playground/src/noop/decode.scala 302:37]
      excep_r_etype <= 2'h0; // @[playground/src/noop/decode.scala 305:25]
    end else if (hs_in & is_compress & _T_7) begin // @[playground/src/noop/decode.scala 199:53]
      excep_r_etype <= 2'h0;
    end else if (hs_in & ~is_compress & ~io_if2id_excep_en) begin // @[playground/src/noop/decode.scala 65:54]
      excep_r_etype <= _GEN_70;
    end
    if (reset) begin // @[playground/src/noop/decode.scala 26:30]
      ctrl_r_aluOp <= 5'h0; // @[playground/src/noop/decode.scala 26:30]
    end else if (hs_in & io_if2id_excep_en) begin // @[playground/src/noop/decode.scala 302:37]
      ctrl_r_aluOp <= 5'h0; // @[playground/src/noop/decode.scala 306:25]
    end else if (hs_in & is_compress & _T_7) begin // @[playground/src/noop/decode.scala 199:53]
      if (_instType_c_T_2) begin // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
        ctrl_r_aluOp <= 5'h3;
      end else begin
        ctrl_r_aluOp <= _instType_c_T_152;
      end
    end else if (hs_in & ~is_compress & ~io_if2id_excep_en) begin // @[playground/src/noop/decode.scala 65:54]
      ctrl_r_aluOp <= instType_1; // @[playground/src/noop/decode.scala 69:27]
    end
    if (reset) begin // @[playground/src/noop/decode.scala 26:30]
      ctrl_r_aluWidth <= 1'h0; // @[playground/src/noop/decode.scala 26:30]
    end else if (hs_in & io_if2id_excep_en) begin // @[playground/src/noop/decode.scala 302:37]
      ctrl_r_aluWidth <= 1'h0; // @[playground/src/noop/decode.scala 306:25]
    end else if (hs_in & is_compress & _T_7) begin // @[playground/src/noop/decode.scala 199:53]
      if (_instType_c_T_2) begin // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
        ctrl_r_aluWidth <= 1'h0;
      end else begin
        ctrl_r_aluWidth <= _instType_c_T_182;
      end
    end else if (hs_in & ~is_compress & ~io_if2id_excep_en) begin // @[playground/src/noop/decode.scala 65:54]
      ctrl_r_aluWidth <= instType_2; // @[playground/src/noop/decode.scala 70:27]
    end
    if (reset) begin // @[playground/src/noop/decode.scala 26:30]
      ctrl_r_dcMode <= 5'h0; // @[playground/src/noop/decode.scala 26:30]
    end else if (hs_in & io_if2id_excep_en) begin // @[playground/src/noop/decode.scala 302:37]
      ctrl_r_dcMode <= 5'h0; // @[playground/src/noop/decode.scala 306:25]
    end else if (hs_in & is_compress & _T_7) begin // @[playground/src/noop/decode.scala 199:53]
      if (_instType_c_T_2) begin // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
        ctrl_r_dcMode <= 5'h0;
      end else begin
        ctrl_r_dcMode <= _instType_c_T_212;
      end
    end else if (hs_in & ~is_compress & ~io_if2id_excep_en) begin // @[playground/src/noop/decode.scala 65:54]
      ctrl_r_dcMode <= instType_3; // @[playground/src/noop/decode.scala 71:27]
    end
    if (reset) begin // @[playground/src/noop/decode.scala 26:30]
      ctrl_r_writeRegEn <= 1'h0; // @[playground/src/noop/decode.scala 26:30]
    end else if (hs_in & io_if2id_excep_en) begin // @[playground/src/noop/decode.scala 302:37]
      ctrl_r_writeRegEn <= 1'h0; // @[playground/src/noop/decode.scala 306:25]
    end else if (hs_in & is_compress & _T_7) begin // @[playground/src/noop/decode.scala 199:53]
      ctrl_r_writeRegEn <= instType_c_5; // @[playground/src/noop/decode.scala 206:27]
    end else if (hs_in & ~is_compress & ~io_if2id_excep_en) begin // @[playground/src/noop/decode.scala 65:54]
      ctrl_r_writeRegEn <= instType_4; // @[playground/src/noop/decode.scala 72:27]
    end
    if (reset) begin // @[playground/src/noop/decode.scala 26:30]
      ctrl_r_writeCSREn <= 1'h0; // @[playground/src/noop/decode.scala 26:30]
    end else if (hs_in & io_if2id_excep_en) begin // @[playground/src/noop/decode.scala 302:37]
      ctrl_r_writeCSREn <= 1'h0; // @[playground/src/noop/decode.scala 306:25]
    end else if (hs_in & is_compress & _T_7) begin // @[playground/src/noop/decode.scala 199:53]
      ctrl_r_writeCSREn <= 1'h0; // @[playground/src/noop/decode.scala 207:27]
    end else if (hs_in & ~is_compress & ~io_if2id_excep_en) begin // @[playground/src/noop/decode.scala 65:54]
      ctrl_r_writeCSREn <= instType_6; // @[playground/src/noop/decode.scala 73:27]
    end
    if (reset) begin // @[playground/src/noop/decode.scala 26:30]
      ctrl_r_brType <= 3'h0; // @[playground/src/noop/decode.scala 26:30]
    end else if (hs_in & io_if2id_excep_en) begin // @[playground/src/noop/decode.scala 302:37]
      ctrl_r_brType <= 3'h0; // @[playground/src/noop/decode.scala 306:25]
    end else if (hs_in & is_compress & _T_7) begin // @[playground/src/noop/decode.scala 199:53]
      if (instType_c_0 == 4'h7) begin // @[playground/src/noop/decode.scala 279:29]
        ctrl_r_brType <= _GEN_172;
      end else begin
        ctrl_r_brType <= _GEN_109;
      end
    end else begin
      ctrl_r_brType <= _GEN_109;
    end
    if (reset) begin // @[playground/src/noop/decode.scala 27:30]
      rs1_r <= 5'h0; // @[playground/src/noop/decode.scala 27:30]
    end else if (hs_in & is_compress & _T_7) begin // @[playground/src/noop/decode.scala 199:53]
      if (instType_c_0 == 4'h7) begin // @[playground/src/noop/decode.scala 279:29]
        rs1_r <= {{1'd0}, _rs1_r_T_4}; // @[playground/src/noop/decode.scala 281:21]
      end else if (instType_c_0 == 4'h6) begin // @[playground/src/noop/decode.scala 268:29]
        rs1_r <= {{1'd0}, _rs1_r_T_4}; // @[playground/src/noop/decode.scala 270:21]
      end else begin
        rs1_r <= _GEN_158;
      end
    end else if (hs_in & ~is_compress & ~io_if2id_excep_en) begin // @[playground/src/noop/decode.scala 65:54]
      rs1_r <= io_if2id_inst[19:15]; // @[playground/src/noop/decode.scala 74:25]
    end
    if (reset) begin // @[playground/src/noop/decode.scala 28:30]
      rrs1_r <= 1'h0; // @[playground/src/noop/decode.scala 28:30]
    end else if (hs_in & io_if2id_excep_en) begin // @[playground/src/noop/decode.scala 302:37]
      rrs1_r <= 1'h0; // @[playground/src/noop/decode.scala 307:25]
    end else if (hs_in & is_compress & _T_7) begin // @[playground/src/noop/decode.scala 199:53]
      rrs1_r <= _GEN_175;
    end else if (hs_in & ~is_compress & ~io_if2id_excep_en) begin // @[playground/src/noop/decode.scala 65:54]
      rrs1_r <= _GEN_40;
    end
    if (reset) begin // @[playground/src/noop/decode.scala 29:30]
      rs1_d_r <= 64'h0; // @[playground/src/noop/decode.scala 29:30]
    end else if (hs_in & is_compress & _T_7) begin // @[playground/src/noop/decode.scala 199:53]
      if (instType_c_0 == 4'h8) begin // @[playground/src/noop/decode.scala 296:29]
        rs1_d_r <= io_if2id_pc; // @[playground/src/noop/decode.scala 297:21]
      end else begin
        rs1_d_r <= _GEN_108;
      end
    end else begin
      rs1_d_r <= _GEN_108;
    end
    if (reset) begin // @[playground/src/noop/decode.scala 30:30]
      rs2_r <= 12'h0; // @[playground/src/noop/decode.scala 30:30]
    end else if (hs_in & is_compress & _T_7) begin // @[playground/src/noop/decode.scala 199:53]
      rs2_r <= {{7'd0}, _GEN_165};
    end else if (hs_in & ~is_compress & ~io_if2id_excep_en) begin // @[playground/src/noop/decode.scala 65:54]
      if (32'h30200073 == io_if2id_inst) begin // @[playground/src/noop/decode.scala 159:37]
        rs2_r <= 12'h341; // @[playground/src/noop/decode.scala 166:25]
      end else begin
        rs2_r <= _GEN_65;
      end
    end
    if (reset) begin // @[playground/src/noop/decode.scala 31:30]
      rrs2_r <= 1'h0; // @[playground/src/noop/decode.scala 31:30]
    end else if (hs_in & io_if2id_excep_en) begin // @[playground/src/noop/decode.scala 302:37]
      rrs2_r <= 1'h0; // @[playground/src/noop/decode.scala 308:25]
    end else if (hs_in & is_compress & _T_7) begin // @[playground/src/noop/decode.scala 199:53]
      rrs2_r <= _GEN_164;
    end else if (hs_in & ~is_compress & ~io_if2id_excep_en) begin // @[playground/src/noop/decode.scala 65:54]
      rrs2_r <= _GEN_41;
    end
    if (reset) begin // @[playground/src/noop/decode.scala 32:30]
      rs2_d_r <= 64'h0; // @[playground/src/noop/decode.scala 32:30]
    end else if (hs_in & is_compress & _T_7) begin // @[playground/src/noop/decode.scala 199:53]
      if (instType_c_0 == 4'h7) begin // @[playground/src/noop/decode.scala 279:29]
        if (_instType_c_T_44) begin // @[playground/src/noop/decode.scala 290:36]
          rs2_d_r <= 64'h0; // @[playground/src/noop/decode.scala 292:29]
        end else begin
          rs2_d_r <= _GEN_170;
        end
      end else if (instType_c_0 == 4'h5) begin // @[playground/src/noop/decode.scala 262:29]
        rs2_d_r <= _rs2_d_r_T_7; // @[playground/src/noop/decode.scala 265:21]
      end else begin
        rs2_d_r <= _GEN_155;
      end
    end else if (hs_in & ~is_compress & ~io_if2id_excep_en) begin // @[playground/src/noop/decode.scala 65:54]
      if (instType_0 == 3'h6) begin // @[playground/src/noop/decode.scala 131:30]
        rs2_d_r <= _rs2_d_r_T_1; // @[playground/src/noop/decode.scala 133:25]
      end else begin
        rs2_d_r <= _GEN_46;
      end
    end
    if (reset) begin // @[playground/src/noop/decode.scala 33:30]
      dst_r <= 5'h0; // @[playground/src/noop/decode.scala 33:30]
    end else if (hs_in & is_compress & _T_7) begin // @[playground/src/noop/decode.scala 199:53]
      if (instType_c_0 == 4'h7) begin // @[playground/src/noop/decode.scala 279:29]
        dst_r <= {{1'd0}, _rs1_r_T_4}; // @[playground/src/noop/decode.scala 284:21]
      end else if (instType_c_0 == 4'h6) begin // @[playground/src/noop/decode.scala 268:29]
        dst_r <= {{1'd0}, _rs1_r_T_4}; // @[playground/src/noop/decode.scala 274:21]
      end else begin
        dst_r <= _GEN_160;
      end
    end else if (hs_in & ~is_compress & ~io_if2id_excep_en) begin // @[playground/src/noop/decode.scala 65:54]
      dst_r <= io_if2id_inst[11:7]; // @[playground/src/noop/decode.scala 78:25]
    end
    if (reset) begin // @[playground/src/noop/decode.scala 34:30]
      dst_d_r <= 64'h0; // @[playground/src/noop/decode.scala 34:30]
    end else if (hs_in & is_compress & _T_7) begin // @[playground/src/noop/decode.scala 199:53]
      if (instType_c_0 == 4'h8) begin // @[playground/src/noop/decode.scala 296:29]
        dst_d_r <= _rs2_d_r_T_7; // @[playground/src/noop/decode.scala 298:21]
      end else if (instType_c_0 == 4'h7) begin // @[playground/src/noop/decode.scala 279:29]
        dst_d_r <= _dst_d_r_T_13; // @[playground/src/noop/decode.scala 283:21]
      end else begin
        dst_d_r <= _GEN_166;
      end
    end else if (hs_in & ~is_compress & ~io_if2id_excep_en) begin // @[playground/src/noop/decode.scala 65:54]
      if (instType_0 == 3'h6) begin // @[playground/src/noop/decode.scala 131:30]
        dst_d_r <= 64'h0; // @[playground/src/noop/decode.scala 134:25]
      end else begin
        dst_d_r <= _GEN_42;
      end
    end
    if (reset) begin // @[playground/src/noop/decode.scala 35:30]
      jmp_type_r <= 2'h0; // @[playground/src/noop/decode.scala 35:30]
    end else if (hs_in & io_if2id_excep_en) begin // @[playground/src/noop/decode.scala 302:37]
      jmp_type_r <= 2'h0; // @[playground/src/noop/decode.scala 309:25]
    end else if (hs_in & is_compress & _T_7) begin // @[playground/src/noop/decode.scala 199:53]
      if (instType_c_0 == 4'h8) begin // @[playground/src/noop/decode.scala 296:29]
        jmp_type_r <= 2'h1; // @[playground/src/noop/decode.scala 299:25]
      end else begin
        jmp_type_r <= _GEN_181;
      end
    end else if (hs_in & ~is_compress & ~io_if2id_excep_en) begin // @[playground/src/noop/decode.scala 65:54]
      jmp_type_r <= _GEN_73;
    end
    if (reset) begin // @[playground/src/noop/decode.scala 36:30]
      special_r <= 2'h0; // @[playground/src/noop/decode.scala 36:30]
    end else if (hs_in & io_if2id_excep_en) begin // @[playground/src/noop/decode.scala 302:37]
      special_r <= 2'h0; // @[playground/src/noop/decode.scala 310:25]
    end else if (hs_in & is_compress & _T_7) begin // @[playground/src/noop/decode.scala 199:53]
      special_r <= 2'h0; // @[playground/src/noop/decode.scala 214:25]
    end else if (hs_in & ~is_compress & ~io_if2id_excep_en) begin // @[playground/src/noop/decode.scala 65:54]
      special_r <= _GEN_80;
    end
    if (reset) begin // @[playground/src/noop/decode.scala 37:30]
      swap_r <= 6'h0; // @[playground/src/noop/decode.scala 37:30]
    end else if (hs_in & io_if2id_excep_en) begin // @[playground/src/noop/decode.scala 302:37]
      swap_r <= 6'h1b; // @[playground/src/noop/decode.scala 312:25]
    end else if (hs_in & is_compress & _T_7) begin // @[playground/src/noop/decode.scala 199:53]
      if (instType_c_0 == 4'h6) begin // @[playground/src/noop/decode.scala 268:29]
        swap_r <= _GEN_161;
      end else begin
        swap_r <= _GEN_152;
      end
    end else if (hs_in & ~is_compress & ~io_if2id_excep_en) begin // @[playground/src/noop/decode.scala 65:54]
      swap_r <= _GEN_38;
    end
    if (reset) begin // @[playground/src/noop/decode.scala 38:30]
      indi_r <= 2'h0; // @[playground/src/noop/decode.scala 38:30]
    end else if (hs_in & io_if2id_excep_en) begin // @[playground/src/noop/decode.scala 302:37]
      indi_r <= 2'h0; // @[playground/src/noop/decode.scala 311:25]
    end else if (hs_in & is_compress & _T_7) begin // @[playground/src/noop/decode.scala 199:53]
      indi_r <= 2'h0; // @[playground/src/noop/decode.scala 215:25]
    end else if (hs_in & ~is_compress & ~io_if2id_excep_en) begin // @[playground/src/noop/decode.scala 65:54]
      indi_r <= _indi_r_T_10; // @[playground/src/noop/decode.scala 81:25]
    end
    if (reset) begin // @[playground/src/noop/decode.scala 39:30]
      recov_r <= 1'h0; // @[playground/src/noop/decode.scala 39:30]
    end else if (hs_in & io_if2id_excep_en) begin // @[playground/src/noop/decode.scala 302:37]
      recov_r <= io_if2id_recov; // @[playground/src/noop/decode.scala 313:25]
    end else if (hs_in & is_compress & _T_7) begin // @[playground/src/noop/decode.scala 199:53]
      recov_r <= _GEN_129;
    end else if (hs_in & ~is_compress & ~io_if2id_excep_en) begin // @[playground/src/noop/decode.scala 65:54]
      recov_r <= _GEN_82;
    end
    if (reset) begin // @[playground/src/noop/decode.scala 40:30]
      valid_r <= 1'h0; // @[playground/src/noop/decode.scala 40:30]
    end else begin
      valid_r <= _GEN_237;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  drop_r = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  stall_r = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  inst_r = _RAND_2[31:0];
  _RAND_3 = {2{`RANDOM}};
  pc_r = _RAND_3[63:0];
  _RAND_4 = {2{`RANDOM}};
  excep_r_cause = _RAND_4[63:0];
  _RAND_5 = {2{`RANDOM}};
  excep_r_tval = _RAND_5[63:0];
  _RAND_6 = {1{`RANDOM}};
  excep_r_en = _RAND_6[0:0];
  _RAND_7 = {2{`RANDOM}};
  excep_r_pc = _RAND_7[63:0];
  _RAND_8 = {1{`RANDOM}};
  excep_r_etype = _RAND_8[1:0];
  _RAND_9 = {1{`RANDOM}};
  ctrl_r_aluOp = _RAND_9[4:0];
  _RAND_10 = {1{`RANDOM}};
  ctrl_r_aluWidth = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  ctrl_r_dcMode = _RAND_11[4:0];
  _RAND_12 = {1{`RANDOM}};
  ctrl_r_writeRegEn = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  ctrl_r_writeCSREn = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  ctrl_r_brType = _RAND_14[2:0];
  _RAND_15 = {1{`RANDOM}};
  rs1_r = _RAND_15[4:0];
  _RAND_16 = {1{`RANDOM}};
  rrs1_r = _RAND_16[0:0];
  _RAND_17 = {2{`RANDOM}};
  rs1_d_r = _RAND_17[63:0];
  _RAND_18 = {1{`RANDOM}};
  rs2_r = _RAND_18[11:0];
  _RAND_19 = {1{`RANDOM}};
  rrs2_r = _RAND_19[0:0];
  _RAND_20 = {2{`RANDOM}};
  rs2_d_r = _RAND_20[63:0];
  _RAND_21 = {1{`RANDOM}};
  dst_r = _RAND_21[4:0];
  _RAND_22 = {2{`RANDOM}};
  dst_d_r = _RAND_22[63:0];
  _RAND_23 = {1{`RANDOM}};
  jmp_type_r = _RAND_23[1:0];
  _RAND_24 = {1{`RANDOM}};
  special_r = _RAND_24[1:0];
  _RAND_25 = {1{`RANDOM}};
  swap_r = _RAND_25[5:0];
  _RAND_26 = {1{`RANDOM}};
  indi_r = _RAND_26[1:0];
  _RAND_27 = {1{`RANDOM}};
  recov_r = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  valid_r = _RAND_28[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Forwarding(
  input         clock,
  input         reset,
  input  [31:0] io_id2df_inst, // @[playground/src/noop/forwading.scala 10:16]
  input  [63:0] io_id2df_pc, // @[playground/src/noop/forwading.scala 10:16]
  input  [63:0] io_id2df_excep_cause, // @[playground/src/noop/forwading.scala 10:16]
  input  [63:0] io_id2df_excep_tval, // @[playground/src/noop/forwading.scala 10:16]
  input         io_id2df_excep_en, // @[playground/src/noop/forwading.scala 10:16]
  input  [63:0] io_id2df_excep_pc, // @[playground/src/noop/forwading.scala 10:16]
  input  [1:0]  io_id2df_excep_etype, // @[playground/src/noop/forwading.scala 10:16]
  input  [4:0]  io_id2df_ctrl_aluOp, // @[playground/src/noop/forwading.scala 10:16]
  input         io_id2df_ctrl_aluWidth, // @[playground/src/noop/forwading.scala 10:16]
  input  [4:0]  io_id2df_ctrl_dcMode, // @[playground/src/noop/forwading.scala 10:16]
  input         io_id2df_ctrl_writeRegEn, // @[playground/src/noop/forwading.scala 10:16]
  input         io_id2df_ctrl_writeCSREn, // @[playground/src/noop/forwading.scala 10:16]
  input  [2:0]  io_id2df_ctrl_brType, // @[playground/src/noop/forwading.scala 10:16]
  input  [4:0]  io_id2df_rs1, // @[playground/src/noop/forwading.scala 10:16]
  input         io_id2df_rrs1, // @[playground/src/noop/forwading.scala 10:16]
  input  [63:0] io_id2df_rs1_d, // @[playground/src/noop/forwading.scala 10:16]
  input  [11:0] io_id2df_rs2, // @[playground/src/noop/forwading.scala 10:16]
  input         io_id2df_rrs2, // @[playground/src/noop/forwading.scala 10:16]
  input  [63:0] io_id2df_rs2_d, // @[playground/src/noop/forwading.scala 10:16]
  input  [4:0]  io_id2df_dst, // @[playground/src/noop/forwading.scala 10:16]
  input  [63:0] io_id2df_dst_d, // @[playground/src/noop/forwading.scala 10:16]
  input  [1:0]  io_id2df_jmp_type, // @[playground/src/noop/forwading.scala 10:16]
  input  [1:0]  io_id2df_special, // @[playground/src/noop/forwading.scala 10:16]
  input  [5:0]  io_id2df_swap, // @[playground/src/noop/forwading.scala 10:16]
  input  [1:0]  io_id2df_indi, // @[playground/src/noop/forwading.scala 10:16]
  output        io_id2df_drop, // @[playground/src/noop/forwading.scala 10:16]
  output        io_id2df_stall, // @[playground/src/noop/forwading.scala 10:16]
  input         io_id2df_recov, // @[playground/src/noop/forwading.scala 10:16]
  input         io_id2df_valid, // @[playground/src/noop/forwading.scala 10:16]
  output        io_id2df_ready, // @[playground/src/noop/forwading.scala 10:16]
  output [31:0] io_df2rr_inst, // @[playground/src/noop/forwading.scala 10:16]
  output [63:0] io_df2rr_pc, // @[playground/src/noop/forwading.scala 10:16]
  output [63:0] io_df2rr_excep_cause, // @[playground/src/noop/forwading.scala 10:16]
  output [63:0] io_df2rr_excep_tval, // @[playground/src/noop/forwading.scala 10:16]
  output        io_df2rr_excep_en, // @[playground/src/noop/forwading.scala 10:16]
  output [63:0] io_df2rr_excep_pc, // @[playground/src/noop/forwading.scala 10:16]
  output [1:0]  io_df2rr_excep_etype, // @[playground/src/noop/forwading.scala 10:16]
  output [4:0]  io_df2rr_ctrl_aluOp, // @[playground/src/noop/forwading.scala 10:16]
  output        io_df2rr_ctrl_aluWidth, // @[playground/src/noop/forwading.scala 10:16]
  output [4:0]  io_df2rr_ctrl_dcMode, // @[playground/src/noop/forwading.scala 10:16]
  output        io_df2rr_ctrl_writeRegEn, // @[playground/src/noop/forwading.scala 10:16]
  output        io_df2rr_ctrl_writeCSREn, // @[playground/src/noop/forwading.scala 10:16]
  output [2:0]  io_df2rr_ctrl_brType, // @[playground/src/noop/forwading.scala 10:16]
  output [4:0]  io_df2rr_rs1, // @[playground/src/noop/forwading.scala 10:16]
  output        io_df2rr_rrs1, // @[playground/src/noop/forwading.scala 10:16]
  output [63:0] io_df2rr_rs1_d, // @[playground/src/noop/forwading.scala 10:16]
  output [11:0] io_df2rr_rs2, // @[playground/src/noop/forwading.scala 10:16]
  output        io_df2rr_rrs2, // @[playground/src/noop/forwading.scala 10:16]
  output [63:0] io_df2rr_rs2_d, // @[playground/src/noop/forwading.scala 10:16]
  output [4:0]  io_df2rr_dst, // @[playground/src/noop/forwading.scala 10:16]
  output [63:0] io_df2rr_dst_d, // @[playground/src/noop/forwading.scala 10:16]
  output [1:0]  io_df2rr_jmp_type, // @[playground/src/noop/forwading.scala 10:16]
  output [1:0]  io_df2rr_special, // @[playground/src/noop/forwading.scala 10:16]
  output [5:0]  io_df2rr_swap, // @[playground/src/noop/forwading.scala 10:16]
  output [1:0]  io_df2rr_indi, // @[playground/src/noop/forwading.scala 10:16]
  input         io_df2rr_drop, // @[playground/src/noop/forwading.scala 10:16]
  input         io_df2rr_stall, // @[playground/src/noop/forwading.scala 10:16]
  output        io_df2rr_recov, // @[playground/src/noop/forwading.scala 10:16]
  output        io_df2rr_valid, // @[playground/src/noop/forwading.scala 10:16]
  input         io_df2rr_ready, // @[playground/src/noop/forwading.scala 10:16]
  input  [4:0]  io_d_rr_id, // @[playground/src/noop/forwading.scala 10:16]
  input  [63:0] io_d_rr_data, // @[playground/src/noop/forwading.scala 10:16]
  input  [1:0]  io_d_rr_state, // @[playground/src/noop/forwading.scala 10:16]
  input  [4:0]  io_d_ex_id, // @[playground/src/noop/forwading.scala 10:16]
  input  [63:0] io_d_ex_data, // @[playground/src/noop/forwading.scala 10:16]
  input  [1:0]  io_d_ex_state, // @[playground/src/noop/forwading.scala 10:16]
  input  [4:0]  io_d_mem1_id, // @[playground/src/noop/forwading.scala 10:16]
  input  [63:0] io_d_mem1_data, // @[playground/src/noop/forwading.scala 10:16]
  input  [1:0]  io_d_mem1_state, // @[playground/src/noop/forwading.scala 10:16]
  input  [4:0]  io_d_mem2_id, // @[playground/src/noop/forwading.scala 10:16]
  input  [63:0] io_d_mem2_data, // @[playground/src/noop/forwading.scala 10:16]
  input  [1:0]  io_d_mem2_state, // @[playground/src/noop/forwading.scala 10:16]
  input  [4:0]  io_d_mem3_id, // @[playground/src/noop/forwading.scala 10:16]
  input  [63:0] io_d_mem3_data, // @[playground/src/noop/forwading.scala 10:16]
  input  [1:0]  io_d_mem3_state // @[playground/src/noop/forwading.scala 10:16]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [63:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [63:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [63:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
`endif // RANDOMIZE_REG_INIT
  wire  _io_id2df_stall_T = ~io_df2rr_drop; // @[playground/src/noop/forwading.scala 23:36]
  reg [31:0] inst_r; // @[playground/src/noop/forwading.scala 24:30]
  reg [63:0] pc_r; // @[playground/src/noop/forwading.scala 25:30]
  reg [63:0] excep_r_cause; // @[playground/src/noop/forwading.scala 26:30]
  reg [63:0] excep_r_tval; // @[playground/src/noop/forwading.scala 26:30]
  reg  excep_r_en; // @[playground/src/noop/forwading.scala 26:30]
  reg [63:0] excep_r_pc; // @[playground/src/noop/forwading.scala 26:30]
  reg [1:0] excep_r_etype; // @[playground/src/noop/forwading.scala 26:30]
  reg [4:0] ctrl_r_aluOp; // @[playground/src/noop/forwading.scala 27:30]
  reg  ctrl_r_aluWidth; // @[playground/src/noop/forwading.scala 27:30]
  reg [4:0] ctrl_r_dcMode; // @[playground/src/noop/forwading.scala 27:30]
  reg  ctrl_r_writeRegEn; // @[playground/src/noop/forwading.scala 27:30]
  reg  ctrl_r_writeCSREn; // @[playground/src/noop/forwading.scala 27:30]
  reg [2:0] ctrl_r_brType; // @[playground/src/noop/forwading.scala 27:30]
  reg [4:0] rs1_r; // @[playground/src/noop/forwading.scala 28:30]
  reg  rrs1_r; // @[playground/src/noop/forwading.scala 29:30]
  reg [63:0] rs1_d_r; // @[playground/src/noop/forwading.scala 30:30]
  reg [11:0] rs2_r; // @[playground/src/noop/forwading.scala 31:30]
  reg  rrs2_r; // @[playground/src/noop/forwading.scala 32:30]
  reg [63:0] rs2_d_r; // @[playground/src/noop/forwading.scala 33:30]
  reg [4:0] dst_r; // @[playground/src/noop/forwading.scala 34:30]
  reg [63:0] dst_d_r; // @[playground/src/noop/forwading.scala 35:30]
  reg [1:0] jmp_type_r; // @[playground/src/noop/forwading.scala 36:30]
  reg [1:0] special_r; // @[playground/src/noop/forwading.scala 37:30]
  reg [1:0] indi_r; // @[playground/src/noop/forwading.scala 38:30]
  reg [5:0] swap_r; // @[playground/src/noop/forwading.scala 39:30]
  reg  recov_r; // @[playground/src/noop/forwading.scala 40:30]
  reg  valid_r; // @[playground/src/noop/forwading.scala 41:30]
  reg [4:0] pre_dst; // @[playground/src/noop/forwading.scala 43:30]
  reg  pre_wr; // @[playground/src/noop/forwading.scala 44:30]
  reg  state; // @[playground/src/noop/forwading.scala 47:24]
  wire  hs_in = io_id2df_ready & io_id2df_valid; // @[playground/src/noop/forwading.scala 48:34]
  wire  hs_out = io_df2rr_ready & io_df2rr_valid; // @[playground/src/noop/forwading.scala 49:34]
  wire [4:0] cur_rs1 = hs_in ? io_id2df_rs1 : rs1_r; // @[playground/src/noop/forwading.scala 59:26]
  wire  cur_rrs1 = hs_in ? io_id2df_rrs1 : rrs1_r; // @[playground/src/noop/forwading.scala 60:26]
  wire [11:0] cur_rs2 = hs_in ? io_id2df_rs2 : rs2_r; // @[playground/src/noop/forwading.scala 61:26]
  wire  cur_rrs2 = hs_in ? io_id2df_rrs2 : rrs2_r; // @[playground/src/noop/forwading.scala 62:26]
  wire  _T_1 = valid_r & pre_wr; // @[playground/src/noop/forwading.scala 67:28]
  wire  _T_5 = io_d_rr_state != 2'h0; // @[playground/src/noop/forwading.scala 69:63]
  wire  _T_7 = io_d_rr_state == 2'h1; // @[playground/src/noop/forwading.scala 70:32]
  wire [63:0] _GEN_0 = io_d_rr_state == 2'h1 ? io_d_rr_data : 64'h0; // @[playground/src/noop/forwading.scala 70:44 71:26 57:62]
  wire  _GEN_2 = io_d_rr_state == 2'h1 ? 1'h0 : 1'h1; // @[playground/src/noop/forwading.scala 57:41 70:44 74:26]
  wire  _T_9 = io_d_ex_state != 2'h0; // @[playground/src/noop/forwading.scala 76:63]
  wire  _T_11 = io_d_ex_state == 2'h1; // @[playground/src/noop/forwading.scala 77:32]
  wire [63:0] _GEN_3 = io_d_ex_state == 2'h1 ? io_d_ex_data : 64'h0; // @[playground/src/noop/forwading.scala 77:44 78:26 57:62]
  wire  _GEN_5 = io_d_ex_state == 2'h1 ? 1'h0 : 1'h1; // @[playground/src/noop/forwading.scala 57:41 77:44 81:26]
  wire  _T_13 = io_d_mem1_state != 2'h0; // @[playground/src/noop/forwading.scala 83:67]
  wire  _T_15 = io_d_mem1_state == 2'h1; // @[playground/src/noop/forwading.scala 84:34]
  wire [63:0] _GEN_6 = io_d_mem1_state == 2'h1 ? io_d_mem1_data : 64'h0; // @[playground/src/noop/forwading.scala 84:46 85:26 57:62]
  wire  _GEN_8 = io_d_mem1_state == 2'h1 ? 1'h0 : 1'h1; // @[playground/src/noop/forwading.scala 57:41 84:46 88:26]
  wire  _T_17 = io_d_mem2_state != 2'h0; // @[playground/src/noop/forwading.scala 90:67]
  wire  _T_19 = io_d_mem2_state == 2'h1; // @[playground/src/noop/forwading.scala 91:34]
  wire [63:0] _GEN_9 = io_d_mem2_state == 2'h1 ? io_d_mem2_data : 64'h0; // @[playground/src/noop/forwading.scala 91:46 92:26 57:62]
  wire  _GEN_11 = io_d_mem2_state == 2'h1 ? 1'h0 : 1'h1; // @[playground/src/noop/forwading.scala 57:41 91:46 95:26]
  wire  _T_21 = io_d_mem3_state != 2'h0; // @[playground/src/noop/forwading.scala 97:67]
  wire  _T_23 = io_d_mem3_state == 2'h1; // @[playground/src/noop/forwading.scala 98:34]
  wire [63:0] _GEN_12 = io_d_mem3_state == 2'h1 ? io_d_mem3_data : 64'h0; // @[playground/src/noop/forwading.scala 98:46 99:26 57:62]
  wire  _GEN_14 = io_d_mem3_state == 2'h1 ? 1'h0 : 1'h1; // @[playground/src/noop/forwading.scala 102:26 57:41 98:46]
  wire [63:0] _GEN_15 = cur_rs1 == io_d_mem3_id & io_d_mem3_state != 2'h0 ? _GEN_12 : 64'h0; // @[playground/src/noop/forwading.scala 57:62 97:82]
  wire  _GEN_16 = cur_rs1 == io_d_mem3_id & io_d_mem3_state != 2'h0 & _T_23; // @[playground/src/noop/forwading.scala 57:15 97:82]
  wire  _GEN_17 = cur_rs1 == io_d_mem3_id & io_d_mem3_state != 2'h0 & _GEN_14; // @[playground/src/noop/forwading.scala 57:41 97:82]
  wire [63:0] _GEN_18 = cur_rs1 == io_d_mem2_id & io_d_mem2_state != 2'h0 ? _GEN_9 : _GEN_15; // @[playground/src/noop/forwading.scala 90:82]
  wire  _GEN_19 = cur_rs1 == io_d_mem2_id & io_d_mem2_state != 2'h0 ? _T_19 : _GEN_16; // @[playground/src/noop/forwading.scala 90:82]
  wire  _GEN_20 = cur_rs1 == io_d_mem2_id & io_d_mem2_state != 2'h0 ? _GEN_11 : _GEN_17; // @[playground/src/noop/forwading.scala 90:82]
  wire [63:0] _GEN_21 = cur_rs1 == io_d_mem1_id & io_d_mem1_state != 2'h0 ? _GEN_6 : _GEN_18; // @[playground/src/noop/forwading.scala 83:82]
  wire  _GEN_22 = cur_rs1 == io_d_mem1_id & io_d_mem1_state != 2'h0 ? _T_15 : _GEN_19; // @[playground/src/noop/forwading.scala 83:82]
  wire  _GEN_23 = cur_rs1 == io_d_mem1_id & io_d_mem1_state != 2'h0 ? _GEN_8 : _GEN_20; // @[playground/src/noop/forwading.scala 83:82]
  wire [63:0] _GEN_24 = cur_rs1 == io_d_ex_id & io_d_ex_state != 2'h0 ? _GEN_3 : _GEN_21; // @[playground/src/noop/forwading.scala 76:78]
  wire  _GEN_25 = cur_rs1 == io_d_ex_id & io_d_ex_state != 2'h0 ? _T_11 : _GEN_22; // @[playground/src/noop/forwading.scala 76:78]
  wire  _GEN_26 = cur_rs1 == io_d_ex_id & io_d_ex_state != 2'h0 ? _GEN_5 : _GEN_23; // @[playground/src/noop/forwading.scala 76:78]
  wire [63:0] _GEN_27 = cur_rs1 == io_d_rr_id & io_d_rr_state != 2'h0 ? _GEN_0 : _GEN_24; // @[playground/src/noop/forwading.scala 69:78]
  wire  _GEN_28 = cur_rs1 == io_d_rr_id & io_d_rr_state != 2'h0 ? _T_7 : _GEN_25; // @[playground/src/noop/forwading.scala 69:78]
  wire  _GEN_29 = cur_rs1 == io_d_rr_id & io_d_rr_state != 2'h0 ? _GEN_2 : _GEN_26; // @[playground/src/noop/forwading.scala 69:78]
  wire  _GEN_30 = valid_r & pre_wr & cur_rs1 == pre_dst | _GEN_29; // @[playground/src/noop/forwading.scala 67:59 68:22]
  wire [63:0] _GEN_31 = valid_r & pre_wr & cur_rs1 == pre_dst ? 64'h0 : _GEN_27; // @[playground/src/noop/forwading.scala 67:59 57:62]
  wire  _GEN_32 = valid_r & pre_wr & cur_rs1 == pre_dst ? 1'h0 : _GEN_28; // @[playground/src/noop/forwading.scala 57:15 67:59]
  wire  _GEN_33 = cur_rs1 == 5'h0 ? 1'h0 : _GEN_30; // @[playground/src/noop/forwading.scala 65:30 66:22]
  wire [63:0] _GEN_34 = cur_rs1 == 5'h0 ? 64'h0 : _GEN_31; // @[playground/src/noop/forwading.scala 65:30 57:62]
  wire  _GEN_35 = cur_rs1 == 5'h0 ? 1'h0 : _GEN_32; // @[playground/src/noop/forwading.scala 57:15 65:30]
  wire  rs1_wait = cur_rrs1 & _GEN_33; // @[playground/src/noop/forwading.scala 63:19 57:41]
  wire  rs1_valid = cur_rrs1 & _GEN_35; // @[playground/src/noop/forwading.scala 57:15 63:19]
  wire [11:0] _GEN_130 = {{7'd0}, pre_dst}; // @[playground/src/noop/forwading.scala 110:48]
  wire [11:0] _GEN_131 = {{7'd0}, io_d_rr_id}; // @[playground/src/noop/forwading.scala 112:29]
  wire [11:0] _GEN_132 = {{7'd0}, io_d_ex_id}; // @[playground/src/noop/forwading.scala 119:29]
  wire [11:0] _GEN_133 = {{7'd0}, io_d_mem1_id}; // @[playground/src/noop/forwading.scala 126:29]
  wire [11:0] _GEN_134 = {{7'd0}, io_d_mem2_id}; // @[playground/src/noop/forwading.scala 133:29]
  wire [11:0] _GEN_135 = {{7'd0}, io_d_mem3_id}; // @[playground/src/noop/forwading.scala 140:29]
  wire [63:0] _GEN_54 = cur_rs2 == _GEN_135 & _T_21 ? _GEN_12 : 64'h0; // @[playground/src/noop/forwading.scala 140:82 58:62]
  wire  _GEN_55 = cur_rs2 == _GEN_135 & _T_21 & _T_23; // @[playground/src/noop/forwading.scala 140:82 58:15]
  wire  _GEN_56 = cur_rs2 == _GEN_135 & _T_21 & _GEN_14; // @[playground/src/noop/forwading.scala 140:82 58:41]
  wire [63:0] _GEN_57 = cur_rs2 == _GEN_134 & _T_17 ? _GEN_9 : _GEN_54; // @[playground/src/noop/forwading.scala 133:82]
  wire  _GEN_58 = cur_rs2 == _GEN_134 & _T_17 ? _T_19 : _GEN_55; // @[playground/src/noop/forwading.scala 133:82]
  wire  _GEN_59 = cur_rs2 == _GEN_134 & _T_17 ? _GEN_11 : _GEN_56; // @[playground/src/noop/forwading.scala 133:82]
  wire [63:0] _GEN_60 = cur_rs2 == _GEN_133 & _T_13 ? _GEN_6 : _GEN_57; // @[playground/src/noop/forwading.scala 126:82]
  wire  _GEN_61 = cur_rs2 == _GEN_133 & _T_13 ? _T_15 : _GEN_58; // @[playground/src/noop/forwading.scala 126:82]
  wire  _GEN_62 = cur_rs2 == _GEN_133 & _T_13 ? _GEN_8 : _GEN_59; // @[playground/src/noop/forwading.scala 126:82]
  wire [63:0] _GEN_63 = cur_rs2 == _GEN_132 & _T_9 ? _GEN_3 : _GEN_60; // @[playground/src/noop/forwading.scala 119:78]
  wire  _GEN_64 = cur_rs2 == _GEN_132 & _T_9 ? _T_11 : _GEN_61; // @[playground/src/noop/forwading.scala 119:78]
  wire  _GEN_65 = cur_rs2 == _GEN_132 & _T_9 ? _GEN_5 : _GEN_62; // @[playground/src/noop/forwading.scala 119:78]
  wire [63:0] _GEN_66 = cur_rs2 == _GEN_131 & _T_5 ? _GEN_0 : _GEN_63; // @[playground/src/noop/forwading.scala 112:78]
  wire  _GEN_67 = cur_rs2 == _GEN_131 & _T_5 ? _T_7 : _GEN_64; // @[playground/src/noop/forwading.scala 112:78]
  wire  _GEN_68 = cur_rs2 == _GEN_131 & _T_5 ? _GEN_2 : _GEN_65; // @[playground/src/noop/forwading.scala 112:78]
  wire  _GEN_69 = _T_1 & cur_rs2 == _GEN_130 | _GEN_68; // @[playground/src/noop/forwading.scala 110:60 111:22]
  wire [63:0] _GEN_70 = _T_1 & cur_rs2 == _GEN_130 ? 64'h0 : _GEN_66; // @[playground/src/noop/forwading.scala 110:60 58:62]
  wire  _GEN_71 = _T_1 & cur_rs2 == _GEN_130 ? 1'h0 : _GEN_67; // @[playground/src/noop/forwading.scala 110:60 58:15]
  wire  _GEN_72 = cur_rs2 == 12'h0 ? 1'h0 : _GEN_69; // @[playground/src/noop/forwading.scala 108:30 109:22]
  wire [63:0] _GEN_73 = cur_rs2 == 12'h0 ? 64'h0 : _GEN_70; // @[playground/src/noop/forwading.scala 108:30 58:62]
  wire  _GEN_74 = cur_rs2 == 12'h0 ? 1'h0 : _GEN_71; // @[playground/src/noop/forwading.scala 108:30 58:15]
  wire  rs2_wait = cur_rrs2 & _GEN_72; // @[playground/src/noop/forwading.scala 106:19 58:41]
  wire  rs2_valid = cur_rrs2 & _GEN_74; // @[playground/src/noop/forwading.scala 106:19 58:15]
  wire [63:0] _GEN_93 = hs_in ? io_id2df_rs1_d : rs1_d_r; // @[playground/src/noop/forwading.scala 150:16 157:21 30:30]
  wire [63:0] _GEN_96 = hs_in ? io_id2df_rs2_d : rs2_d_r; // @[playground/src/noop/forwading.scala 150:16 160:21 33:30]
  wire  _GEN_116 = (valid_r | state) & ~hs_out ? 1'h0 : io_id2df_valid; // @[playground/src/noop/forwading.scala 189:20 191:54]
  wire  _GEN_117 = hs_out ? 1'h0 : valid_r; // @[playground/src/noop/forwading.scala 202:31 203:25 41:30]
  wire  _GEN_118 = hs_in | _GEN_117; // @[playground/src/noop/forwading.scala 200:30 201:25]
  wire  _GEN_119 = hs_in & (rs1_wait | rs2_wait) | state; // @[playground/src/noop/forwading.scala 197:50 198:23 47:24]
  wire  _GEN_120 = hs_in & (rs1_wait | rs2_wait) ? 1'h0 : _GEN_118; // @[playground/src/noop/forwading.scala 197:50 199:25]
  wire  _GEN_121 = ~state ? _GEN_119 : state; // @[playground/src/noop/forwading.scala 196:30 47:24]
  wire  _GEN_122 = ~state ? _GEN_120 : valid_r; // @[playground/src/noop/forwading.scala 196:30 41:30]
  wire  _GEN_123 = ~rs1_wait & ~rs2_wait ? 1'h0 : _GEN_121; // @[playground/src/noop/forwading.scala 207:43 208:23]
  wire  _GEN_124 = ~rs1_wait & ~rs2_wait | _GEN_122; // @[playground/src/noop/forwading.scala 207:43 209:25]
  wire  _GEN_125 = state ? _GEN_123 : _GEN_121; // @[playground/src/noop/forwading.scala 206:30]
  wire  _GEN_126 = state ? _GEN_124 : _GEN_122; // @[playground/src/noop/forwading.scala 206:30]
  wire  _GEN_128 = _io_id2df_stall_T & _GEN_125; // @[playground/src/noop/forwading.scala 190:25 214:21]
  wire  _GEN_129 = _io_id2df_stall_T & _GEN_126; // @[playground/src/noop/forwading.scala 190:25 215:21]
  assign io_id2df_drop = io_df2rr_drop; // @[playground/src/noop/forwading.scala 22:31]
  assign io_id2df_stall = io_df2rr_stall; // @[playground/src/noop/forwading.scala 23:52]
  assign io_id2df_ready = _io_id2df_stall_T & _GEN_116; // @[playground/src/noop/forwading.scala 189:20 190:25]
  assign io_df2rr_inst = inst_r; // @[playground/src/noop/forwading.scala 217:25]
  assign io_df2rr_pc = pc_r; // @[playground/src/noop/forwading.scala 218:25]
  assign io_df2rr_excep_cause = excep_r_cause; // @[playground/src/noop/forwading.scala 219:25]
  assign io_df2rr_excep_tval = excep_r_tval; // @[playground/src/noop/forwading.scala 219:25]
  assign io_df2rr_excep_en = excep_r_en; // @[playground/src/noop/forwading.scala 219:25]
  assign io_df2rr_excep_pc = excep_r_pc; // @[playground/src/noop/forwading.scala 219:25]
  assign io_df2rr_excep_etype = excep_r_etype; // @[playground/src/noop/forwading.scala 219:25]
  assign io_df2rr_ctrl_aluOp = ctrl_r_aluOp; // @[playground/src/noop/forwading.scala 220:25]
  assign io_df2rr_ctrl_aluWidth = ctrl_r_aluWidth; // @[playground/src/noop/forwading.scala 220:25]
  assign io_df2rr_ctrl_dcMode = ctrl_r_dcMode; // @[playground/src/noop/forwading.scala 220:25]
  assign io_df2rr_ctrl_writeRegEn = ctrl_r_writeRegEn; // @[playground/src/noop/forwading.scala 220:25]
  assign io_df2rr_ctrl_writeCSREn = ctrl_r_writeCSREn; // @[playground/src/noop/forwading.scala 220:25]
  assign io_df2rr_ctrl_brType = ctrl_r_brType; // @[playground/src/noop/forwading.scala 220:25]
  assign io_df2rr_rs1 = rs1_r; // @[playground/src/noop/forwading.scala 221:25]
  assign io_df2rr_rrs1 = rrs1_r; // @[playground/src/noop/forwading.scala 222:25]
  assign io_df2rr_rs1_d = rs1_d_r; // @[playground/src/noop/forwading.scala 223:25]
  assign io_df2rr_rs2 = rs2_r; // @[playground/src/noop/forwading.scala 224:25]
  assign io_df2rr_rrs2 = rrs2_r; // @[playground/src/noop/forwading.scala 225:25]
  assign io_df2rr_rs2_d = rs2_d_r; // @[playground/src/noop/forwading.scala 226:25]
  assign io_df2rr_dst = dst_r; // @[playground/src/noop/forwading.scala 227:25]
  assign io_df2rr_dst_d = dst_d_r; // @[playground/src/noop/forwading.scala 228:25]
  assign io_df2rr_jmp_type = jmp_type_r; // @[playground/src/noop/forwading.scala 229:25]
  assign io_df2rr_special = special_r; // @[playground/src/noop/forwading.scala 230:25]
  assign io_df2rr_swap = swap_r; // @[playground/src/noop/forwading.scala 232:25]
  assign io_df2rr_indi = indi_r; // @[playground/src/noop/forwading.scala 231:25]
  assign io_df2rr_recov = recov_r; // @[playground/src/noop/forwading.scala 233:25]
  assign io_df2rr_valid = valid_r; // @[playground/src/noop/forwading.scala 234:25]
  always @(posedge clock) begin
    if (reset) begin // @[playground/src/noop/forwading.scala 24:30]
      inst_r <= 32'h0; // @[playground/src/noop/forwading.scala 24:30]
    end else if (hs_in) begin // @[playground/src/noop/forwading.scala 150:16]
      inst_r <= io_id2df_inst; // @[playground/src/noop/forwading.scala 151:21]
    end
    if (reset) begin // @[playground/src/noop/forwading.scala 25:30]
      pc_r <= 64'h0; // @[playground/src/noop/forwading.scala 25:30]
    end else if (hs_in) begin // @[playground/src/noop/forwading.scala 150:16]
      pc_r <= io_id2df_pc; // @[playground/src/noop/forwading.scala 152:21]
    end
    if (reset) begin // @[playground/src/noop/forwading.scala 26:30]
      excep_r_cause <= 64'h0; // @[playground/src/noop/forwading.scala 26:30]
    end else if (hs_in) begin // @[playground/src/noop/forwading.scala 150:16]
      excep_r_cause <= io_id2df_excep_cause; // @[playground/src/noop/forwading.scala 153:21]
    end
    if (reset) begin // @[playground/src/noop/forwading.scala 26:30]
      excep_r_tval <= 64'h0; // @[playground/src/noop/forwading.scala 26:30]
    end else if (hs_in) begin // @[playground/src/noop/forwading.scala 150:16]
      excep_r_tval <= io_id2df_excep_tval; // @[playground/src/noop/forwading.scala 153:21]
    end
    if (reset) begin // @[playground/src/noop/forwading.scala 26:30]
      excep_r_en <= 1'h0; // @[playground/src/noop/forwading.scala 26:30]
    end else if (hs_in) begin // @[playground/src/noop/forwading.scala 150:16]
      excep_r_en <= io_id2df_excep_en; // @[playground/src/noop/forwading.scala 153:21]
    end
    if (reset) begin // @[playground/src/noop/forwading.scala 26:30]
      excep_r_pc <= 64'h0; // @[playground/src/noop/forwading.scala 26:30]
    end else if (hs_in) begin // @[playground/src/noop/forwading.scala 150:16]
      excep_r_pc <= io_id2df_excep_pc; // @[playground/src/noop/forwading.scala 153:21]
    end
    if (reset) begin // @[playground/src/noop/forwading.scala 26:30]
      excep_r_etype <= 2'h0; // @[playground/src/noop/forwading.scala 26:30]
    end else if (hs_in) begin // @[playground/src/noop/forwading.scala 150:16]
      excep_r_etype <= io_id2df_excep_etype; // @[playground/src/noop/forwading.scala 153:21]
    end
    if (reset) begin // @[playground/src/noop/forwading.scala 27:30]
      ctrl_r_aluOp <= 5'h0; // @[playground/src/noop/forwading.scala 27:30]
    end else if (hs_in) begin // @[playground/src/noop/forwading.scala 150:16]
      ctrl_r_aluOp <= io_id2df_ctrl_aluOp; // @[playground/src/noop/forwading.scala 154:21]
    end
    if (reset) begin // @[playground/src/noop/forwading.scala 27:30]
      ctrl_r_aluWidth <= 1'h0; // @[playground/src/noop/forwading.scala 27:30]
    end else if (hs_in) begin // @[playground/src/noop/forwading.scala 150:16]
      ctrl_r_aluWidth <= io_id2df_ctrl_aluWidth; // @[playground/src/noop/forwading.scala 154:21]
    end
    if (reset) begin // @[playground/src/noop/forwading.scala 27:30]
      ctrl_r_dcMode <= 5'h0; // @[playground/src/noop/forwading.scala 27:30]
    end else if (hs_in) begin // @[playground/src/noop/forwading.scala 150:16]
      ctrl_r_dcMode <= io_id2df_ctrl_dcMode; // @[playground/src/noop/forwading.scala 154:21]
    end
    if (reset) begin // @[playground/src/noop/forwading.scala 27:30]
      ctrl_r_writeRegEn <= 1'h0; // @[playground/src/noop/forwading.scala 27:30]
    end else if (hs_in) begin // @[playground/src/noop/forwading.scala 150:16]
      ctrl_r_writeRegEn <= io_id2df_ctrl_writeRegEn; // @[playground/src/noop/forwading.scala 154:21]
    end
    if (reset) begin // @[playground/src/noop/forwading.scala 27:30]
      ctrl_r_writeCSREn <= 1'h0; // @[playground/src/noop/forwading.scala 27:30]
    end else if (hs_in) begin // @[playground/src/noop/forwading.scala 150:16]
      ctrl_r_writeCSREn <= io_id2df_ctrl_writeCSREn; // @[playground/src/noop/forwading.scala 154:21]
    end
    if (reset) begin // @[playground/src/noop/forwading.scala 27:30]
      ctrl_r_brType <= 3'h0; // @[playground/src/noop/forwading.scala 27:30]
    end else if (hs_in) begin // @[playground/src/noop/forwading.scala 150:16]
      ctrl_r_brType <= io_id2df_ctrl_brType; // @[playground/src/noop/forwading.scala 154:21]
    end
    if (reset) begin // @[playground/src/noop/forwading.scala 28:30]
      rs1_r <= 5'h0; // @[playground/src/noop/forwading.scala 28:30]
    end else if (hs_in) begin // @[playground/src/noop/forwading.scala 59:26]
      rs1_r <= io_id2df_rs1;
    end
    if (reset) begin // @[playground/src/noop/forwading.scala 29:30]
      rrs1_r <= 1'h0; // @[playground/src/noop/forwading.scala 29:30]
    end else if (hs_in | state) begin // @[playground/src/noop/forwading.scala 170:37]
      if (rs1_valid & cur_rrs1) begin // @[playground/src/noop/forwading.scala 171:36]
        rrs1_r <= 1'h0; // @[playground/src/noop/forwading.scala 172:21]
      end else begin
        rrs1_r <= cur_rrs1;
      end
    end else begin
      rrs1_r <= cur_rrs1;
    end
    if (reset) begin // @[playground/src/noop/forwading.scala 30:30]
      rs1_d_r <= 64'h0; // @[playground/src/noop/forwading.scala 30:30]
    end else if (hs_in | state) begin // @[playground/src/noop/forwading.scala 170:37]
      if (rs1_valid & cur_rrs1) begin // @[playground/src/noop/forwading.scala 171:36]
        if (cur_rrs1) begin // @[playground/src/noop/forwading.scala 63:19]
          rs1_d_r <= _GEN_34;
        end else begin
          rs1_d_r <= 64'h0; // @[playground/src/noop/forwading.scala 57:62]
        end
      end else begin
        rs1_d_r <= _GEN_93;
      end
    end else begin
      rs1_d_r <= _GEN_93;
    end
    if (reset) begin // @[playground/src/noop/forwading.scala 31:30]
      rs2_r <= 12'h0; // @[playground/src/noop/forwading.scala 31:30]
    end else if (hs_in) begin // @[playground/src/noop/forwading.scala 61:26]
      rs2_r <= io_id2df_rs2;
    end
    if (reset) begin // @[playground/src/noop/forwading.scala 32:30]
      rrs2_r <= 1'h0; // @[playground/src/noop/forwading.scala 32:30]
    end else if (hs_in | state) begin // @[playground/src/noop/forwading.scala 170:37]
      if (rs2_valid & cur_rrs2) begin // @[playground/src/noop/forwading.scala 175:36]
        rrs2_r <= 1'h0; // @[playground/src/noop/forwading.scala 176:21]
      end else begin
        rrs2_r <= cur_rrs2;
      end
    end else begin
      rrs2_r <= cur_rrs2;
    end
    if (reset) begin // @[playground/src/noop/forwading.scala 33:30]
      rs2_d_r <= 64'h0; // @[playground/src/noop/forwading.scala 33:30]
    end else if (hs_in | state) begin // @[playground/src/noop/forwading.scala 170:37]
      if (rs2_valid & cur_rrs2) begin // @[playground/src/noop/forwading.scala 175:36]
        if (cur_rrs2) begin // @[playground/src/noop/forwading.scala 106:19]
          rs2_d_r <= _GEN_73;
        end else begin
          rs2_d_r <= 64'h0; // @[playground/src/noop/forwading.scala 58:62]
        end
      end else begin
        rs2_d_r <= _GEN_96;
      end
    end else begin
      rs2_d_r <= _GEN_96;
    end
    if (reset) begin // @[playground/src/noop/forwading.scala 34:30]
      dst_r <= 5'h0; // @[playground/src/noop/forwading.scala 34:30]
    end else if (hs_in) begin // @[playground/src/noop/forwading.scala 150:16]
      dst_r <= io_id2df_dst; // @[playground/src/noop/forwading.scala 161:21]
    end
    if (reset) begin // @[playground/src/noop/forwading.scala 35:30]
      dst_d_r <= 64'h0; // @[playground/src/noop/forwading.scala 35:30]
    end else if (hs_in) begin // @[playground/src/noop/forwading.scala 150:16]
      dst_d_r <= io_id2df_dst_d; // @[playground/src/noop/forwading.scala 162:21]
    end
    if (reset) begin // @[playground/src/noop/forwading.scala 36:30]
      jmp_type_r <= 2'h0; // @[playground/src/noop/forwading.scala 36:30]
    end else if (hs_in) begin // @[playground/src/noop/forwading.scala 150:16]
      jmp_type_r <= io_id2df_jmp_type; // @[playground/src/noop/forwading.scala 163:21]
    end
    if (reset) begin // @[playground/src/noop/forwading.scala 37:30]
      special_r <= 2'h0; // @[playground/src/noop/forwading.scala 37:30]
    end else if (hs_in) begin // @[playground/src/noop/forwading.scala 150:16]
      special_r <= io_id2df_special; // @[playground/src/noop/forwading.scala 164:21]
    end
    if (reset) begin // @[playground/src/noop/forwading.scala 38:30]
      indi_r <= 2'h0; // @[playground/src/noop/forwading.scala 38:30]
    end else if (hs_in) begin // @[playground/src/noop/forwading.scala 150:16]
      indi_r <= io_id2df_indi; // @[playground/src/noop/forwading.scala 165:21]
    end
    if (reset) begin // @[playground/src/noop/forwading.scala 39:30]
      swap_r <= 6'h0; // @[playground/src/noop/forwading.scala 39:30]
    end else if (hs_in) begin // @[playground/src/noop/forwading.scala 150:16]
      swap_r <= io_id2df_swap; // @[playground/src/noop/forwading.scala 166:21]
    end
    if (reset) begin // @[playground/src/noop/forwading.scala 40:30]
      recov_r <= 1'h0; // @[playground/src/noop/forwading.scala 40:30]
    end else if (hs_in) begin // @[playground/src/noop/forwading.scala 150:16]
      recov_r <= io_id2df_recov; // @[playground/src/noop/forwading.scala 167:21]
    end
    if (reset) begin // @[playground/src/noop/forwading.scala 41:30]
      valid_r <= 1'h0; // @[playground/src/noop/forwading.scala 41:30]
    end else begin
      valid_r <= _GEN_129;
    end
    if (reset) begin // @[playground/src/noop/forwading.scala 43:30]
      pre_dst <= 5'h0; // @[playground/src/noop/forwading.scala 43:30]
    end else if (hs_in) begin // @[playground/src/noop/forwading.scala 181:16]
      pre_dst <= io_id2df_dst; // @[playground/src/noop/forwading.scala 182:17]
    end
    if (reset) begin // @[playground/src/noop/forwading.scala 44:30]
      pre_wr <= 1'h0; // @[playground/src/noop/forwading.scala 44:30]
    end else if (hs_in) begin // @[playground/src/noop/forwading.scala 181:16]
      pre_wr <= io_id2df_ctrl_writeRegEn; // @[playground/src/noop/forwading.scala 183:17]
    end else if (hs_out) begin // @[playground/src/noop/forwading.scala 184:23]
      pre_wr <= 1'h0; // @[playground/src/noop/forwading.scala 185:17]
    end
    if (reset) begin // @[playground/src/noop/forwading.scala 47:24]
      state <= 1'h0; // @[playground/src/noop/forwading.scala 47:24]
    end else begin
      state <= _GEN_128;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  inst_r = _RAND_0[31:0];
  _RAND_1 = {2{`RANDOM}};
  pc_r = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  excep_r_cause = _RAND_2[63:0];
  _RAND_3 = {2{`RANDOM}};
  excep_r_tval = _RAND_3[63:0];
  _RAND_4 = {1{`RANDOM}};
  excep_r_en = _RAND_4[0:0];
  _RAND_5 = {2{`RANDOM}};
  excep_r_pc = _RAND_5[63:0];
  _RAND_6 = {1{`RANDOM}};
  excep_r_etype = _RAND_6[1:0];
  _RAND_7 = {1{`RANDOM}};
  ctrl_r_aluOp = _RAND_7[4:0];
  _RAND_8 = {1{`RANDOM}};
  ctrl_r_aluWidth = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  ctrl_r_dcMode = _RAND_9[4:0];
  _RAND_10 = {1{`RANDOM}};
  ctrl_r_writeRegEn = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  ctrl_r_writeCSREn = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  ctrl_r_brType = _RAND_12[2:0];
  _RAND_13 = {1{`RANDOM}};
  rs1_r = _RAND_13[4:0];
  _RAND_14 = {1{`RANDOM}};
  rrs1_r = _RAND_14[0:0];
  _RAND_15 = {2{`RANDOM}};
  rs1_d_r = _RAND_15[63:0];
  _RAND_16 = {1{`RANDOM}};
  rs2_r = _RAND_16[11:0];
  _RAND_17 = {1{`RANDOM}};
  rrs2_r = _RAND_17[0:0];
  _RAND_18 = {2{`RANDOM}};
  rs2_d_r = _RAND_18[63:0];
  _RAND_19 = {1{`RANDOM}};
  dst_r = _RAND_19[4:0];
  _RAND_20 = {2{`RANDOM}};
  dst_d_r = _RAND_20[63:0];
  _RAND_21 = {1{`RANDOM}};
  jmp_type_r = _RAND_21[1:0];
  _RAND_22 = {1{`RANDOM}};
  special_r = _RAND_22[1:0];
  _RAND_23 = {1{`RANDOM}};
  indi_r = _RAND_23[1:0];
  _RAND_24 = {1{`RANDOM}};
  swap_r = _RAND_24[5:0];
  _RAND_25 = {1{`RANDOM}};
  recov_r = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  valid_r = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  pre_dst = _RAND_27[4:0];
  _RAND_28 = {1{`RANDOM}};
  pre_wr = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  state = _RAND_29[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ReadRegs(
  input         clock,
  input         reset,
  input  [31:0] io_df2rr_inst, // @[playground/src/noop/readregs.scala 10:16]
  input  [63:0] io_df2rr_pc, // @[playground/src/noop/readregs.scala 10:16]
  input  [63:0] io_df2rr_excep_cause, // @[playground/src/noop/readregs.scala 10:16]
  input  [63:0] io_df2rr_excep_tval, // @[playground/src/noop/readregs.scala 10:16]
  input         io_df2rr_excep_en, // @[playground/src/noop/readregs.scala 10:16]
  input  [63:0] io_df2rr_excep_pc, // @[playground/src/noop/readregs.scala 10:16]
  input  [1:0]  io_df2rr_excep_etype, // @[playground/src/noop/readregs.scala 10:16]
  input  [4:0]  io_df2rr_ctrl_aluOp, // @[playground/src/noop/readregs.scala 10:16]
  input         io_df2rr_ctrl_aluWidth, // @[playground/src/noop/readregs.scala 10:16]
  input  [4:0]  io_df2rr_ctrl_dcMode, // @[playground/src/noop/readregs.scala 10:16]
  input         io_df2rr_ctrl_writeRegEn, // @[playground/src/noop/readregs.scala 10:16]
  input         io_df2rr_ctrl_writeCSREn, // @[playground/src/noop/readregs.scala 10:16]
  input  [2:0]  io_df2rr_ctrl_brType, // @[playground/src/noop/readregs.scala 10:16]
  input  [4:0]  io_df2rr_rs1, // @[playground/src/noop/readregs.scala 10:16]
  input         io_df2rr_rrs1, // @[playground/src/noop/readregs.scala 10:16]
  input  [63:0] io_df2rr_rs1_d, // @[playground/src/noop/readregs.scala 10:16]
  input  [11:0] io_df2rr_rs2, // @[playground/src/noop/readregs.scala 10:16]
  input         io_df2rr_rrs2, // @[playground/src/noop/readregs.scala 10:16]
  input  [63:0] io_df2rr_rs2_d, // @[playground/src/noop/readregs.scala 10:16]
  input  [4:0]  io_df2rr_dst, // @[playground/src/noop/readregs.scala 10:16]
  input  [63:0] io_df2rr_dst_d, // @[playground/src/noop/readregs.scala 10:16]
  input  [1:0]  io_df2rr_jmp_type, // @[playground/src/noop/readregs.scala 10:16]
  input  [1:0]  io_df2rr_special, // @[playground/src/noop/readregs.scala 10:16]
  input  [5:0]  io_df2rr_swap, // @[playground/src/noop/readregs.scala 10:16]
  input  [1:0]  io_df2rr_indi, // @[playground/src/noop/readregs.scala 10:16]
  output        io_df2rr_drop, // @[playground/src/noop/readregs.scala 10:16]
  output        io_df2rr_stall, // @[playground/src/noop/readregs.scala 10:16]
  input         io_df2rr_recov, // @[playground/src/noop/readregs.scala 10:16]
  input         io_df2rr_valid, // @[playground/src/noop/readregs.scala 10:16]
  output        io_df2rr_ready, // @[playground/src/noop/readregs.scala 10:16]
  output [31:0] io_rr2ex_inst, // @[playground/src/noop/readregs.scala 10:16]
  output [63:0] io_rr2ex_pc, // @[playground/src/noop/readregs.scala 10:16]
  output [63:0] io_rr2ex_excep_cause, // @[playground/src/noop/readregs.scala 10:16]
  output [63:0] io_rr2ex_excep_tval, // @[playground/src/noop/readregs.scala 10:16]
  output        io_rr2ex_excep_en, // @[playground/src/noop/readregs.scala 10:16]
  output [63:0] io_rr2ex_excep_pc, // @[playground/src/noop/readregs.scala 10:16]
  output [1:0]  io_rr2ex_excep_etype, // @[playground/src/noop/readregs.scala 10:16]
  output [4:0]  io_rr2ex_ctrl_aluOp, // @[playground/src/noop/readregs.scala 10:16]
  output        io_rr2ex_ctrl_aluWidth, // @[playground/src/noop/readregs.scala 10:16]
  output [4:0]  io_rr2ex_ctrl_dcMode, // @[playground/src/noop/readregs.scala 10:16]
  output        io_rr2ex_ctrl_writeRegEn, // @[playground/src/noop/readregs.scala 10:16]
  output        io_rr2ex_ctrl_writeCSREn, // @[playground/src/noop/readregs.scala 10:16]
  output [2:0]  io_rr2ex_ctrl_brType, // @[playground/src/noop/readregs.scala 10:16]
  output [63:0] io_rr2ex_rs1_d, // @[playground/src/noop/readregs.scala 10:16]
  output [11:0] io_rr2ex_rs2, // @[playground/src/noop/readregs.scala 10:16]
  output [63:0] io_rr2ex_rs2_d, // @[playground/src/noop/readregs.scala 10:16]
  output [4:0]  io_rr2ex_dst, // @[playground/src/noop/readregs.scala 10:16]
  output [63:0] io_rr2ex_dst_d, // @[playground/src/noop/readregs.scala 10:16]
  output [11:0] io_rr2ex_rcsr_id, // @[playground/src/noop/readregs.scala 10:16]
  output [1:0]  io_rr2ex_jmp_type, // @[playground/src/noop/readregs.scala 10:16]
  output [1:0]  io_rr2ex_special, // @[playground/src/noop/readregs.scala 10:16]
  output [1:0]  io_rr2ex_indi, // @[playground/src/noop/readregs.scala 10:16]
  input         io_rr2ex_drop, // @[playground/src/noop/readregs.scala 10:16]
  input         io_rr2ex_stall, // @[playground/src/noop/readregs.scala 10:16]
  output        io_rr2ex_recov, // @[playground/src/noop/readregs.scala 10:16]
  output        io_rr2ex_valid, // @[playground/src/noop/readregs.scala 10:16]
  input         io_rr2ex_ready, // @[playground/src/noop/readregs.scala 10:16]
  output [4:0]  io_rs1Read_id, // @[playground/src/noop/readregs.scala 10:16]
  input  [63:0] io_rs1Read_data, // @[playground/src/noop/readregs.scala 10:16]
  output [4:0]  io_rs2Read_id, // @[playground/src/noop/readregs.scala 10:16]
  input  [63:0] io_rs2Read_data, // @[playground/src/noop/readregs.scala 10:16]
  output [11:0] io_csrRead_id, // @[playground/src/noop/readregs.scala 10:16]
  input  [63:0] io_csrRead_data, // @[playground/src/noop/readregs.scala 10:16]
  input         io_csrRead_is_err, // @[playground/src/noop/readregs.scala 10:16]
  output [4:0]  io_d_rr_id, // @[playground/src/noop/readregs.scala 10:16]
  output [63:0] io_d_rr_data, // @[playground/src/noop/readregs.scala 10:16]
  output [1:0]  io_d_rr_state // @[playground/src/noop/readregs.scala 10:16]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [63:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [63:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [63:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
`endif // RANDOMIZE_REG_INIT
  reg  drop_r; // @[playground/src/noop/readregs.scala 18:30]
  reg  stall_r; // @[playground/src/noop/readregs.scala 20:30]
  reg  recov_r; // @[playground/src/noop/readregs.scala 22:30]
  wire  drop_in = io_rr2ex_drop | drop_r; // @[playground/src/noop/readregs.scala 26:37]
  wire  _io_df2rr_stall_T = ~io_rr2ex_drop; // @[playground/src/noop/readregs.scala 28:36]
  reg [31:0] inst_r; // @[playground/src/noop/readregs.scala 29:30]
  reg [63:0] pc_r; // @[playground/src/noop/readregs.scala 30:30]
  reg [63:0] excep_r_cause; // @[playground/src/noop/readregs.scala 31:30]
  reg [63:0] excep_r_tval; // @[playground/src/noop/readregs.scala 31:30]
  reg  excep_r_en; // @[playground/src/noop/readregs.scala 31:30]
  reg [63:0] excep_r_pc; // @[playground/src/noop/readregs.scala 31:30]
  reg [1:0] excep_r_etype; // @[playground/src/noop/readregs.scala 31:30]
  reg [4:0] ctrl_r_aluOp; // @[playground/src/noop/readregs.scala 32:30]
  reg  ctrl_r_aluWidth; // @[playground/src/noop/readregs.scala 32:30]
  reg [4:0] ctrl_r_dcMode; // @[playground/src/noop/readregs.scala 32:30]
  reg  ctrl_r_writeRegEn; // @[playground/src/noop/readregs.scala 32:30]
  reg  ctrl_r_writeCSREn; // @[playground/src/noop/readregs.scala 32:30]
  reg [2:0] ctrl_r_brType; // @[playground/src/noop/readregs.scala 32:30]
  reg [63:0] rs1_d_r; // @[playground/src/noop/readregs.scala 34:30]
  reg [11:0] rs2_r; // @[playground/src/noop/readregs.scala 35:30]
  reg [63:0] rs2_d_r; // @[playground/src/noop/readregs.scala 36:30]
  reg [4:0] dst_r; // @[playground/src/noop/readregs.scala 37:30]
  reg [63:0] dst_d_r; // @[playground/src/noop/readregs.scala 38:30]
  reg [11:0] rcsr_id_r; // @[playground/src/noop/readregs.scala 39:30]
  reg [1:0] jmp_type_r; // @[playground/src/noop/readregs.scala 40:30]
  reg [1:0] special_r; // @[playground/src/noop/readregs.scala 41:30]
  reg [1:0] indi_r; // @[playground/src/noop/readregs.scala 42:30]
  reg  valid_r; // @[playground/src/noop/readregs.scala 44:30]
  wire  hs_in = io_df2rr_ready & io_df2rr_valid; // @[playground/src/noop/readregs.scala 46:34]
  wire  hs_out = io_rr2ex_ready & io_rr2ex_valid; // @[playground/src/noop/readregs.scala 47:34]
  wire [63:0] rs1_bef = io_df2rr_rrs1 ? io_rs1Read_data : io_df2rr_rs1_d; // @[playground/src/noop/readregs.scala 52:22]
  wire [63:0] _rs2_bef_T_2 = io_df2rr_rrs2 ? io_rs2Read_data : io_df2rr_rs2_d; // @[playground/src/noop/readregs.scala 53:98]
  wire [63:0] rs2_bef = io_df2rr_ctrl_writeCSREn | io_df2rr_excep_en ? io_csrRead_data : _rs2_bef_T_2; // @[playground/src/noop/readregs.scala 53:22]
  wire [63:0] _rs1_d_r_T_2 = 2'h1 == io_df2rr_swap[5:4] ? rs1_bef : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 81:58]
  wire [63:0] _rs2_d_r_T_2 = 2'h1 == io_df2rr_swap[3:2] ? rs1_bef : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 81:58]
  wire [63:0] _dst_d_r_T_2 = 2'h1 == io_df2rr_swap[1:0] ? rs1_bef : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 81:58]
  wire  _T = io_df2rr_ctrl_writeCSREn & io_csrRead_is_err; // @[playground/src/noop/readregs.scala 78:39]
  wire  _GEN_2 = io_df2rr_ctrl_writeCSREn & io_csrRead_is_err | io_df2rr_excep_en; // @[playground/src/noop/readregs.scala 65:21 78:60 81:29]
  wire  _GEN_6 = io_df2rr_ctrl_writeCSREn & io_csrRead_is_err | io_df2rr_recov; // @[playground/src/noop/readregs.scala 24:57 77:21 78:60]
  wire  _GEN_39 = hs_in & _T; // @[playground/src/noop/readregs.scala 62:16 19:21]
  wire  _GEN_41 = valid_r & ~hs_out ? 1'h0 : io_df2rr_valid; // @[playground/src/noop/readregs.scala 90:20 92:33]
  wire  _GEN_43 = hs_out ? 1'h0 : valid_r; // @[playground/src/noop/readregs.scala 100:27 101:21 44:30]
  wire  _GEN_44 = hs_in | _GEN_43; // @[playground/src/noop/readregs.scala 98:20 99:21]
  wire  _GEN_45 = _io_df2rr_stall_T & _GEN_44; // @[playground/src/noop/readregs.scala 104:17 97:25]
  assign io_df2rr_drop = io_rr2ex_drop | drop_r; // @[playground/src/noop/readregs.scala 26:37]
  assign io_df2rr_stall = stall_r & ~io_rr2ex_drop | io_rr2ex_stall; // @[playground/src/noop/readregs.scala 28:52]
  assign io_df2rr_ready = ~drop_in & _GEN_41; // @[playground/src/noop/readregs.scala 91:19 90:20]
  assign io_rr2ex_inst = inst_r; // @[playground/src/noop/readregs.scala 106:25]
  assign io_rr2ex_pc = pc_r; // @[playground/src/noop/readregs.scala 107:25]
  assign io_rr2ex_excep_cause = excep_r_cause; // @[playground/src/noop/readregs.scala 108:25]
  assign io_rr2ex_excep_tval = excep_r_tval; // @[playground/src/noop/readregs.scala 108:25]
  assign io_rr2ex_excep_en = excep_r_en; // @[playground/src/noop/readregs.scala 108:25]
  assign io_rr2ex_excep_pc = excep_r_pc; // @[playground/src/noop/readregs.scala 108:25]
  assign io_rr2ex_excep_etype = excep_r_etype; // @[playground/src/noop/readregs.scala 108:25]
  assign io_rr2ex_ctrl_aluOp = ctrl_r_aluOp; // @[playground/src/noop/readregs.scala 109:25]
  assign io_rr2ex_ctrl_aluWidth = ctrl_r_aluWidth; // @[playground/src/noop/readregs.scala 109:25]
  assign io_rr2ex_ctrl_dcMode = ctrl_r_dcMode; // @[playground/src/noop/readregs.scala 109:25]
  assign io_rr2ex_ctrl_writeRegEn = ctrl_r_writeRegEn; // @[playground/src/noop/readregs.scala 109:25]
  assign io_rr2ex_ctrl_writeCSREn = ctrl_r_writeCSREn; // @[playground/src/noop/readregs.scala 109:25]
  assign io_rr2ex_ctrl_brType = ctrl_r_brType; // @[playground/src/noop/readregs.scala 109:25]
  assign io_rr2ex_rs1_d = rs1_d_r; // @[playground/src/noop/readregs.scala 111:25]
  assign io_rr2ex_rs2 = rs2_r; // @[playground/src/noop/readregs.scala 112:25]
  assign io_rr2ex_rs2_d = rs2_d_r; // @[playground/src/noop/readregs.scala 113:25]
  assign io_rr2ex_dst = dst_r; // @[playground/src/noop/readregs.scala 114:25]
  assign io_rr2ex_dst_d = dst_d_r; // @[playground/src/noop/readregs.scala 115:25]
  assign io_rr2ex_rcsr_id = rcsr_id_r; // @[playground/src/noop/readregs.scala 116:25]
  assign io_rr2ex_jmp_type = jmp_type_r; // @[playground/src/noop/readregs.scala 117:25]
  assign io_rr2ex_special = special_r; // @[playground/src/noop/readregs.scala 118:25]
  assign io_rr2ex_indi = indi_r; // @[playground/src/noop/readregs.scala 119:25]
  assign io_rr2ex_recov = recov_r; // @[playground/src/noop/readregs.scala 120:25]
  assign io_rr2ex_valid = valid_r; // @[playground/src/noop/readregs.scala 121:25]
  assign io_rs1Read_id = io_df2rr_rs1; // @[playground/src/noop/readregs.scala 49:19]
  assign io_rs2Read_id = io_df2rr_rs2[4:0]; // @[playground/src/noop/readregs.scala 50:34]
  assign io_csrRead_id = io_df2rr_rs2; // @[playground/src/noop/readregs.scala 51:19]
  assign io_d_rr_id = dst_r; // @[playground/src/noop/readregs.scala 123:21]
  assign io_d_rr_data = dst_d_r; // @[playground/src/noop/readregs.scala 124:21]
  assign io_d_rr_state = valid_r ? 2'h2 : 2'h0; // @[playground/src/noop/readregs.scala 125:27]
  always @(posedge clock) begin
    if (reset) begin // @[playground/src/noop/readregs.scala 18:30]
      drop_r <= 1'h0; // @[playground/src/noop/readregs.scala 18:30]
    end else begin
      drop_r <= _GEN_39;
    end
    if (reset) begin // @[playground/src/noop/readregs.scala 20:30]
      stall_r <= 1'h0; // @[playground/src/noop/readregs.scala 20:30]
    end else begin
      stall_r <= _GEN_39;
    end
    if (reset) begin // @[playground/src/noop/readregs.scala 22:30]
      recov_r <= 1'h0; // @[playground/src/noop/readregs.scala 22:30]
    end else if (hs_in) begin // @[playground/src/noop/readregs.scala 62:16]
      recov_r <= _GEN_6;
    end
    if (reset) begin // @[playground/src/noop/readregs.scala 29:30]
      inst_r <= 32'h0; // @[playground/src/noop/readregs.scala 29:30]
    end else if (hs_in) begin // @[playground/src/noop/readregs.scala 62:16]
      inst_r <= io_df2rr_inst; // @[playground/src/noop/readregs.scala 63:21]
    end
    if (reset) begin // @[playground/src/noop/readregs.scala 30:30]
      pc_r <= 64'h0; // @[playground/src/noop/readregs.scala 30:30]
    end else if (hs_in) begin // @[playground/src/noop/readregs.scala 62:16]
      pc_r <= io_df2rr_pc; // @[playground/src/noop/readregs.scala 64:21]
    end
    if (reset) begin // @[playground/src/noop/readregs.scala 31:30]
      excep_r_cause <= 64'h0; // @[playground/src/noop/readregs.scala 31:30]
    end else if (hs_in) begin // @[playground/src/noop/readregs.scala 62:16]
      if (io_df2rr_ctrl_writeCSREn & io_csrRead_is_err) begin // @[playground/src/noop/readregs.scala 78:60]
        excep_r_cause <= 64'h2; // @[playground/src/noop/readregs.scala 79:29]
      end else begin
        excep_r_cause <= io_df2rr_excep_cause; // @[playground/src/noop/readregs.scala 65:21]
      end
    end
    if (reset) begin // @[playground/src/noop/readregs.scala 31:30]
      excep_r_tval <= 64'h0; // @[playground/src/noop/readregs.scala 31:30]
    end else if (hs_in) begin // @[playground/src/noop/readregs.scala 62:16]
      if (io_df2rr_ctrl_writeCSREn & io_csrRead_is_err) begin // @[playground/src/noop/readregs.scala 78:60]
        excep_r_tval <= {{32'd0}, io_df2rr_inst}; // @[playground/src/noop/readregs.scala 80:29]
      end else begin
        excep_r_tval <= io_df2rr_excep_tval; // @[playground/src/noop/readregs.scala 65:21]
      end
    end
    if (reset) begin // @[playground/src/noop/readregs.scala 31:30]
      excep_r_en <= 1'h0; // @[playground/src/noop/readregs.scala 31:30]
    end else if (hs_in) begin // @[playground/src/noop/readregs.scala 62:16]
      excep_r_en <= _GEN_2;
    end
    if (reset) begin // @[playground/src/noop/readregs.scala 31:30]
      excep_r_pc <= 64'h0; // @[playground/src/noop/readregs.scala 31:30]
    end else if (hs_in) begin // @[playground/src/noop/readregs.scala 62:16]
      if (io_df2rr_ctrl_writeCSREn & io_csrRead_is_err) begin // @[playground/src/noop/readregs.scala 78:60]
        excep_r_pc <= io_df2rr_pc; // @[playground/src/noop/readregs.scala 82:29]
      end else begin
        excep_r_pc <= io_df2rr_excep_pc; // @[playground/src/noop/readregs.scala 65:21]
      end
    end
    if (reset) begin // @[playground/src/noop/readregs.scala 31:30]
      excep_r_etype <= 2'h0; // @[playground/src/noop/readregs.scala 31:30]
    end else if (hs_in) begin // @[playground/src/noop/readregs.scala 62:16]
      if (io_df2rr_ctrl_writeCSREn & io_csrRead_is_err) begin // @[playground/src/noop/readregs.scala 78:60]
        excep_r_etype <= 2'h0; // @[playground/src/noop/readregs.scala 83:29]
      end else begin
        excep_r_etype <= io_df2rr_excep_etype; // @[playground/src/noop/readregs.scala 65:21]
      end
    end
    if (reset) begin // @[playground/src/noop/readregs.scala 32:30]
      ctrl_r_aluOp <= 5'h0; // @[playground/src/noop/readregs.scala 32:30]
    end else if (hs_in) begin // @[playground/src/noop/readregs.scala 62:16]
      if (io_df2rr_ctrl_writeCSREn & io_csrRead_is_err) begin // @[playground/src/noop/readregs.scala 78:60]
        ctrl_r_aluOp <= 5'h0; // @[playground/src/noop/readregs.scala 85:25]
      end else begin
        ctrl_r_aluOp <= io_df2rr_ctrl_aluOp; // @[playground/src/noop/readregs.scala 66:21]
      end
    end
    if (reset) begin // @[playground/src/noop/readregs.scala 32:30]
      ctrl_r_aluWidth <= 1'h0; // @[playground/src/noop/readregs.scala 32:30]
    end else if (hs_in) begin // @[playground/src/noop/readregs.scala 62:16]
      if (io_df2rr_ctrl_writeCSREn & io_csrRead_is_err) begin // @[playground/src/noop/readregs.scala 78:60]
        ctrl_r_aluWidth <= 1'h0; // @[playground/src/noop/readregs.scala 85:25]
      end else begin
        ctrl_r_aluWidth <= io_df2rr_ctrl_aluWidth; // @[playground/src/noop/readregs.scala 66:21]
      end
    end
    if (reset) begin // @[playground/src/noop/readregs.scala 32:30]
      ctrl_r_dcMode <= 5'h0; // @[playground/src/noop/readregs.scala 32:30]
    end else if (hs_in) begin // @[playground/src/noop/readregs.scala 62:16]
      if (io_df2rr_ctrl_writeCSREn & io_csrRead_is_err) begin // @[playground/src/noop/readregs.scala 78:60]
        ctrl_r_dcMode <= 5'h0; // @[playground/src/noop/readregs.scala 85:25]
      end else begin
        ctrl_r_dcMode <= io_df2rr_ctrl_dcMode; // @[playground/src/noop/readregs.scala 66:21]
      end
    end
    if (reset) begin // @[playground/src/noop/readregs.scala 32:30]
      ctrl_r_writeRegEn <= 1'h0; // @[playground/src/noop/readregs.scala 32:30]
    end else if (hs_in) begin // @[playground/src/noop/readregs.scala 62:16]
      if (io_df2rr_ctrl_writeCSREn & io_csrRead_is_err) begin // @[playground/src/noop/readregs.scala 78:60]
        ctrl_r_writeRegEn <= 1'h0; // @[playground/src/noop/readregs.scala 85:25]
      end else begin
        ctrl_r_writeRegEn <= io_df2rr_ctrl_writeRegEn; // @[playground/src/noop/readregs.scala 66:21]
      end
    end
    if (reset) begin // @[playground/src/noop/readregs.scala 32:30]
      ctrl_r_writeCSREn <= 1'h0; // @[playground/src/noop/readregs.scala 32:30]
    end else if (hs_in) begin // @[playground/src/noop/readregs.scala 62:16]
      if (io_df2rr_ctrl_writeCSREn & io_csrRead_is_err) begin // @[playground/src/noop/readregs.scala 78:60]
        ctrl_r_writeCSREn <= 1'h0; // @[playground/src/noop/readregs.scala 85:25]
      end else begin
        ctrl_r_writeCSREn <= io_df2rr_ctrl_writeCSREn; // @[playground/src/noop/readregs.scala 66:21]
      end
    end
    if (reset) begin // @[playground/src/noop/readregs.scala 32:30]
      ctrl_r_brType <= 3'h0; // @[playground/src/noop/readregs.scala 32:30]
    end else if (hs_in) begin // @[playground/src/noop/readregs.scala 62:16]
      if (io_df2rr_ctrl_writeCSREn & io_csrRead_is_err) begin // @[playground/src/noop/readregs.scala 78:60]
        ctrl_r_brType <= 3'h0; // @[playground/src/noop/readregs.scala 85:25]
      end else begin
        ctrl_r_brType <= io_df2rr_ctrl_brType; // @[playground/src/noop/readregs.scala 66:21]
      end
    end
    if (reset) begin // @[playground/src/noop/readregs.scala 34:30]
      rs1_d_r <= 64'h0; // @[playground/src/noop/readregs.scala 34:30]
    end else if (hs_in) begin // @[playground/src/noop/readregs.scala 62:16]
      if (2'h3 == io_df2rr_swap[5:4]) begin // @[src/main/scala/chisel3/util/Mux.scala 81:58]
        rs1_d_r <= io_df2rr_dst_d;
      end else if (2'h2 == io_df2rr_swap[5:4]) begin // @[src/main/scala/chisel3/util/Mux.scala 81:58]
        rs1_d_r <= rs2_bef;
      end else begin
        rs1_d_r <= _rs1_d_r_T_2;
      end
    end
    if (reset) begin // @[playground/src/noop/readregs.scala 35:30]
      rs2_r <= 12'h0; // @[playground/src/noop/readregs.scala 35:30]
    end else if (hs_in) begin // @[playground/src/noop/readregs.scala 62:16]
      rs2_r <= io_df2rr_rs2; // @[playground/src/noop/readregs.scala 69:21]
    end
    if (reset) begin // @[playground/src/noop/readregs.scala 36:30]
      rs2_d_r <= 64'h0; // @[playground/src/noop/readregs.scala 36:30]
    end else if (hs_in) begin // @[playground/src/noop/readregs.scala 62:16]
      if (2'h3 == io_df2rr_swap[3:2]) begin // @[src/main/scala/chisel3/util/Mux.scala 81:58]
        rs2_d_r <= io_df2rr_dst_d;
      end else if (2'h2 == io_df2rr_swap[3:2]) begin // @[src/main/scala/chisel3/util/Mux.scala 81:58]
        rs2_d_r <= rs2_bef;
      end else begin
        rs2_d_r <= _rs2_d_r_T_2;
      end
    end
    if (reset) begin // @[playground/src/noop/readregs.scala 37:30]
      dst_r <= 5'h0; // @[playground/src/noop/readregs.scala 37:30]
    end else if (hs_in) begin // @[playground/src/noop/readregs.scala 62:16]
      dst_r <= io_df2rr_dst; // @[playground/src/noop/readregs.scala 71:21]
    end
    if (reset) begin // @[playground/src/noop/readregs.scala 38:30]
      dst_d_r <= 64'h0; // @[playground/src/noop/readregs.scala 38:30]
    end else if (hs_in) begin // @[playground/src/noop/readregs.scala 62:16]
      if (2'h3 == io_df2rr_swap[1:0]) begin // @[src/main/scala/chisel3/util/Mux.scala 81:58]
        dst_d_r <= io_df2rr_dst_d;
      end else if (2'h2 == io_df2rr_swap[1:0]) begin // @[src/main/scala/chisel3/util/Mux.scala 81:58]
        dst_d_r <= rs2_bef;
      end else begin
        dst_d_r <= _dst_d_r_T_2;
      end
    end
    if (reset) begin // @[playground/src/noop/readregs.scala 39:30]
      rcsr_id_r <= 12'h0; // @[playground/src/noop/readregs.scala 39:30]
    end else if (hs_in) begin // @[playground/src/noop/readregs.scala 62:16]
      if (io_df2rr_ctrl_writeCSREn) begin // @[playground/src/noop/readregs.scala 73:27]
        rcsr_id_r <= io_df2rr_rs2;
      end else begin
        rcsr_id_r <= 12'h0;
      end
    end
    if (reset) begin // @[playground/src/noop/readregs.scala 40:30]
      jmp_type_r <= 2'h0; // @[playground/src/noop/readregs.scala 40:30]
    end else if (hs_in) begin // @[playground/src/noop/readregs.scala 62:16]
      if (io_df2rr_ctrl_writeCSREn & io_csrRead_is_err) begin // @[playground/src/noop/readregs.scala 78:60]
        jmp_type_r <= 2'h0; // @[playground/src/noop/readregs.scala 86:25]
      end else begin
        jmp_type_r <= io_df2rr_jmp_type; // @[playground/src/noop/readregs.scala 74:21]
      end
    end
    if (reset) begin // @[playground/src/noop/readregs.scala 41:30]
      special_r <= 2'h0; // @[playground/src/noop/readregs.scala 41:30]
    end else if (hs_in) begin // @[playground/src/noop/readregs.scala 62:16]
      if (io_df2rr_ctrl_writeCSREn & io_csrRead_is_err) begin // @[playground/src/noop/readregs.scala 78:60]
        special_r <= 2'h0; // @[playground/src/noop/readregs.scala 87:25]
      end else begin
        special_r <= io_df2rr_special; // @[playground/src/noop/readregs.scala 75:21]
      end
    end
    if (reset) begin // @[playground/src/noop/readregs.scala 42:30]
      indi_r <= 2'h0; // @[playground/src/noop/readregs.scala 42:30]
    end else if (hs_in) begin // @[playground/src/noop/readregs.scala 62:16]
      indi_r <= io_df2rr_indi; // @[playground/src/noop/readregs.scala 76:21]
    end
    if (reset) begin // @[playground/src/noop/readregs.scala 44:30]
      valid_r <= 1'h0; // @[playground/src/noop/readregs.scala 44:30]
    end else begin
      valid_r <= _GEN_45;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  drop_r = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  stall_r = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  recov_r = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  inst_r = _RAND_3[31:0];
  _RAND_4 = {2{`RANDOM}};
  pc_r = _RAND_4[63:0];
  _RAND_5 = {2{`RANDOM}};
  excep_r_cause = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  excep_r_tval = _RAND_6[63:0];
  _RAND_7 = {1{`RANDOM}};
  excep_r_en = _RAND_7[0:0];
  _RAND_8 = {2{`RANDOM}};
  excep_r_pc = _RAND_8[63:0];
  _RAND_9 = {1{`RANDOM}};
  excep_r_etype = _RAND_9[1:0];
  _RAND_10 = {1{`RANDOM}};
  ctrl_r_aluOp = _RAND_10[4:0];
  _RAND_11 = {1{`RANDOM}};
  ctrl_r_aluWidth = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  ctrl_r_dcMode = _RAND_12[4:0];
  _RAND_13 = {1{`RANDOM}};
  ctrl_r_writeRegEn = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  ctrl_r_writeCSREn = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  ctrl_r_brType = _RAND_15[2:0];
  _RAND_16 = {2{`RANDOM}};
  rs1_d_r = _RAND_16[63:0];
  _RAND_17 = {1{`RANDOM}};
  rs2_r = _RAND_17[11:0];
  _RAND_18 = {2{`RANDOM}};
  rs2_d_r = _RAND_18[63:0];
  _RAND_19 = {1{`RANDOM}};
  dst_r = _RAND_19[4:0];
  _RAND_20 = {2{`RANDOM}};
  dst_d_r = _RAND_20[63:0];
  _RAND_21 = {1{`RANDOM}};
  rcsr_id_r = _RAND_21[11:0];
  _RAND_22 = {1{`RANDOM}};
  jmp_type_r = _RAND_22[1:0];
  _RAND_23 = {1{`RANDOM}};
  special_r = _RAND_23[1:0];
  _RAND_24 = {1{`RANDOM}};
  indi_r = _RAND_24[1:0];
  _RAND_25 = {1{`RANDOM}};
  valid_r = _RAND_25[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module MUL(
  input         clock,
  input         reset,
  input  [63:0] io_a, // @[playground/src/noop/muldiv.scala 18:16]
  input  [63:0] io_b, // @[playground/src/noop/muldiv.scala 18:16]
  input  [4:0]  io_aluop, // @[playground/src/noop/muldiv.scala 18:16]
  input         io_en, // @[playground/src/noop/muldiv.scala 18:16]
  output [63:0] io_out, // @[playground/src/noop/muldiv.scala 18:16]
  output        io_valid // @[playground/src/noop/muldiv.scala 18:16]
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
`endif // RANDOMIZE_REG_INIT
  reg [63:0] out_r; // @[playground/src/noop/muldiv.scala 20:30]
  reg [63:0] val1; // @[playground/src/noop/muldiv.scala 21:30]
  reg [63:0] val2; // @[playground/src/noop/muldiv.scala 22:30]
  reg [4:0] aluop_r; // @[playground/src/noop/muldiv.scala 23:33]
  reg  valid_r; // @[playground/src/noop/muldiv.scala 24:30]
  reg [1:0] state; // @[playground/src/noop/muldiv.scala 26:24]
  wire [127:0] _out_r_T = val1 * val2; // @[playground/src/noop/muldiv.scala 42:34]
  wire [127:0] _out_r_T_4 = $signed(val1) * $signed(val2); // @[playground/src/noop/muldiv.scala 43:42]
  wire [64:0] _out_r_T_9 = {1'b0,$signed(val2)}; // @[playground/src/noop/muldiv.scala 45:41]
  wire [128:0] _out_r_T_10 = $signed(val1) * $signed(_out_r_T_9); // @[playground/src/noop/muldiv.scala 45:41]
  wire [127:0] _out_r_T_12 = _out_r_T_10[127:0]; // @[playground/src/noop/muldiv.scala 45:41]
  wire [63:0] _out_r_T_15 = _out_r_T_12[127:64]; // @[playground/src/noop/muldiv.scala 45:65]
  wire [63:0] _out_r_T_17 = 5'hd == aluop_r ? _out_r_T[63:0] : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 81:58]
  wire [63:0] _out_r_T_19 = 5'he == aluop_r ? _out_r_T_4[127:64] : _out_r_T_17; // @[src/main/scala/chisel3/util/Mux.scala 81:58]
  wire [63:0] _out_r_T_21 = 5'hf == aluop_r ? _out_r_T[127:64] : _out_r_T_19; // @[src/main/scala/chisel3/util/Mux.scala 81:58]
  wire  _GEN_5 = 2'h1 == state | valid_r; // @[playground/src/noop/muldiv.scala 30:18 47:21 24:30]
  assign io_out = out_r; // @[playground/src/noop/muldiv.scala 28:12]
  assign io_valid = valid_r; // @[playground/src/noop/muldiv.scala 29:14]
  always @(posedge clock) begin
    if (reset) begin // @[playground/src/noop/muldiv.scala 20:30]
      out_r <= 64'h0; // @[playground/src/noop/muldiv.scala 20:30]
    end else if (!(2'h0 == state)) begin // @[playground/src/noop/muldiv.scala 30:18]
      if (2'h1 == state) begin // @[playground/src/noop/muldiv.scala 30:18]
        if (5'h10 == aluop_r) begin // @[src/main/scala/chisel3/util/Mux.scala 81:58]
          out_r <= _out_r_T_15;
        end else begin
          out_r <= _out_r_T_21;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/muldiv.scala 21:30]
      val1 <= 64'h0; // @[playground/src/noop/muldiv.scala 21:30]
    end else if (2'h0 == state) begin // @[playground/src/noop/muldiv.scala 30:18]
      if (io_en) begin // @[playground/src/noop/muldiv.scala 33:24]
        val1 <= io_a; // @[playground/src/noop/muldiv.scala 35:22]
      end
    end
    if (reset) begin // @[playground/src/noop/muldiv.scala 22:30]
      val2 <= 64'h0; // @[playground/src/noop/muldiv.scala 22:30]
    end else if (2'h0 == state) begin // @[playground/src/noop/muldiv.scala 30:18]
      if (io_en) begin // @[playground/src/noop/muldiv.scala 33:24]
        val2 <= io_b; // @[playground/src/noop/muldiv.scala 36:22]
      end
    end
    if (reset) begin // @[playground/src/noop/muldiv.scala 23:33]
      aluop_r <= 5'h0; // @[playground/src/noop/muldiv.scala 23:33]
    end else if (2'h0 == state) begin // @[playground/src/noop/muldiv.scala 30:18]
      if (io_en) begin // @[playground/src/noop/muldiv.scala 33:24]
        aluop_r <= io_aluop; // @[playground/src/noop/muldiv.scala 37:25]
      end
    end
    if (reset) begin // @[playground/src/noop/muldiv.scala 24:30]
      valid_r <= 1'h0; // @[playground/src/noop/muldiv.scala 24:30]
    end else if (2'h0 == state) begin // @[playground/src/noop/muldiv.scala 30:18]
      valid_r <= 1'h0; // @[playground/src/noop/muldiv.scala 32:21]
    end else begin
      valid_r <= _GEN_5;
    end
    if (reset) begin // @[playground/src/noop/muldiv.scala 26:24]
      state <= 2'h0; // @[playground/src/noop/muldiv.scala 26:24]
    end else if (2'h0 == state) begin // @[playground/src/noop/muldiv.scala 30:18]
      if (io_en) begin // @[playground/src/noop/muldiv.scala 33:24]
        state <= 2'h1; // @[playground/src/noop/muldiv.scala 34:23]
      end
    end else if (2'h1 == state) begin // @[playground/src/noop/muldiv.scala 30:18]
      state <= 2'h0; // @[playground/src/noop/muldiv.scala 48:19]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  out_r = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  val1 = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  val2 = _RAND_2[63:0];
  _RAND_3 = {1{`RANDOM}};
  aluop_r = _RAND_3[4:0];
  _RAND_4 = {1{`RANDOM}};
  valid_r = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  state = _RAND_5[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module DIV(
  input         clock,
  input         reset,
  input         io_alu64, // @[playground/src/noop/muldiv.scala 66:16]
  input  [63:0] io_a, // @[playground/src/noop/muldiv.scala 66:16]
  input  [63:0] io_b, // @[playground/src/noop/muldiv.scala 66:16]
  input         io_sign, // @[playground/src/noop/muldiv.scala 66:16]
  input         io_en, // @[playground/src/noop/muldiv.scala 66:16]
  output [63:0] io_qua, // @[playground/src/noop/muldiv.scala 66:16]
  output [63:0] io_rem, // @[playground/src/noop/muldiv.scala 66:16]
  output        io_valid // @[playground/src/noop/muldiv.scala 66:16]
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [127:0] _RAND_1;
  reg [127:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
`endif // RANDOMIZE_REG_INIT
  reg [63:0] quatient; // @[playground/src/noop/muldiv.scala 67:27]
  reg [127:0] val1; // @[playground/src/noop/muldiv.scala 68:26]
  reg [127:0] val2; // @[playground/src/noop/muldiv.scala 69:26]
  reg  qua_sign; // @[playground/src/noop/muldiv.scala 70:27]
  reg  rem_sign; // @[playground/src/noop/muldiv.scala 71:27]
  reg [6:0] iter; // @[playground/src/noop/muldiv.scala 72:26]
  reg  pre_alu64; // @[playground/src/noop/muldiv.scala 73:28]
  reg [1:0] state; // @[playground/src/noop/muldiv.scala 75:24]
  wire  _val1_T_3 = io_sign & io_a[63]; // @[playground/src/noop/muldiv.scala 84:61]
  wire [63:0] _val1_T_4 = ~io_a; // @[playground/src/noop/muldiv.scala 84:82]
  wire [63:0] _val1_T_6 = _val1_T_4 + 64'h1; // @[playground/src/noop/muldiv.scala 84:87]
  wire [63:0] _val1_T_7 = io_sign & io_a[63] ? _val1_T_6 : io_a; // @[playground/src/noop/muldiv.scala 84:52]
  wire [127:0] _val1_T_8 = {64'h0,_val1_T_7}; // @[playground/src/noop/muldiv.scala 84:28]
  wire [63:0] _val2_T_3 = ~io_b; // @[playground/src/noop/muldiv.scala 85:62]
  wire [63:0] _val2_T_5 = _val2_T_3 + 64'h1; // @[playground/src/noop/muldiv.scala 85:67]
  wire [63:0] _val2_T_6 = io_sign & io_b[63] ? _val2_T_5 : io_b; // @[playground/src/noop/muldiv.scala 85:32]
  wire [127:0] _val2_T_8 = {_val2_T_6,64'h0}; // @[playground/src/noop/muldiv.scala 85:28]
  wire [6:0] _iter_T_1 = iter + 7'h1; // @[playground/src/noop/muldiv.scala 95:30]
  wire [63:0] _quatient_T_1 = {quatient[62:0],1'h1}; // @[playground/src/noop/muldiv.scala 97:36]
  wire [127:0] _val1_T_10 = val1 - val2; // @[playground/src/noop/muldiv.scala 98:34]
  wire [127:0] _val2_T_9 = {{1'd0}, val2[127:1]}; // @[playground/src/noop/muldiv.scala 99:34]
  wire [63:0] _quatient_T_3 = {quatient[62:0],1'h0}; // @[playground/src/noop/muldiv.scala 101:36]
  wire [63:0] _GEN_8 = val1 >= val2 ? _quatient_T_1 : _quatient_T_3; // @[playground/src/noop/muldiv.scala 101:30 96:35 97:30]
  wire [127:0] _GEN_9 = val1 >= val2 ? _val1_T_10 : val1; // @[playground/src/noop/muldiv.scala 68:26 96:35 98:26]
  wire [127:0] _GEN_10 = val1 >= val2 ? _val2_T_9 : _val2_T_9; // @[playground/src/noop/muldiv.scala 102:26 96:35 99:26]
  wire [63:0] _sign_qua_T = ~quatient; // @[playground/src/noop/muldiv.scala 107:46]
  wire [63:0] _sign_qua_T_2 = _sign_qua_T + 64'h1; // @[playground/src/noop/muldiv.scala 107:56]
  wire [63:0] sign_qua = qua_sign ? _sign_qua_T_2 : quatient; // @[playground/src/noop/muldiv.scala 107:35]
  wire [63:0] _sign_rem_T_1 = ~val1[63:0]; // @[playground/src/noop/muldiv.scala 108:46]
  wire [63:0] _sign_rem_T_3 = _sign_rem_T_1 + 64'h1; // @[playground/src/noop/muldiv.scala 108:58]
  wire [63:0] sign_rem = rem_sign ? _sign_rem_T_3 : val1[63:0]; // @[playground/src/noop/muldiv.scala 108:35]
  wire [31:0] _io_qua_T_2 = sign_qua[31] ? 32'hffffffff : 32'h0; // @[playground/src/noop/muldiv.scala 109:62]
  wire [63:0] _io_qua_T_4 = {_io_qua_T_2,sign_qua[31:0]}; // @[playground/src/noop/muldiv.scala 109:57]
  wire [63:0] _io_qua_T_5 = pre_alu64 ? sign_qua : _io_qua_T_4; // @[playground/src/noop/muldiv.scala 109:32]
  wire [31:0] _io_rem_T_2 = sign_rem[31] ? 32'hffffffff : 32'h0; // @[playground/src/noop/muldiv.scala 110:62]
  wire [63:0] _io_rem_T_4 = {_io_rem_T_2,sign_rem[31:0]}; // @[playground/src/noop/muldiv.scala 110:57]
  wire [63:0] _io_rem_T_5 = pre_alu64 ? sign_rem : _io_rem_T_4; // @[playground/src/noop/muldiv.scala 110:32]
  wire  _GEN_16 = iter <= 7'h40 ? 1'h0 : 1'h1; // @[playground/src/noop/muldiv.scala 79:14 106:26 94:39]
  wire [63:0] _GEN_17 = iter <= 7'h40 ? 64'h0 : _io_qua_T_5; // @[playground/src/noop/muldiv.scala 77:12 109:26 94:39]
  wire [63:0] _GEN_18 = iter <= 7'h40 ? 64'h0 : _io_rem_T_5; // @[playground/src/noop/muldiv.scala 78:12 110:26 94:39]
  wire [63:0] _GEN_25 = 2'h1 == state ? _GEN_17 : 64'h0; // @[playground/src/noop/muldiv.scala 77:12 80:18]
  wire [63:0] _GEN_26 = 2'h1 == state ? _GEN_18 : 64'h0; // @[playground/src/noop/muldiv.scala 78:12 80:18]
  assign io_qua = 2'h0 == state ? 64'h0 : _GEN_25; // @[playground/src/noop/muldiv.scala 77:12 80:18]
  assign io_rem = 2'h0 == state ? 64'h0 : _GEN_26; // @[playground/src/noop/muldiv.scala 78:12 80:18]
  assign io_valid = 2'h0 == state ? 1'h0 : 2'h1 == state & _GEN_16; // @[playground/src/noop/muldiv.scala 79:14 80:18]
  always @(posedge clock) begin
    if (reset) begin // @[playground/src/noop/muldiv.scala 67:27]
      quatient <= 64'h0; // @[playground/src/noop/muldiv.scala 67:27]
    end else if (2'h0 == state) begin // @[playground/src/noop/muldiv.scala 80:18]
      if (io_en) begin // @[playground/src/noop/muldiv.scala 82:24]
        quatient <= 64'h0; // @[playground/src/noop/muldiv.scala 89:26]
      end
    end else if (2'h1 == state) begin // @[playground/src/noop/muldiv.scala 80:18]
      if (iter <= 7'h40) begin // @[playground/src/noop/muldiv.scala 94:39]
        quatient <= _GEN_8;
      end
    end
    if (reset) begin // @[playground/src/noop/muldiv.scala 68:26]
      val1 <= 128'h0; // @[playground/src/noop/muldiv.scala 68:26]
    end else if (2'h0 == state) begin // @[playground/src/noop/muldiv.scala 80:18]
      if (io_en) begin // @[playground/src/noop/muldiv.scala 82:24]
        val1 <= _val1_T_8; // @[playground/src/noop/muldiv.scala 84:22]
      end
    end else if (2'h1 == state) begin // @[playground/src/noop/muldiv.scala 80:18]
      if (iter <= 7'h40) begin // @[playground/src/noop/muldiv.scala 94:39]
        val1 <= _GEN_9;
      end
    end
    if (reset) begin // @[playground/src/noop/muldiv.scala 69:26]
      val2 <= 128'h0; // @[playground/src/noop/muldiv.scala 69:26]
    end else if (2'h0 == state) begin // @[playground/src/noop/muldiv.scala 80:18]
      if (io_en) begin // @[playground/src/noop/muldiv.scala 82:24]
        val2 <= _val2_T_8; // @[playground/src/noop/muldiv.scala 85:22]
      end
    end else if (2'h1 == state) begin // @[playground/src/noop/muldiv.scala 80:18]
      if (iter <= 7'h40) begin // @[playground/src/noop/muldiv.scala 94:39]
        val2 <= _GEN_10;
      end
    end
    if (reset) begin // @[playground/src/noop/muldiv.scala 70:27]
      qua_sign <= 1'h0; // @[playground/src/noop/muldiv.scala 70:27]
    end else if (2'h0 == state) begin // @[playground/src/noop/muldiv.scala 80:18]
      if (io_en) begin // @[playground/src/noop/muldiv.scala 82:24]
        qua_sign <= io_sign & (io_a[63] != io_b[63] & io_b != 64'h0); // @[playground/src/noop/muldiv.scala 86:26]
      end
    end
    if (reset) begin // @[playground/src/noop/muldiv.scala 71:27]
      rem_sign <= 1'h0; // @[playground/src/noop/muldiv.scala 71:27]
    end else if (2'h0 == state) begin // @[playground/src/noop/muldiv.scala 80:18]
      if (io_en) begin // @[playground/src/noop/muldiv.scala 82:24]
        rem_sign <= _val1_T_3; // @[playground/src/noop/muldiv.scala 87:26]
      end
    end
    if (reset) begin // @[playground/src/noop/muldiv.scala 72:26]
      iter <= 7'h0; // @[playground/src/noop/muldiv.scala 72:26]
    end else if (2'h0 == state) begin // @[playground/src/noop/muldiv.scala 80:18]
      if (io_en) begin // @[playground/src/noop/muldiv.scala 82:24]
        iter <= 7'h0; // @[playground/src/noop/muldiv.scala 90:22]
      end
    end else if (2'h1 == state) begin // @[playground/src/noop/muldiv.scala 80:18]
      if (iter <= 7'h40) begin // @[playground/src/noop/muldiv.scala 94:39]
        iter <= _iter_T_1; // @[playground/src/noop/muldiv.scala 95:22]
      end
    end
    if (reset) begin // @[playground/src/noop/muldiv.scala 73:28]
      pre_alu64 <= 1'h0; // @[playground/src/noop/muldiv.scala 73:28]
    end else if (2'h0 == state) begin // @[playground/src/noop/muldiv.scala 80:18]
      if (io_en) begin // @[playground/src/noop/muldiv.scala 82:24]
        pre_alu64 <= io_alu64; // @[playground/src/noop/muldiv.scala 88:27]
      end
    end
    if (reset) begin // @[playground/src/noop/muldiv.scala 75:24]
      state <= 2'h0; // @[playground/src/noop/muldiv.scala 75:24]
    end else if (2'h0 == state) begin // @[playground/src/noop/muldiv.scala 80:18]
      if (io_en) begin // @[playground/src/noop/muldiv.scala 82:24]
        state <= 2'h1; // @[playground/src/noop/muldiv.scala 83:23]
      end
    end else if (2'h1 == state) begin // @[playground/src/noop/muldiv.scala 80:18]
      if (!(iter <= 7'h40)) begin // @[playground/src/noop/muldiv.scala 94:39]
        state <= 2'h0; // @[playground/src/noop/muldiv.scala 105:23]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  quatient = _RAND_0[63:0];
  _RAND_1 = {4{`RANDOM}};
  val1 = _RAND_1[127:0];
  _RAND_2 = {4{`RANDOM}};
  val2 = _RAND_2[127:0];
  _RAND_3 = {1{`RANDOM}};
  qua_sign = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  rem_sign = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  iter = _RAND_5[6:0];
  _RAND_6 = {1{`RANDOM}};
  pre_alu64 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  state = _RAND_7[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ALU(
  input         clock,
  input         reset,
  input  [4:0]  io_alu_op, // @[playground/src/noop/alu.scala 39:16]
  input  [63:0] io_val1, // @[playground/src/noop/alu.scala 39:16]
  input  [63:0] io_val2, // @[playground/src/noop/alu.scala 39:16]
  input         io_alu64, // @[playground/src/noop/alu.scala 39:16]
  input         io_en, // @[playground/src/noop/alu.scala 39:16]
  output [63:0] io_out, // @[playground/src/noop/alu.scala 39:16]
  output        io_valid // @[playground/src/noop/alu.scala 39:16]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  wire  multiplier_clock; // @[playground/src/noop/alu.scala 40:28]
  wire  multiplier_reset; // @[playground/src/noop/alu.scala 40:28]
  wire [63:0] multiplier_io_a; // @[playground/src/noop/alu.scala 40:28]
  wire [63:0] multiplier_io_b; // @[playground/src/noop/alu.scala 40:28]
  wire [4:0] multiplier_io_aluop; // @[playground/src/noop/alu.scala 40:28]
  wire  multiplier_io_en; // @[playground/src/noop/alu.scala 40:28]
  wire [63:0] multiplier_io_out; // @[playground/src/noop/alu.scala 40:28]
  wire  multiplier_io_valid; // @[playground/src/noop/alu.scala 40:28]
  wire  divider_clock; // @[playground/src/noop/alu.scala 41:28]
  wire  divider_reset; // @[playground/src/noop/alu.scala 41:28]
  wire  divider_io_alu64; // @[playground/src/noop/alu.scala 41:28]
  wire [63:0] divider_io_a; // @[playground/src/noop/alu.scala 41:28]
  wire [63:0] divider_io_b; // @[playground/src/noop/alu.scala 41:28]
  wire  divider_io_sign; // @[playground/src/noop/alu.scala 41:28]
  wire  divider_io_en; // @[playground/src/noop/alu.scala 41:28]
  wire [63:0] divider_io_qua; // @[playground/src/noop/alu.scala 41:28]
  wire [63:0] divider_io_rem; // @[playground/src/noop/alu.scala 41:28]
  wire  divider_io_valid; // @[playground/src/noop/alu.scala 41:28]
  reg [4:0] pre_aluop; // @[playground/src/noop/alu.scala 43:28]
  reg [1:0] state; // @[playground/src/noop/alu.scala 44:24]
  wire  _div_type_T_1 = 5'h11 == io_alu_op; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _div_type_T_3 = 5'h12 == io_alu_op; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _div_type_T_5 = 5'h13 == io_alu_op; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _div_type_T_13 = _div_type_T_3 ? 1'h0 : _div_type_T_5; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  _T_7 = io_alu_op == 5'hd | io_alu_op == 5'he | io_alu_op == 5'hf | io_alu_op == 5'h10; // @[playground/src/noop/alu.scala 63:97]
  wire  _T_14 = io_alu_op == 5'h11 | io_alu_op == 5'h12 | io_alu_op == 5'h13 | io_alu_op == 5'h14; // @[playground/src/noop/alu.scala 66:102]
  wire [63:0] _alu_val_T_1 = io_val1 + io_val2; // @[playground/src/noop/alu.scala 75:49]
  wire [63:0] _alu_val_T_2 = io_val1 ^ io_val2; // @[playground/src/noop/alu.scala 76:49]
  wire [63:0] _alu_val_T_3 = io_val1 | io_val2; // @[playground/src/noop/alu.scala 77:49]
  wire [63:0] _alu_val_T_4 = io_val1 & io_val2; // @[playground/src/noop/alu.scala 78:49]
  wire [126:0] _GEN_33 = {{63'd0}, io_val1}; // @[playground/src/noop/alu.scala 79:49]
  wire [126:0] _alu_val_T_6 = _GEN_33 << io_val2[5:0]; // @[playground/src/noop/alu.scala 79:49]
  wire [63:0] _alu_val_T_8 = io_val1 >> io_val2[5:0]; // @[playground/src/noop/alu.scala 80:63]
  wire [31:0] _alu_val_T_11 = io_val1[31:0] >> io_val2[5:0]; // @[playground/src/noop/alu.scala 80:104]
  wire [63:0] _alu_val_T_12 = io_alu64 ? _alu_val_T_8 : {{32'd0}, _alu_val_T_11}; // @[playground/src/noop/alu.scala 80:43]
  wire [63:0] _alu_val_T_16 = $signed(io_val1) >>> io_val2[5:0]; // @[playground/src/noop/alu.scala 81:87]
  wire [31:0] _alu_val_T_18 = io_val1[31:0]; // @[playground/src/noop/alu.scala 81:112]
  wire [31:0] _alu_val_T_21 = $signed(_alu_val_T_18) >>> io_val2[5:0]; // @[playground/src/noop/alu.scala 81:136]
  wire [63:0] _alu_val_T_22 = io_alu64 ? _alu_val_T_16 : {{32'd0}, _alu_val_T_21}; // @[playground/src/noop/alu.scala 81:43]
  wire [63:0] _alu_val_T_24 = io_val1 - io_val2; // @[playground/src/noop/alu.scala 82:49]
  wire  _alu_val_T_27 = $signed(io_val1) < $signed(io_val2); // @[playground/src/noop/alu.scala 83:59]
  wire  _alu_val_T_29 = io_val1 < io_val2; // @[playground/src/noop/alu.scala 84:52]
  wire [63:0] _alu_val_T_31 = ~io_val1; // @[playground/src/noop/alu.scala 85:42]
  wire [63:0] _alu_val_T_32 = _alu_val_T_31 & io_val2; // @[playground/src/noop/alu.scala 85:52]
  wire [63:0] _alu_val_T_36 = 5'h1 == io_alu_op ? io_val1 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 81:58]
  wire [63:0] _alu_val_T_38 = 5'h2 == io_alu_op ? io_val2 : _alu_val_T_36; // @[src/main/scala/chisel3/util/Mux.scala 81:58]
  wire [63:0] _alu_val_T_40 = 5'h3 == io_alu_op ? _alu_val_T_1 : _alu_val_T_38; // @[src/main/scala/chisel3/util/Mux.scala 81:58]
  wire [63:0] _alu_val_T_42 = 5'h4 == io_alu_op ? _alu_val_T_2 : _alu_val_T_40; // @[src/main/scala/chisel3/util/Mux.scala 81:58]
  wire [63:0] _alu_val_T_44 = 5'h5 == io_alu_op ? _alu_val_T_3 : _alu_val_T_42; // @[src/main/scala/chisel3/util/Mux.scala 81:58]
  wire [63:0] _alu_val_T_46 = 5'h6 == io_alu_op ? _alu_val_T_4 : _alu_val_T_44; // @[src/main/scala/chisel3/util/Mux.scala 81:58]
  wire [126:0] _alu_val_T_48 = 5'h7 == io_alu_op ? _alu_val_T_6 : {{63'd0}, _alu_val_T_46}; // @[src/main/scala/chisel3/util/Mux.scala 81:58]
  wire [126:0] _alu_val_T_50 = 5'h8 == io_alu_op ? {{63'd0}, _alu_val_T_12} : _alu_val_T_48; // @[src/main/scala/chisel3/util/Mux.scala 81:58]
  wire [126:0] _alu_val_T_52 = 5'h9 == io_alu_op ? {{63'd0}, _alu_val_T_22} : _alu_val_T_50; // @[src/main/scala/chisel3/util/Mux.scala 81:58]
  wire [126:0] _alu_val_T_54 = 5'ha == io_alu_op ? {{63'd0}, _alu_val_T_24} : _alu_val_T_52; // @[src/main/scala/chisel3/util/Mux.scala 81:58]
  wire [126:0] _alu_val_T_56 = 5'hb == io_alu_op ? {{126'd0}, _alu_val_T_27} : _alu_val_T_54; // @[src/main/scala/chisel3/util/Mux.scala 81:58]
  wire [126:0] _alu_val_T_58 = 5'hc == io_alu_op ? {{126'd0}, _alu_val_T_29} : _alu_val_T_56; // @[src/main/scala/chisel3/util/Mux.scala 81:58]
  wire [126:0] alu_val = 5'h15 == io_alu_op ? {{63'd0}, _alu_val_T_32} : _alu_val_T_58; // @[src/main/scala/chisel3/util/Mux.scala 81:58]
  wire [1:0] _GEN_1 = io_alu_op == 5'h11 | io_alu_op == 5'h12 | io_alu_op == 5'h13 | io_alu_op == 5'h14 ? 2'h2 : state; // @[playground/src/noop/alu.scala 66:129 44:24 68:27]
  wire [126:0] _GEN_2 = io_alu_op == 5'h11 | io_alu_op == 5'h12 | io_alu_op == 5'h13 | io_alu_op == 5'h14 ? 127'h0 :
    alu_val; // @[playground/src/noop/alu.scala 66:129 57:14 87:28]
  wire  _GEN_3 = io_alu_op == 5'h11 | io_alu_op == 5'h12 | io_alu_op == 5'h13 | io_alu_op == 5'h14 ? 1'h0 : 1'h1; // @[playground/src/noop/alu.scala 66:129 56:14 88:30]
  wire  _GEN_6 = io_alu_op == 5'hd | io_alu_op == 5'he | io_alu_op == 5'hf | io_alu_op == 5'h10 ? 1'h0 : _T_14; // @[playground/src/noop/alu.scala 63:125 55:25]
  wire [126:0] _GEN_7 = io_alu_op == 5'hd | io_alu_op == 5'he | io_alu_op == 5'hf | io_alu_op == 5'h10 ? 127'h0 : _GEN_2
    ; // @[playground/src/noop/alu.scala 63:125 57:14]
  wire  _GEN_8 = io_alu_op == 5'hd | io_alu_op == 5'he | io_alu_op == 5'hf | io_alu_op == 5'h10 ? 1'h0 : _GEN_3; // @[playground/src/noop/alu.scala 63:125 56:14]
  wire  _GEN_10 = io_en & _T_7; // @[playground/src/noop/alu.scala 61:24 48:25]
  wire  _GEN_12 = io_en & _GEN_6; // @[playground/src/noop/alu.scala 61:24 55:25]
  wire [126:0] _GEN_13 = io_en ? _GEN_7 : 127'h0; // @[playground/src/noop/alu.scala 57:14 61:24]
  wire  _GEN_14 = io_en & _GEN_8; // @[playground/src/noop/alu.scala 56:14 61:24]
  wire [63:0] _GEN_15 = multiplier_io_valid ? multiplier_io_out : 64'h0; // @[playground/src/noop/alu.scala 57:14 93:38 94:24]
  wire  _GEN_16 = multiplier_io_valid; // @[playground/src/noop/alu.scala 56:14 93:38 95:26]
  wire [63:0] _io_out_T_3 = pre_aluop == 5'h11 | pre_aluop == 5'h12 ? divider_io_qua : divider_io_rem; // @[playground/src/noop/alu.scala 101:30]
  wire [63:0] _GEN_18 = divider_io_valid ? _io_out_T_3 : 64'h0; // @[playground/src/noop/alu.scala 100:35 101:24 57:14]
  wire  _GEN_19 = divider_io_valid; // @[playground/src/noop/alu.scala 100:35 102:26 56:14]
  wire [1:0] _GEN_20 = divider_io_valid ? 2'h0 : state; // @[playground/src/noop/alu.scala 100:35 103:23 44:24]
  wire [63:0] _GEN_21 = 2'h2 == state ? _GEN_18 : 64'h0; // @[playground/src/noop/alu.scala 57:14 59:18]
  wire  _GEN_22 = 2'h2 == state & _GEN_19; // @[playground/src/noop/alu.scala 56:14 59:18]
  wire [63:0] _GEN_24 = 2'h1 == state ? _GEN_15 : _GEN_21; // @[playground/src/noop/alu.scala 59:18]
  wire  _GEN_25 = 2'h1 == state ? _GEN_16 : _GEN_22; // @[playground/src/noop/alu.scala 59:18]
  wire [126:0] _GEN_31 = 2'h0 == state ? _GEN_13 : {{63'd0}, _GEN_24}; // @[playground/src/noop/alu.scala 59:18]
  MUL multiplier ( // @[playground/src/noop/alu.scala 40:28]
    .clock(multiplier_clock),
    .reset(multiplier_reset),
    .io_a(multiplier_io_a),
    .io_b(multiplier_io_b),
    .io_aluop(multiplier_io_aluop),
    .io_en(multiplier_io_en),
    .io_out(multiplier_io_out),
    .io_valid(multiplier_io_valid)
  );
  DIV divider ( // @[playground/src/noop/alu.scala 41:28]
    .clock(divider_clock),
    .reset(divider_reset),
    .io_alu64(divider_io_alu64),
    .io_a(divider_io_a),
    .io_b(divider_io_b),
    .io_sign(divider_io_sign),
    .io_en(divider_io_en),
    .io_qua(divider_io_qua),
    .io_rem(divider_io_rem),
    .io_valid(divider_io_valid)
  );
  assign io_out = _GEN_31[63:0];
  assign io_valid = 2'h0 == state ? _GEN_14 : _GEN_25; // @[playground/src/noop/alu.scala 59:18]
  assign multiplier_clock = clock;
  assign multiplier_reset = reset;
  assign multiplier_io_a = io_val1; // @[playground/src/noop/alu.scala 46:25]
  assign multiplier_io_b = io_val2; // @[playground/src/noop/alu.scala 47:25]
  assign multiplier_io_aluop = io_alu_op; // @[playground/src/noop/alu.scala 49:26]
  assign multiplier_io_en = 2'h0 == state & _GEN_10; // @[playground/src/noop/alu.scala 59:18 48:25]
  assign divider_clock = clock;
  assign divider_reset = reset;
  assign divider_io_alu64 = io_alu64; // @[playground/src/noop/alu.scala 51:25]
  assign divider_io_a = io_val1; // @[playground/src/noop/alu.scala 52:25]
  assign divider_io_b = io_val2; // @[playground/src/noop/alu.scala 53:25]
  assign divider_io_sign = _div_type_T_1 | _div_type_T_13; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  assign divider_io_en = 2'h0 == state & _GEN_12; // @[playground/src/noop/alu.scala 59:18 55:25]
  always @(posedge clock) begin
    if (reset) begin // @[playground/src/noop/alu.scala 43:28]
      pre_aluop <= 5'h0; // @[playground/src/noop/alu.scala 43:28]
    end else if (2'h0 == state) begin // @[playground/src/noop/alu.scala 59:18]
      if (io_en) begin // @[playground/src/noop/alu.scala 61:24]
        pre_aluop <= io_alu_op; // @[playground/src/noop/alu.scala 62:27]
      end
    end
    if (reset) begin // @[playground/src/noop/alu.scala 44:24]
      state <= 2'h0; // @[playground/src/noop/alu.scala 44:24]
    end else if (2'h0 == state) begin // @[playground/src/noop/alu.scala 59:18]
      if (io_en) begin // @[playground/src/noop/alu.scala 61:24]
        if (io_alu_op == 5'hd | io_alu_op == 5'he | io_alu_op == 5'hf | io_alu_op == 5'h10) begin // @[playground/src/noop/alu.scala 63:125]
          state <= 2'h1; // @[playground/src/noop/alu.scala 65:27]
        end else begin
          state <= _GEN_1;
        end
      end
    end else if (2'h1 == state) begin // @[playground/src/noop/alu.scala 59:18]
      if (multiplier_io_valid) begin // @[playground/src/noop/alu.scala 93:38]
        state <= 2'h0; // @[playground/src/noop/alu.scala 96:23]
      end
    end else if (2'h2 == state) begin // @[playground/src/noop/alu.scala 59:18]
      state <= _GEN_20;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  pre_aluop = _RAND_0[4:0];
  _RAND_1 = {1{`RANDOM}};
  state = _RAND_1[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module BranchALU(
  input  [63:0] io_val1, // @[playground/src/noop/alu.scala 117:16]
  input  [63:0] io_val2, // @[playground/src/noop/alu.scala 117:16]
  input  [2:0]  io_brType, // @[playground/src/noop/alu.scala 117:16]
  output        io_is_jmp // @[playground/src/noop/alu.scala 117:16]
);
  wire  _io_is_jmp_T = io_val1 == io_val2; // @[playground/src/noop/alu.scala 119:29]
  wire  _io_is_jmp_T_1 = io_val1 != io_val2; // @[playground/src/noop/alu.scala 120:29]
  wire  _io_is_jmp_T_4 = $signed(io_val1) < $signed(io_val2); // @[playground/src/noop/alu.scala 121:36]
  wire  _io_is_jmp_T_7 = $signed(io_val1) >= $signed(io_val2); // @[playground/src/noop/alu.scala 122:36]
  wire  _io_is_jmp_T_8 = io_val1 < io_val2; // @[playground/src/noop/alu.scala 123:29]
  wire  _io_is_jmp_T_9 = io_val1 >= io_val2; // @[playground/src/noop/alu.scala 124:29]
  wire  _io_is_jmp_T_13 = 3'h1 == io_brType ? _io_is_jmp_T_1 : 3'h0 == io_brType & _io_is_jmp_T; // @[src/main/scala/chisel3/util/Mux.scala 81:58]
  wire  _io_is_jmp_T_15 = 3'h4 == io_brType ? _io_is_jmp_T_4 : _io_is_jmp_T_13; // @[src/main/scala/chisel3/util/Mux.scala 81:58]
  wire  _io_is_jmp_T_17 = 3'h5 == io_brType ? _io_is_jmp_T_7 : _io_is_jmp_T_15; // @[src/main/scala/chisel3/util/Mux.scala 81:58]
  wire  _io_is_jmp_T_19 = 3'h6 == io_brType ? _io_is_jmp_T_8 : _io_is_jmp_T_17; // @[src/main/scala/chisel3/util/Mux.scala 81:58]
  assign io_is_jmp = 3'h7 == io_brType ? _io_is_jmp_T_9 : _io_is_jmp_T_19; // @[src/main/scala/chisel3/util/Mux.scala 81:58]
endmodule
module Execute(
  input         clock,
  input         reset,
  input  [31:0] io_rr2ex_inst, // @[playground/src/noop/execute.scala 14:16]
  input  [63:0] io_rr2ex_pc, // @[playground/src/noop/execute.scala 14:16]
  input  [63:0] io_rr2ex_excep_cause, // @[playground/src/noop/execute.scala 14:16]
  input  [63:0] io_rr2ex_excep_tval, // @[playground/src/noop/execute.scala 14:16]
  input         io_rr2ex_excep_en, // @[playground/src/noop/execute.scala 14:16]
  input  [63:0] io_rr2ex_excep_pc, // @[playground/src/noop/execute.scala 14:16]
  input  [1:0]  io_rr2ex_excep_etype, // @[playground/src/noop/execute.scala 14:16]
  input  [4:0]  io_rr2ex_ctrl_aluOp, // @[playground/src/noop/execute.scala 14:16]
  input         io_rr2ex_ctrl_aluWidth, // @[playground/src/noop/execute.scala 14:16]
  input  [4:0]  io_rr2ex_ctrl_dcMode, // @[playground/src/noop/execute.scala 14:16]
  input         io_rr2ex_ctrl_writeRegEn, // @[playground/src/noop/execute.scala 14:16]
  input         io_rr2ex_ctrl_writeCSREn, // @[playground/src/noop/execute.scala 14:16]
  input  [2:0]  io_rr2ex_ctrl_brType, // @[playground/src/noop/execute.scala 14:16]
  input  [63:0] io_rr2ex_rs1_d, // @[playground/src/noop/execute.scala 14:16]
  input  [11:0] io_rr2ex_rs2, // @[playground/src/noop/execute.scala 14:16]
  input  [63:0] io_rr2ex_rs2_d, // @[playground/src/noop/execute.scala 14:16]
  input  [4:0]  io_rr2ex_dst, // @[playground/src/noop/execute.scala 14:16]
  input  [63:0] io_rr2ex_dst_d, // @[playground/src/noop/execute.scala 14:16]
  input  [11:0] io_rr2ex_rcsr_id, // @[playground/src/noop/execute.scala 14:16]
  input  [1:0]  io_rr2ex_jmp_type, // @[playground/src/noop/execute.scala 14:16]
  input  [1:0]  io_rr2ex_special, // @[playground/src/noop/execute.scala 14:16]
  input  [1:0]  io_rr2ex_indi, // @[playground/src/noop/execute.scala 14:16]
  output        io_rr2ex_drop, // @[playground/src/noop/execute.scala 14:16]
  output        io_rr2ex_stall, // @[playground/src/noop/execute.scala 14:16]
  input         io_rr2ex_recov, // @[playground/src/noop/execute.scala 14:16]
  input         io_rr2ex_valid, // @[playground/src/noop/execute.scala 14:16]
  output        io_rr2ex_ready, // @[playground/src/noop/execute.scala 14:16]
  output [31:0] io_ex2mem_inst, // @[playground/src/noop/execute.scala 14:16]
  output [63:0] io_ex2mem_pc, // @[playground/src/noop/execute.scala 14:16]
  output [63:0] io_ex2mem_excep_cause, // @[playground/src/noop/execute.scala 14:16]
  output [63:0] io_ex2mem_excep_tval, // @[playground/src/noop/execute.scala 14:16]
  output        io_ex2mem_excep_en, // @[playground/src/noop/execute.scala 14:16]
  output [63:0] io_ex2mem_excep_pc, // @[playground/src/noop/execute.scala 14:16]
  output [1:0]  io_ex2mem_excep_etype, // @[playground/src/noop/execute.scala 14:16]
  output [4:0]  io_ex2mem_ctrl_dcMode, // @[playground/src/noop/execute.scala 14:16]
  output        io_ex2mem_ctrl_writeRegEn, // @[playground/src/noop/execute.scala 14:16]
  output        io_ex2mem_ctrl_writeCSREn, // @[playground/src/noop/execute.scala 14:16]
  output [63:0] io_ex2mem_mem_addr, // @[playground/src/noop/execute.scala 14:16]
  output [63:0] io_ex2mem_mem_data, // @[playground/src/noop/execute.scala 14:16]
  output [11:0] io_ex2mem_csr_id, // @[playground/src/noop/execute.scala 14:16]
  output [63:0] io_ex2mem_csr_d, // @[playground/src/noop/execute.scala 14:16]
  output [4:0]  io_ex2mem_dst, // @[playground/src/noop/execute.scala 14:16]
  output [63:0] io_ex2mem_dst_d, // @[playground/src/noop/execute.scala 14:16]
  output [11:0] io_ex2mem_rcsr_id, // @[playground/src/noop/execute.scala 14:16]
  output [1:0]  io_ex2mem_special, // @[playground/src/noop/execute.scala 14:16]
  output [1:0]  io_ex2mem_indi, // @[playground/src/noop/execute.scala 14:16]
  input         io_ex2mem_drop, // @[playground/src/noop/execute.scala 14:16]
  input         io_ex2mem_stall, // @[playground/src/noop/execute.scala 14:16]
  output        io_ex2mem_recov, // @[playground/src/noop/execute.scala 14:16]
  output        io_ex2mem_valid, // @[playground/src/noop/execute.scala 14:16]
  input         io_ex2mem_ready, // @[playground/src/noop/execute.scala 14:16]
  output [4:0]  io_d_ex_id, // @[playground/src/noop/execute.scala 14:16]
  output [63:0] io_d_ex_data, // @[playground/src/noop/execute.scala 14:16]
  output [1:0]  io_d_ex_state, // @[playground/src/noop/execute.scala 14:16]
  output [63:0] io_ex2if_seq_pc, // @[playground/src/noop/execute.scala 14:16]
  output        io_ex2if_valid, // @[playground/src/noop/execute.scala 14:16]
  input  [63:0] io_updateNextPc_seq_pc, // @[playground/src/noop/execute.scala 14:16]
  input         io_updateNextPc_valid // @[playground/src/noop/execute.scala 14:16]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [63:0] _RAND_12;
  reg [63:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [63:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [63:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [63:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [63:0] _RAND_27;
  reg [31:0] _RAND_28;
`endif // RANDOMIZE_REG_INIT
  wire  alu_clock; // @[playground/src/noop/execute.scala 27:25]
  wire  alu_reset; // @[playground/src/noop/execute.scala 27:25]
  wire [4:0] alu_io_alu_op; // @[playground/src/noop/execute.scala 27:25]
  wire [63:0] alu_io_val1; // @[playground/src/noop/execute.scala 27:25]
  wire [63:0] alu_io_val2; // @[playground/src/noop/execute.scala 27:25]
  wire  alu_io_alu64; // @[playground/src/noop/execute.scala 27:25]
  wire  alu_io_en; // @[playground/src/noop/execute.scala 27:25]
  wire [63:0] alu_io_out; // @[playground/src/noop/execute.scala 27:25]
  wire  alu_io_valid; // @[playground/src/noop/execute.scala 27:25]
  wire [63:0] branchAlu_io_val1; // @[playground/src/noop/execute.scala 153:27]
  wire [63:0] branchAlu_io_val2; // @[playground/src/noop/execute.scala 153:27]
  wire [2:0] branchAlu_io_brType; // @[playground/src/noop/execute.scala 153:27]
  wire  branchAlu_io_is_jmp; // @[playground/src/noop/execute.scala 153:27]
  reg  drop_r; // @[playground/src/noop/execute.scala 21:25]
  reg  stall_r; // @[playground/src/noop/execute.scala 22:26]
  wire  drop_in = drop_r | io_ex2mem_drop; // @[playground/src/noop/execute.scala 24:26]
  wire  _io_rr2ex_stall_T = ~io_ex2mem_drop; // @[playground/src/noop/execute.scala 26:55]
  reg [31:0] inst_r; // @[playground/src/noop/execute.scala 28:30]
  reg [63:0] pc_r; // @[playground/src/noop/execute.scala 29:30]
  reg [63:0] excep_r_cause; // @[playground/src/noop/execute.scala 30:30]
  reg [63:0] excep_r_tval; // @[playground/src/noop/execute.scala 30:30]
  reg  excep_r_en; // @[playground/src/noop/execute.scala 30:30]
  reg [63:0] excep_r_pc; // @[playground/src/noop/execute.scala 30:30]
  reg [1:0] excep_r_etype; // @[playground/src/noop/execute.scala 30:30]
  reg [4:0] ctrl_r_dcMode; // @[playground/src/noop/execute.scala 31:30]
  reg  ctrl_r_writeRegEn; // @[playground/src/noop/execute.scala 31:30]
  reg  ctrl_r_writeCSREn; // @[playground/src/noop/execute.scala 31:30]
  reg [63:0] mem_addr_r; // @[playground/src/noop/execute.scala 32:30]
  reg [63:0] mem_data_r; // @[playground/src/noop/execute.scala 33:30]
  reg [11:0] csr_id_r; // @[playground/src/noop/execute.scala 34:30]
  reg [63:0] csr_d_r; // @[playground/src/noop/execute.scala 35:30]
  reg [4:0] dst_r; // @[playground/src/noop/execute.scala 36:30]
  reg [63:0] dst_d_r; // @[playground/src/noop/execute.scala 37:30]
  reg [11:0] rcsr_id_r; // @[playground/src/noop/execute.scala 38:30]
  reg [1:0] special_r; // @[playground/src/noop/execute.scala 39:30]
  reg  alu64_r; // @[playground/src/noop/execute.scala 40:30]
  reg [1:0] indi_r; // @[playground/src/noop/execute.scala 41:30]
  reg [63:0] next_pc_r; // @[playground/src/noop/execute.scala 42:30]
  reg  recov_r; // @[playground/src/noop/execute.scala 43:30]
  reg  valid_r; // @[playground/src/noop/execute.scala 44:30]
  wire  hs_in = io_rr2ex_ready & io_rr2ex_valid; // @[playground/src/noop/execute.scala 46:34]
  wire  hs_out = io_ex2mem_ready & io_ex2mem_valid; // @[playground/src/noop/execute.scala 47:35]
  wire  alu64 = ~io_rr2ex_ctrl_aluWidth; // @[playground/src/noop/execute.scala 48:40]
  wire  _signed_dr_T = ~alu64; // @[playground/src/noop/execute.scala 51:23]
  wire  signed_dr = ~alu64 & (io_rr2ex_ctrl_aluOp == 5'h11 | io_rr2ex_ctrl_aluOp == 5'h13); // @[playground/src/noop/execute.scala 51:30]
  wire  unsigned_dr = _signed_dr_T & (io_rr2ex_ctrl_aluOp == 5'h12 | io_rr2ex_ctrl_aluOp == 5'h14); // @[playground/src/noop/execute.scala 52:30]
  wire [63:0] _val1_T_1 = {32'h0,io_rr2ex_rs1_d[31:0]}; // @[playground/src/noop/common.scala 712:12]
  wire [31:0] _val1_T_4 = io_rr2ex_rs1_d[31] ? 32'hffffffff : 32'h0; // @[playground/src/noop/common.scala 709:18]
  wire [63:0] _val1_T_6 = {_val1_T_4,io_rr2ex_rs1_d[31:0]}; // @[playground/src/noop/common.scala 709:13]
  wire [63:0] _val1_T_7 = signed_dr ? _val1_T_6 : io_rr2ex_rs1_d; // @[src/main/scala/chisel3/util/Mux.scala 47:70]
  wire  is_shift = io_rr2ex_ctrl_aluOp == 5'h7 | io_rr2ex_ctrl_aluOp == 5'h8 | io_rr2ex_ctrl_aluOp == 5'h9; // @[playground/src/noop/execute.scala 58:59]
  wire [63:0] _val2_T_1 = {32'h0,io_rr2ex_rs2_d[31:0]}; // @[playground/src/noop/common.scala 712:12]
  wire [31:0] _val2_T_4 = io_rr2ex_rs2_d[31] ? 32'hffffffff : 32'h0; // @[playground/src/noop/common.scala 709:18]
  wire [63:0] _val2_T_6 = {_val2_T_4,io_rr2ex_rs2_d[31:0]}; // @[playground/src/noop/common.scala 709:13]
  wire [5:0] _val2_T_9 = {1'h0,io_rr2ex_rs2_d[4:0]}; // @[playground/src/noop/execute.scala 62:60]
  wire [5:0] _val2_T_10 = alu64 ? io_rr2ex_rs2_d[5:0] : _val2_T_9; // @[playground/src/noop/execute.scala 62:28]
  wire [63:0] _val2_T_11 = is_shift ? {{58'd0}, _val2_T_10} : io_rr2ex_rs2_d; // @[src/main/scala/chisel3/util/Mux.scala 47:70]
  wire [63:0] _val2_T_12 = signed_dr ? _val2_T_6 : _val2_T_11; // @[src/main/scala/chisel3/util/Mux.scala 47:70]
  wire  cur_alu64 = hs_in ? alu64 : alu64_r; // @[playground/src/noop/execute.scala 70:26]
  wire [63:0] _alu_out_T = alu_io_out; // @[playground/src/noop/execute.scala 71:44]
  wire [31:0] _alu_out_T_3 = alu_io_out[31] ? 32'hffffffff : 32'h0; // @[playground/src/noop/common.scala 709:18]
  wire [63:0] _alu_out_T_5 = {_alu_out_T_3,alu_io_out[31:0]}; // @[playground/src/noop/common.scala 709:13]
  wire [63:0] alu_out = cur_alu64 ? _alu_out_T : _alu_out_T_5; // @[playground/src/noop/execute.scala 71:22]
  wire [63:0] _wdata_T_1 = io_rr2ex_ctrl_writeCSREn ? io_rr2ex_rs2_d : alu_out; // @[src/main/scala/chisel3/util/Mux.scala 47:70]
  wire [63:0] wdata = io_rr2ex_ctrl_dcMode[3] ? io_rr2ex_dst_d : _wdata_T_1; // @[src/main/scala/chisel3/util/Mux.scala 47:70]
  wire [63:0] _memAlign_ans_T = alu_out & 64'h1; // @[playground/src/noop/common.scala 329:27]
  wire  _memAlign_ans_T_1 = _memAlign_ans_T == 64'h0; // @[playground/src/noop/common.scala 329:36]
  wire [63:0] _memAlign_ans_T_2 = alu_out & 64'h3; // @[playground/src/noop/common.scala 330:27]
  wire  _memAlign_ans_T_3 = _memAlign_ans_T_2 == 64'h0; // @[playground/src/noop/common.scala 330:36]
  wire [63:0] _memAlign_ans_T_4 = alu_out & 64'h7; // @[playground/src/noop/common.scala 331:27]
  wire  _memAlign_ans_T_5 = _memAlign_ans_T_4 == 64'h0; // @[playground/src/noop/common.scala 331:36]
  wire  _memAlign_ans_T_7 = 2'h1 == io_rr2ex_ctrl_dcMode[1:0] ? _memAlign_ans_T_1 : 1'h1; // @[src/main/scala/chisel3/util/Mux.scala 81:58]
  wire  _memAlign_ans_T_9 = 2'h2 == io_rr2ex_ctrl_dcMode[1:0] ? _memAlign_ans_T_3 : _memAlign_ans_T_7; // @[src/main/scala/chisel3/util/Mux.scala 81:58]
  wire  memAlign_ans = 2'h3 == io_rr2ex_ctrl_dcMode[1:0] ? _memAlign_ans_T_5 : _memAlign_ans_T_9; // @[src/main/scala/chisel3/util/Mux.scala 81:58]
  wire  memAlign = io_rr2ex_ctrl_dcMode == 5'h0 | memAlign_ans; // @[playground/src/noop/execute.scala 85:54]
  wire  _T_1 = ~memAlign; // @[playground/src/noop/execute.scala 105:14]
  wire [2:0] _excep_r_cause_T_1 = io_rr2ex_ctrl_dcMode[3] ? 3'h6 : 3'h4; // @[playground/src/noop/execute.scala 108:33]
  wire  _GEN_11 = ~memAlign | io_rr2ex_excep_en; // @[playground/src/noop/execute.scala 105:24 110:25 89:21]
  wire  _GEN_15 = ~memAlign | io_rr2ex_recov; // @[playground/src/noop/execute.scala 101:21 105:24 83:54]
  wire [63:0] _GEN_34 = hs_in ? wdata : dst_d_r; // @[playground/src/noop/execute.scala 86:16 96:21 37:30]
  wire  _GEN_40 = hs_in & _T_1; // @[playground/src/noop/execute.scala 23:12 86:16]
  reg  state; // @[playground/src/noop/execute.scala 118:24]
  reg  drop_alu; // @[playground/src/noop/execute.scala 119:27]
  wire  _T_2 = ~drop_in; // @[playground/src/noop/execute.scala 120:10]
  wire  _GEN_42 = (valid_r | state) & ~hs_out ? 1'h0 : io_rr2ex_valid; // @[playground/src/noop/execute.scala 116:21 121:54]
  wire  _GEN_44 = hs_out ? 1'h0 : valid_r; // @[playground/src/noop/execute.scala 134:31 135:25 44:30]
  wire  _GEN_45 = hs_in | _GEN_44; // @[playground/src/noop/execute.scala 132:30 133:25]
  wire  _GEN_46 = hs_in & ~alu_io_valid ? 1'h0 : _GEN_45; // @[playground/src/noop/execute.scala 129:41 130:25]
  wire  _GEN_47 = hs_in & ~alu_io_valid | state; // @[playground/src/noop/execute.scala 129:41 131:23 118:24]
  wire  _GEN_48 = ~state ? _GEN_46 : valid_r; // @[playground/src/noop/execute.scala 128:30 44:30]
  wire  _GEN_49 = ~state ? _GEN_47 : state; // @[playground/src/noop/execute.scala 118:24 128:30]
  wire  _GEN_52 = alu_io_valid ? ~drop_alu : _GEN_48; // @[playground/src/noop/execute.scala 139:31 142:29]
  wire  _GEN_56 = state ? _GEN_52 : _GEN_48; // @[playground/src/noop/execute.scala 138:33]
  wire  _GEN_58 = state | drop_alu; // @[playground/src/noop/execute.scala 148:30 149:22 119:27]
  wire  _GEN_59 = _io_rr2ex_stall_T & _GEN_56; // @[playground/src/noop/execute.scala 127:26 147:17]
  reg [63:0] forceJmp_seq_pc; // @[playground/src/noop/execute.scala 154:27]
  reg  forceJmp_valid; // @[playground/src/noop/execute.scala 154:27]
  wire  real_is_target = 2'h2 == io_rr2ex_jmp_type ? branchAlu_io_is_jmp : 2'h1 == io_rr2ex_jmp_type; // @[src/main/scala/chisel3/util/Mux.scala 81:58]
  wire  _real_target_T = io_rr2ex_jmp_type == 2'h3; // @[playground/src/noop/execute.scala 164:28]
  wire  _real_target_T_1 = ~real_is_target; // @[playground/src/noop/execute.scala 165:10]
  wire [2:0] _real_target_T_4 = io_rr2ex_inst[1:0] == 2'h3 ? 3'h4 : 3'h2; // @[playground/src/noop/execute.scala 165:62]
  wire [63:0] _GEN_2 = {{61'd0}, _real_target_T_4}; // @[playground/src/noop/execute.scala 165:57]
  wire [63:0] _real_target_T_6 = io_rr2ex_pc + _GEN_2; // @[playground/src/noop/execute.scala 165:57]
  wire  _real_target_T_7 = io_rr2ex_jmp_type == 2'h1; // @[playground/src/noop/execute.scala 166:28]
  wire [63:0] _real_target_T_9 = io_rr2ex_rs1_d + io_rr2ex_dst_d; // @[playground/src/noop/execute.scala 166:60]
  wire [63:0] _real_target_T_10 = _real_target_T_7 ? _real_target_T_9 : io_rr2ex_dst_d; // @[src/main/scala/chisel3/util/Mux.scala 47:70]
  wire [63:0] _real_target_T_11 = _real_target_T_1 ? _real_target_T_6 : _real_target_T_10; // @[src/main/scala/chisel3/util/Mux.scala 47:70]
  wire  _T_18 = hs_in & ~io_rr2ex_excep_en & real_is_target & io_rr2ex_jmp_type != 2'h0; // @[playground/src/noop/execute.scala 174:60]
  wire  _GEN_66 = hs_in & ~io_rr2ex_excep_en & real_is_target & io_rr2ex_jmp_type != 2'h0 | _GEN_40; // @[playground/src/noop/execute.scala 174:92 177:21]
  wire  _GEN_68 = _T_2 & _T_18; // @[playground/src/noop/execute.scala 173:19 155:20]
  wire [1:0] _io_d_ex_state_T_3 = ctrl_r_writeRegEn ? 2'h1 : 2'h0; // @[playground/src/noop/execute.scala 189:91]
  wire [1:0] _io_d_ex_state_T_4 = ctrl_r_dcMode[2] | indi_r[1] ? 2'h2 : _io_d_ex_state_T_3; // @[playground/src/noop/execute.scala 189:31]
  wire [1:0] _GEN_70 = state ? 2'h2 : 2'h0; // @[playground/src/noop/execute.scala 187:20 190:32 191:25]
  ALU alu ( // @[playground/src/noop/execute.scala 27:25]
    .clock(alu_clock),
    .reset(alu_reset),
    .io_alu_op(alu_io_alu_op),
    .io_val1(alu_io_val1),
    .io_val2(alu_io_val2),
    .io_alu64(alu_io_alu64),
    .io_en(alu_io_en),
    .io_out(alu_io_out),
    .io_valid(alu_io_valid)
  );
  BranchALU branchAlu ( // @[playground/src/noop/execute.scala 153:27]
    .io_val1(branchAlu_io_val1),
    .io_val2(branchAlu_io_val2),
    .io_brType(branchAlu_io_brType),
    .io_is_jmp(branchAlu_io_is_jmp)
  );
  assign io_rr2ex_drop = drop_r | io_ex2mem_drop; // @[playground/src/noop/execute.scala 24:26]
  assign io_rr2ex_stall = io_ex2mem_stall | stall_r & ~io_ex2mem_drop; // @[playground/src/noop/execute.scala 26:40]
  assign io_rr2ex_ready = ~drop_in & _GEN_42; // @[playground/src/noop/execute.scala 120:19 116:21]
  assign io_ex2mem_inst = inst_r; // @[playground/src/noop/execute.scala 195:25]
  assign io_ex2mem_pc = pc_r; // @[playground/src/noop/execute.scala 196:25]
  assign io_ex2mem_excep_cause = excep_r_cause; // @[playground/src/noop/execute.scala 197:25]
  assign io_ex2mem_excep_tval = excep_r_tval; // @[playground/src/noop/execute.scala 197:25]
  assign io_ex2mem_excep_en = excep_r_en; // @[playground/src/noop/execute.scala 197:25]
  assign io_ex2mem_excep_pc = excep_r_pc; // @[playground/src/noop/execute.scala 197:25]
  assign io_ex2mem_excep_etype = excep_r_etype; // @[playground/src/noop/execute.scala 197:25]
  assign io_ex2mem_ctrl_dcMode = ctrl_r_dcMode; // @[playground/src/noop/execute.scala 198:25]
  assign io_ex2mem_ctrl_writeRegEn = ctrl_r_writeRegEn; // @[playground/src/noop/execute.scala 198:25]
  assign io_ex2mem_ctrl_writeCSREn = ctrl_r_writeCSREn; // @[playground/src/noop/execute.scala 198:25]
  assign io_ex2mem_mem_addr = mem_addr_r; // @[playground/src/noop/execute.scala 199:25]
  assign io_ex2mem_mem_data = mem_data_r; // @[playground/src/noop/execute.scala 200:25]
  assign io_ex2mem_csr_id = csr_id_r; // @[playground/src/noop/execute.scala 201:25]
  assign io_ex2mem_csr_d = csr_d_r; // @[playground/src/noop/execute.scala 202:25]
  assign io_ex2mem_dst = dst_r; // @[playground/src/noop/execute.scala 203:25]
  assign io_ex2mem_dst_d = dst_d_r; // @[playground/src/noop/execute.scala 204:25]
  assign io_ex2mem_rcsr_id = rcsr_id_r; // @[playground/src/noop/execute.scala 205:25]
  assign io_ex2mem_special = special_r; // @[playground/src/noop/execute.scala 206:25]
  assign io_ex2mem_indi = indi_r; // @[playground/src/noop/execute.scala 207:25]
  assign io_ex2mem_recov = recov_r; // @[playground/src/noop/execute.scala 209:25]
  assign io_ex2mem_valid = valid_r; // @[playground/src/noop/execute.scala 208:25]
  assign io_d_ex_id = dst_r; // @[playground/src/noop/execute.scala 185:20]
  assign io_d_ex_data = dst_d_r; // @[playground/src/noop/execute.scala 186:20]
  assign io_d_ex_state = valid_r ? _io_d_ex_state_T_4 : _GEN_70; // @[playground/src/noop/execute.scala 188:18 189:25]
  assign io_ex2if_seq_pc = forceJmp_seq_pc; // @[playground/src/noop/execute.scala 180:21]
  assign io_ex2if_valid = forceJmp_valid & _io_rr2ex_stall_T; // @[playground/src/noop/execute.scala 181:39]
  assign alu_clock = clock;
  assign alu_reset = reset;
  assign alu_io_alu_op = io_rr2ex_ctrl_aluOp; // @[playground/src/noop/execute.scala 65:21]
  assign alu_io_val1 = unsigned_dr ? _val1_T_1 : _val1_T_7; // @[src/main/scala/chisel3/util/Mux.scala 47:70]
  assign alu_io_val2 = unsigned_dr ? _val2_T_1 : _val2_T_12; // @[src/main/scala/chisel3/util/Mux.scala 47:70]
  assign alu_io_alu64 = ~io_rr2ex_ctrl_aluWidth; // @[playground/src/noop/execute.scala 48:40]
  assign alu_io_en = ~drop_in & _GEN_42; // @[playground/src/noop/execute.scala 120:19 116:21]
  assign branchAlu_io_val1 = unsigned_dr ? _val1_T_1 : _val1_T_7; // @[src/main/scala/chisel3/util/Mux.scala 47:70]
  assign branchAlu_io_val2 = unsigned_dr ? _val2_T_1 : _val2_T_12; // @[src/main/scala/chisel3/util/Mux.scala 47:70]
  assign branchAlu_io_brType = io_rr2ex_ctrl_brType; // @[playground/src/noop/execute.scala 158:25]
  always @(posedge clock) begin
    if (reset) begin // @[playground/src/noop/execute.scala 21:25]
      drop_r <= 1'h0; // @[playground/src/noop/execute.scala 21:25]
    end else if (_T_2) begin // @[playground/src/noop/execute.scala 173:19]
      drop_r <= _GEN_66;
    end else begin
      drop_r <= _GEN_40;
    end
    if (reset) begin // @[playground/src/noop/execute.scala 22:26]
      stall_r <= 1'h0; // @[playground/src/noop/execute.scala 22:26]
    end else begin
      stall_r <= _GEN_40;
    end
    if (reset) begin // @[playground/src/noop/execute.scala 28:30]
      inst_r <= 32'h0; // @[playground/src/noop/execute.scala 28:30]
    end else if (hs_in) begin // @[playground/src/noop/execute.scala 86:16]
      inst_r <= io_rr2ex_inst; // @[playground/src/noop/execute.scala 87:21]
    end
    if (reset) begin // @[playground/src/noop/execute.scala 29:30]
      pc_r <= 64'h0; // @[playground/src/noop/execute.scala 29:30]
    end else if (hs_in) begin // @[playground/src/noop/execute.scala 86:16]
      pc_r <= io_rr2ex_pc; // @[playground/src/noop/execute.scala 88:21]
    end
    if (reset) begin // @[playground/src/noop/execute.scala 30:30]
      excep_r_cause <= 64'h0; // @[playground/src/noop/execute.scala 30:30]
    end else if (hs_in) begin // @[playground/src/noop/execute.scala 86:16]
      if (~memAlign) begin // @[playground/src/noop/execute.scala 105:24]
        excep_r_cause <= {{61'd0}, _excep_r_cause_T_1}; // @[playground/src/noop/execute.scala 108:27]
      end else begin
        excep_r_cause <= io_rr2ex_excep_cause; // @[playground/src/noop/execute.scala 89:21]
      end
    end
    if (reset) begin // @[playground/src/noop/execute.scala 30:30]
      excep_r_tval <= 64'h0; // @[playground/src/noop/execute.scala 30:30]
    end else if (hs_in) begin // @[playground/src/noop/execute.scala 86:16]
      if (~memAlign) begin // @[playground/src/noop/execute.scala 105:24]
        if (cur_alu64) begin // @[playground/src/noop/execute.scala 71:22]
          excep_r_tval <= _alu_out_T;
        end else begin
          excep_r_tval <= _alu_out_T_5;
        end
      end else begin
        excep_r_tval <= io_rr2ex_excep_tval; // @[playground/src/noop/execute.scala 89:21]
      end
    end
    if (reset) begin // @[playground/src/noop/execute.scala 30:30]
      excep_r_en <= 1'h0; // @[playground/src/noop/execute.scala 30:30]
    end else if (hs_in) begin // @[playground/src/noop/execute.scala 86:16]
      excep_r_en <= _GEN_11;
    end
    if (reset) begin // @[playground/src/noop/execute.scala 30:30]
      excep_r_pc <= 64'h0; // @[playground/src/noop/execute.scala 30:30]
    end else if (hs_in) begin // @[playground/src/noop/execute.scala 86:16]
      if (~memAlign) begin // @[playground/src/noop/execute.scala 105:24]
        excep_r_pc <= io_rr2ex_pc; // @[playground/src/noop/execute.scala 111:25]
      end else if (io_rr2ex_excep_cause[63]) begin // @[playground/src/noop/execute.scala 102:39]
        excep_r_pc <= next_pc_r; // @[playground/src/noop/execute.scala 103:24]
      end else begin
        excep_r_pc <= io_rr2ex_excep_pc; // @[playground/src/noop/execute.scala 89:21]
      end
    end
    if (reset) begin // @[playground/src/noop/execute.scala 30:30]
      excep_r_etype <= 2'h0; // @[playground/src/noop/execute.scala 30:30]
    end else if (hs_in) begin // @[playground/src/noop/execute.scala 86:16]
      if (~memAlign) begin // @[playground/src/noop/execute.scala 105:24]
        excep_r_etype <= 2'h0; // @[playground/src/noop/execute.scala 112:27]
      end else begin
        excep_r_etype <= io_rr2ex_excep_etype; // @[playground/src/noop/execute.scala 89:21]
      end
    end
    if (reset) begin // @[playground/src/noop/execute.scala 31:30]
      ctrl_r_dcMode <= 5'h0; // @[playground/src/noop/execute.scala 31:30]
    end else if (hs_in) begin // @[playground/src/noop/execute.scala 86:16]
      if (~memAlign) begin // @[playground/src/noop/execute.scala 105:24]
        ctrl_r_dcMode <= 5'h0; // @[playground/src/noop/execute.scala 106:20]
      end else begin
        ctrl_r_dcMode <= io_rr2ex_ctrl_dcMode; // @[playground/src/noop/execute.scala 90:21]
      end
    end
    if (reset) begin // @[playground/src/noop/execute.scala 31:30]
      ctrl_r_writeRegEn <= 1'h0; // @[playground/src/noop/execute.scala 31:30]
    end else if (hs_in) begin // @[playground/src/noop/execute.scala 86:16]
      if (~memAlign) begin // @[playground/src/noop/execute.scala 105:24]
        ctrl_r_writeRegEn <= 1'h0; // @[playground/src/noop/execute.scala 106:20]
      end else begin
        ctrl_r_writeRegEn <= io_rr2ex_ctrl_writeRegEn; // @[playground/src/noop/execute.scala 90:21]
      end
    end
    if (reset) begin // @[playground/src/noop/execute.scala 31:30]
      ctrl_r_writeCSREn <= 1'h0; // @[playground/src/noop/execute.scala 31:30]
    end else if (hs_in) begin // @[playground/src/noop/execute.scala 86:16]
      if (~memAlign) begin // @[playground/src/noop/execute.scala 105:24]
        ctrl_r_writeCSREn <= 1'h0; // @[playground/src/noop/execute.scala 106:20]
      end else begin
        ctrl_r_writeCSREn <= io_rr2ex_ctrl_writeCSREn; // @[playground/src/noop/execute.scala 90:21]
      end
    end
    if (reset) begin // @[playground/src/noop/execute.scala 32:30]
      mem_addr_r <= 64'h0; // @[playground/src/noop/execute.scala 32:30]
    end else if (hs_in) begin // @[playground/src/noop/execute.scala 86:16]
      if (cur_alu64) begin // @[playground/src/noop/execute.scala 71:22]
        mem_addr_r <= _alu_out_T;
      end else begin
        mem_addr_r <= _alu_out_T_5;
      end
    end
    if (reset) begin // @[playground/src/noop/execute.scala 33:30]
      mem_data_r <= 64'h0; // @[playground/src/noop/execute.scala 33:30]
    end else if (hs_in) begin // @[playground/src/noop/execute.scala 86:16]
      if (io_rr2ex_ctrl_dcMode[3]) begin // @[src/main/scala/chisel3/util/Mux.scala 47:70]
        mem_data_r <= io_rr2ex_dst_d;
      end else if (io_rr2ex_ctrl_writeCSREn) begin // @[src/main/scala/chisel3/util/Mux.scala 47:70]
        mem_data_r <= io_rr2ex_rs2_d;
      end else begin
        mem_data_r <= alu_out;
      end
    end
    if (reset) begin // @[playground/src/noop/execute.scala 34:30]
      csr_id_r <= 12'h0; // @[playground/src/noop/execute.scala 34:30]
    end else if (hs_in) begin // @[playground/src/noop/execute.scala 86:16]
      csr_id_r <= io_rr2ex_rs2; // @[playground/src/noop/execute.scala 93:21]
    end
    if (reset) begin // @[playground/src/noop/execute.scala 35:30]
      csr_d_r <= 64'h0; // @[playground/src/noop/execute.scala 35:30]
    end else if (hs_in) begin // @[playground/src/noop/execute.scala 86:16]
      if (cur_alu64) begin // @[playground/src/noop/execute.scala 71:22]
        csr_d_r <= _alu_out_T;
      end else begin
        csr_d_r <= _alu_out_T_5;
      end
    end
    if (reset) begin // @[playground/src/noop/execute.scala 36:30]
      dst_r <= 5'h0; // @[playground/src/noop/execute.scala 36:30]
    end else if (hs_in) begin // @[playground/src/noop/execute.scala 86:16]
      dst_r <= io_rr2ex_dst; // @[playground/src/noop/execute.scala 95:21]
    end
    if (reset) begin // @[playground/src/noop/execute.scala 37:30]
      dst_d_r <= 64'h0; // @[playground/src/noop/execute.scala 37:30]
    end else if (_io_rr2ex_stall_T) begin // @[playground/src/noop/execute.scala 127:26]
      if (state) begin // @[playground/src/noop/execute.scala 138:33]
        if (alu_io_valid) begin // @[playground/src/noop/execute.scala 139:31]
          dst_d_r <= alu_out; // @[playground/src/noop/execute.scala 141:29]
        end else begin
          dst_d_r <= _GEN_34;
        end
      end else begin
        dst_d_r <= _GEN_34;
      end
    end else begin
      dst_d_r <= _GEN_34;
    end
    if (reset) begin // @[playground/src/noop/execute.scala 38:30]
      rcsr_id_r <= 12'h0; // @[playground/src/noop/execute.scala 38:30]
    end else if (hs_in) begin // @[playground/src/noop/execute.scala 86:16]
      rcsr_id_r <= io_rr2ex_rcsr_id; // @[playground/src/noop/execute.scala 97:21]
    end
    if (reset) begin // @[playground/src/noop/execute.scala 39:30]
      special_r <= 2'h0; // @[playground/src/noop/execute.scala 39:30]
    end else if (hs_in) begin // @[playground/src/noop/execute.scala 86:16]
      special_r <= io_rr2ex_special; // @[playground/src/noop/execute.scala 98:21]
    end
    if (reset) begin // @[playground/src/noop/execute.scala 40:30]
      alu64_r <= 1'h0; // @[playground/src/noop/execute.scala 40:30]
    end else if (hs_in) begin // @[playground/src/noop/execute.scala 70:26]
      alu64_r <= alu64;
    end
    if (reset) begin // @[playground/src/noop/execute.scala 41:30]
      indi_r <= 2'h0; // @[playground/src/noop/execute.scala 41:30]
    end else if (hs_in) begin // @[playground/src/noop/execute.scala 86:16]
      if (~memAlign) begin // @[playground/src/noop/execute.scala 105:24]
        indi_r <= 2'h0; // @[playground/src/noop/execute.scala 107:20]
      end else begin
        indi_r <= io_rr2ex_indi; // @[playground/src/noop/execute.scala 99:21]
      end
    end
    if (reset) begin // @[playground/src/noop/execute.scala 42:30]
      next_pc_r <= 64'h0; // @[playground/src/noop/execute.scala 42:30]
    end else if (hs_in) begin // @[playground/src/noop/execute.scala 170:16]
      if (_real_target_T) begin // @[src/main/scala/chisel3/util/Mux.scala 47:70]
        next_pc_r <= io_rr2ex_rs2_d;
      end else if (_real_target_T_1) begin // @[src/main/scala/chisel3/util/Mux.scala 47:70]
        next_pc_r <= _real_target_T_6;
      end else begin
        next_pc_r <= _real_target_T_10;
      end
    end else if (io_updateNextPc_valid) begin // @[playground/src/noop/execute.scala 78:32]
      next_pc_r <= io_updateNextPc_seq_pc; // @[playground/src/noop/execute.scala 79:19]
    end
    if (reset) begin // @[playground/src/noop/execute.scala 43:30]
      recov_r <= 1'h0; // @[playground/src/noop/execute.scala 43:30]
    end else if (hs_in) begin // @[playground/src/noop/execute.scala 86:16]
      recov_r <= _GEN_15;
    end
    if (reset) begin // @[playground/src/noop/execute.scala 44:30]
      valid_r <= 1'h0; // @[playground/src/noop/execute.scala 44:30]
    end else begin
      valid_r <= _GEN_59;
    end
    if (reset) begin // @[playground/src/noop/execute.scala 118:24]
      state <= 1'h0; // @[playground/src/noop/execute.scala 118:24]
    end else if (_io_rr2ex_stall_T) begin // @[playground/src/noop/execute.scala 127:26]
      if (state) begin // @[playground/src/noop/execute.scala 138:33]
        if (alu_io_valid) begin // @[playground/src/noop/execute.scala 139:31]
          state <= 1'h0; // @[playground/src/noop/execute.scala 140:29]
        end else begin
          state <= _GEN_49;
        end
      end else begin
        state <= _GEN_49;
      end
    end
    if (reset) begin // @[playground/src/noop/execute.scala 119:27]
      drop_alu <= 1'h0; // @[playground/src/noop/execute.scala 119:27]
    end else if (_io_rr2ex_stall_T) begin // @[playground/src/noop/execute.scala 127:26]
      if (state) begin // @[playground/src/noop/execute.scala 138:33]
        if (alu_io_valid) begin // @[playground/src/noop/execute.scala 139:31]
          drop_alu <= 1'h0; // @[playground/src/noop/execute.scala 143:29]
        end
      end
    end else begin
      drop_alu <= _GEN_58;
    end
    if (reset) begin // @[playground/src/noop/execute.scala 154:27]
      forceJmp_seq_pc <= 64'h0; // @[playground/src/noop/execute.scala 154:27]
    end else if (_T_2) begin // @[playground/src/noop/execute.scala 173:19]
      if (hs_in & ~io_rr2ex_excep_en & real_is_target & io_rr2ex_jmp_type != 2'h0) begin // @[playground/src/noop/execute.scala 174:92]
        if (_real_target_T) begin // @[src/main/scala/chisel3/util/Mux.scala 47:70]
          forceJmp_seq_pc <= io_rr2ex_rs2_d;
        end else begin
          forceJmp_seq_pc <= _real_target_T_11;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/execute.scala 154:27]
      forceJmp_valid <= 1'h0; // @[playground/src/noop/execute.scala 154:27]
    end else begin
      forceJmp_valid <= _GEN_68;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  drop_r = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  stall_r = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  inst_r = _RAND_2[31:0];
  _RAND_3 = {2{`RANDOM}};
  pc_r = _RAND_3[63:0];
  _RAND_4 = {2{`RANDOM}};
  excep_r_cause = _RAND_4[63:0];
  _RAND_5 = {2{`RANDOM}};
  excep_r_tval = _RAND_5[63:0];
  _RAND_6 = {1{`RANDOM}};
  excep_r_en = _RAND_6[0:0];
  _RAND_7 = {2{`RANDOM}};
  excep_r_pc = _RAND_7[63:0];
  _RAND_8 = {1{`RANDOM}};
  excep_r_etype = _RAND_8[1:0];
  _RAND_9 = {1{`RANDOM}};
  ctrl_r_dcMode = _RAND_9[4:0];
  _RAND_10 = {1{`RANDOM}};
  ctrl_r_writeRegEn = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  ctrl_r_writeCSREn = _RAND_11[0:0];
  _RAND_12 = {2{`RANDOM}};
  mem_addr_r = _RAND_12[63:0];
  _RAND_13 = {2{`RANDOM}};
  mem_data_r = _RAND_13[63:0];
  _RAND_14 = {1{`RANDOM}};
  csr_id_r = _RAND_14[11:0];
  _RAND_15 = {2{`RANDOM}};
  csr_d_r = _RAND_15[63:0];
  _RAND_16 = {1{`RANDOM}};
  dst_r = _RAND_16[4:0];
  _RAND_17 = {2{`RANDOM}};
  dst_d_r = _RAND_17[63:0];
  _RAND_18 = {1{`RANDOM}};
  rcsr_id_r = _RAND_18[11:0];
  _RAND_19 = {1{`RANDOM}};
  special_r = _RAND_19[1:0];
  _RAND_20 = {1{`RANDOM}};
  alu64_r = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  indi_r = _RAND_21[1:0];
  _RAND_22 = {2{`RANDOM}};
  next_pc_r = _RAND_22[63:0];
  _RAND_23 = {1{`RANDOM}};
  recov_r = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  valid_r = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  state = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  drop_alu = _RAND_26[0:0];
  _RAND_27 = {2{`RANDOM}};
  forceJmp_seq_pc = _RAND_27[63:0];
  _RAND_28 = {1{`RANDOM}};
  forceJmp_valid = _RAND_28[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Memory(
  input         clock,
  input         reset,
  input  [31:0] io_ex2mem_inst, // @[playground/src/noop/memory.scala 85:16]
  input  [63:0] io_ex2mem_pc, // @[playground/src/noop/memory.scala 85:16]
  input  [63:0] io_ex2mem_excep_cause, // @[playground/src/noop/memory.scala 85:16]
  input  [63:0] io_ex2mem_excep_tval, // @[playground/src/noop/memory.scala 85:16]
  input         io_ex2mem_excep_en, // @[playground/src/noop/memory.scala 85:16]
  input  [63:0] io_ex2mem_excep_pc, // @[playground/src/noop/memory.scala 85:16]
  input  [1:0]  io_ex2mem_excep_etype, // @[playground/src/noop/memory.scala 85:16]
  input  [4:0]  io_ex2mem_ctrl_dcMode, // @[playground/src/noop/memory.scala 85:16]
  input         io_ex2mem_ctrl_writeRegEn, // @[playground/src/noop/memory.scala 85:16]
  input         io_ex2mem_ctrl_writeCSREn, // @[playground/src/noop/memory.scala 85:16]
  input  [63:0] io_ex2mem_mem_addr, // @[playground/src/noop/memory.scala 85:16]
  input  [63:0] io_ex2mem_mem_data, // @[playground/src/noop/memory.scala 85:16]
  input  [11:0] io_ex2mem_csr_id, // @[playground/src/noop/memory.scala 85:16]
  input  [63:0] io_ex2mem_csr_d, // @[playground/src/noop/memory.scala 85:16]
  input  [4:0]  io_ex2mem_dst, // @[playground/src/noop/memory.scala 85:16]
  input  [63:0] io_ex2mem_dst_d, // @[playground/src/noop/memory.scala 85:16]
  input  [11:0] io_ex2mem_rcsr_id, // @[playground/src/noop/memory.scala 85:16]
  input  [1:0]  io_ex2mem_special, // @[playground/src/noop/memory.scala 85:16]
  input  [1:0]  io_ex2mem_indi, // @[playground/src/noop/memory.scala 85:16]
  output        io_ex2mem_drop, // @[playground/src/noop/memory.scala 85:16]
  output        io_ex2mem_stall, // @[playground/src/noop/memory.scala 85:16]
  input         io_ex2mem_recov, // @[playground/src/noop/memory.scala 85:16]
  input         io_ex2mem_valid, // @[playground/src/noop/memory.scala 85:16]
  output        io_ex2mem_ready, // @[playground/src/noop/memory.scala 85:16]
  output [31:0] io_mem2rb_inst, // @[playground/src/noop/memory.scala 85:16]
  output [63:0] io_mem2rb_pc, // @[playground/src/noop/memory.scala 85:16]
  output [63:0] io_mem2rb_excep_cause, // @[playground/src/noop/memory.scala 85:16]
  output [63:0] io_mem2rb_excep_tval, // @[playground/src/noop/memory.scala 85:16]
  output        io_mem2rb_excep_en, // @[playground/src/noop/memory.scala 85:16]
  output [63:0] io_mem2rb_excep_pc, // @[playground/src/noop/memory.scala 85:16]
  output [1:0]  io_mem2rb_excep_etype, // @[playground/src/noop/memory.scala 85:16]
  output [11:0] io_mem2rb_csr_id, // @[playground/src/noop/memory.scala 85:16]
  output [63:0] io_mem2rb_csr_d, // @[playground/src/noop/memory.scala 85:16]
  output        io_mem2rb_csr_en, // @[playground/src/noop/memory.scala 85:16]
  output [4:0]  io_mem2rb_dst, // @[playground/src/noop/memory.scala 85:16]
  output [63:0] io_mem2rb_dst_d, // @[playground/src/noop/memory.scala 85:16]
  output        io_mem2rb_dst_en, // @[playground/src/noop/memory.scala 85:16]
  output [11:0] io_mem2rb_rcsr_id, // @[playground/src/noop/memory.scala 85:16]
  output [1:0]  io_mem2rb_special, // @[playground/src/noop/memory.scala 85:16]
  output        io_mem2rb_is_mmio, // @[playground/src/noop/memory.scala 85:16]
  input         io_mem2rb_drop, // @[playground/src/noop/memory.scala 85:16]
  input         io_mem2rb_stall, // @[playground/src/noop/memory.scala 85:16]
  output        io_mem2rb_recov, // @[playground/src/noop/memory.scala 85:16]
  output        io_mem2rb_valid, // @[playground/src/noop/memory.scala 85:16]
  input         io_mem2rb_ready, // @[playground/src/noop/memory.scala 85:16]
  output [31:0] io_dataRW_addr, // @[playground/src/noop/memory.scala 85:16]
  input  [63:0] io_dataRW_rdata, // @[playground/src/noop/memory.scala 85:16]
  input         io_dataRW_rvalid, // @[playground/src/noop/memory.scala 85:16]
  output [63:0] io_dataRW_wdata, // @[playground/src/noop/memory.scala 85:16]
  output [4:0]  io_dataRW_dc_mode, // @[playground/src/noop/memory.scala 85:16]
  output [4:0]  io_dataRW_amo, // @[playground/src/noop/memory.scala 85:16]
  input         io_dataRW_ready, // @[playground/src/noop/memory.scala 85:16]
  output [63:0] io_va2pa_vaddr, // @[playground/src/noop/memory.scala 85:16]
  output        io_va2pa_vvalid, // @[playground/src/noop/memory.scala 85:16]
  output [1:0]  io_va2pa_m_type, // @[playground/src/noop/memory.scala 85:16]
  input  [31:0] io_va2pa_paddr, // @[playground/src/noop/memory.scala 85:16]
  input         io_va2pa_pvalid, // @[playground/src/noop/memory.scala 85:16]
  input  [63:0] io_va2pa_tlb_excep_cause, // @[playground/src/noop/memory.scala 85:16]
  input  [63:0] io_va2pa_tlb_excep_tval, // @[playground/src/noop/memory.scala 85:16]
  input         io_va2pa_tlb_excep_en, // @[playground/src/noop/memory.scala 85:16]
  output [4:0]  io_d_mem1_id, // @[playground/src/noop/memory.scala 85:16]
  output [63:0] io_d_mem1_data, // @[playground/src/noop/memory.scala 85:16]
  output [1:0]  io_d_mem1_state, // @[playground/src/noop/memory.scala 85:16]
  output [4:0]  io_d_mem2_id, // @[playground/src/noop/memory.scala 85:16]
  output [63:0] io_d_mem2_data, // @[playground/src/noop/memory.scala 85:16]
  output [1:0]  io_d_mem2_state, // @[playground/src/noop/memory.scala 85:16]
  output [4:0]  io_d_mem3_id, // @[playground/src/noop/memory.scala 85:16]
  output [63:0] io_d_mem3_data, // @[playground/src/noop/memory.scala 85:16]
  output [1:0]  io_d_mem3_state // @[playground/src/noop/memory.scala 85:16]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [63:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [63:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [63:0] _RAND_30;
  reg [63:0] _RAND_31;
  reg [63:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [63:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [63:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [63:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [63:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [63:0] _RAND_51;
  reg [63:0] _RAND_52;
  reg [63:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [63:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [63:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [63:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
`endif // RANDOMIZE_REG_INIT
  reg  drop2_r; // @[playground/src/noop/memory.scala 95:26]
  reg  stall2_r; // @[playground/src/noop/memory.scala 98:27]
  wire  drop2_in = drop2_r | io_mem2rb_drop; // @[playground/src/noop/memory.scala 103:31]
  wire  _stall3_in_T = ~io_mem2rb_drop; // @[playground/src/noop/memory.scala 105:34]
  wire  _stall1_in_T = ~drop2_in; // @[playground/src/noop/memory.scala 107:34]
  reg [31:0] inst1_r; // @[playground/src/noop/memory.scala 111:30]
  reg [63:0] pc1_r; // @[playground/src/noop/memory.scala 112:30]
  reg [63:0] excep1_r_cause; // @[playground/src/noop/memory.scala 113:30]
  reg [63:0] excep1_r_tval; // @[playground/src/noop/memory.scala 113:30]
  reg  excep1_r_en; // @[playground/src/noop/memory.scala 113:30]
  reg [63:0] excep1_r_pc; // @[playground/src/noop/memory.scala 113:30]
  reg [1:0] excep1_r_etype; // @[playground/src/noop/memory.scala 113:30]
  reg [4:0] ctrl1_r_dcMode; // @[playground/src/noop/memory.scala 114:30]
  reg [63:0] mem_addr1_r; // @[playground/src/noop/memory.scala 115:30]
  reg [63:0] mem_data1_r; // @[playground/src/noop/memory.scala 116:30]
  reg [4:0] dst1_r; // @[playground/src/noop/memory.scala 117:30]
  reg [63:0] dst_d1_r; // @[playground/src/noop/memory.scala 118:30]
  reg  dst_en1_r; // @[playground/src/noop/memory.scala 119:30]
  reg [11:0] csr_id1_r; // @[playground/src/noop/memory.scala 120:30]
  reg [63:0] csr_d1_r; // @[playground/src/noop/memory.scala 121:30]
  reg  csr_en1_r; // @[playground/src/noop/memory.scala 122:30]
  reg [11:0] rcsr_id1_r; // @[playground/src/noop/memory.scala 123:30]
  reg [1:0] special1_r; // @[playground/src/noop/memory.scala 124:30]
  reg [1:0] indi1_r; // @[playground/src/noop/memory.scala 125:30]
  reg  recov1_r; // @[playground/src/noop/memory.scala 126:30]
  reg  valid1_r; // @[playground/src/noop/memory.scala 128:30]
  reg  is_tlb_r; // @[playground/src/noop/memory.scala 134:30]
  reg  drop_tlb; // @[playground/src/noop/memory.scala 135:30]
  wire  hs_in = io_ex2mem_ready & io_ex2mem_valid; // @[playground/src/noop/memory.scala 137:35]
  wire [4:0] _GEN_9 = hs_in ? io_ex2mem_ctrl_dcMode : ctrl1_r_dcMode; // @[playground/src/noop/memory.scala 142:16 146:21 114:30]
  wire  access_tlb = io_ex2mem_ctrl_dcMode != 5'h0; // @[playground/src/noop/memory.scala 160:45]
  reg  valid2_r; // @[playground/src/noop/memory.scala 214:30]
  reg  valid3_r; // @[playground/src/noop/memory.scala 343:30]
  reg [4:0] ctrl2_r_dcMode; // @[playground/src/noop/memory.scala 201:30]
  wire  is_dc_r = ctrl2_r_dcMode != 5'h0; // @[playground/src/noop/memory.scala 254:39]
  wire  _dc_valid3_T = ~is_dc_r; // @[playground/src/noop/memory.scala 367:21]
  reg  drop_dc; // @[playground/src/noop/memory.scala 255:30]
  wire  dc_valid3 = ~is_dc_r | io_dataRW_rvalid & ~drop_dc; // @[playground/src/noop/memory.scala 367:30]
  wire  _T_34 = valid2_r & dc_valid3; // @[playground/src/noop/memory.scala 370:29]
  wire  _GEN_167 = valid3_r & ~io_mem2rb_ready ? 1'h0 : _T_34; // @[playground/src/noop/memory.scala 141:25 369:34]
  wire  hs2 = _stall3_in_T & _GEN_167; // @[playground/src/noop/memory.scala 368:20 141:25]
  wire  inp_tlb_valid2 = io_va2pa_pvalid | io_va2pa_tlb_excep_en; // @[playground/src/noop/memory.scala 260:42]
  wire  _tlb_valid2_T_1 = ~drop_tlb; // @[playground/src/noop/memory.scala 282:55]
  wire  tlb_valid2 = ~is_tlb_r | inp_tlb_valid2 & ~drop_tlb; // @[playground/src/noop/memory.scala 282:33]
  wire  _T_23 = valid1_r & tlb_valid2; // @[playground/src/noop/memory.scala 289:29]
  wire  _GEN_89 = valid2_r & ~hs2 ? 1'h0 : _T_23; // @[playground/src/noop/memory.scala 288:31 141:9]
  wire  hs1 = _stall1_in_T & _GEN_89; // @[playground/src/noop/memory.scala 287:20 141:9]
  wire  _io_va2pa_vvalid_T_2 = ~hs1; // @[playground/src/noop/memory.scala 162:49]
  wire  _GEN_26 = valid1_r & _io_va2pa_vvalid_T_2 ? 1'h0 : io_ex2mem_valid; // @[playground/src/noop/memory.scala 165:21 167:31]
  wire  _GEN_28 = hs1 ? 1'h0 : valid1_r; // @[playground/src/noop/memory.scala 177:24 178:22 128:30]
  wire  _GEN_29 = hs1 ? 1'h0 : is_tlb_r; // @[playground/src/noop/memory.scala 177:24 179:22 134:30]
  wire  _GEN_30 = hs_in | _GEN_28; // @[playground/src/noop/memory.scala 173:20 174:22]
  wire  _GEN_31 = hs_in ? access_tlb : _GEN_29; // @[playground/src/noop/memory.scala 173:20 175:22]
  wire  _GEN_32 = hs_in ? access_tlb : _stall1_in_T & is_tlb_r & ~hs1; // @[playground/src/noop/memory.scala 173:20 162:21 176:29]
  wire  _GEN_33 = _stall1_in_T & _GEN_30; // @[playground/src/noop/memory.scala 172:20 182:18]
  wire  _GEN_34 = _stall1_in_T & _GEN_31; // @[playground/src/noop/memory.scala 172:20 184:18]
  wire [1:0] _GEN_37 = valid1_r ? 2'h2 : 2'h0; // @[playground/src/noop/memory.scala 192:25 193:25 195:25]
  wire [1:0] _GEN_38 = valid1_r & ~(ctrl1_r_dcMode[2] | indi1_r[1]) ? 2'h1 : _GEN_37; // @[playground/src/noop/memory.scala 190:80 191:25]
  reg [31:0] inst2_r; // @[playground/src/noop/memory.scala 198:30]
  reg [63:0] pc2_r; // @[playground/src/noop/memory.scala 199:30]
  reg [63:0] excep2_r_cause; // @[playground/src/noop/memory.scala 200:30]
  reg [63:0] excep2_r_tval; // @[playground/src/noop/memory.scala 200:30]
  reg  excep2_r_en; // @[playground/src/noop/memory.scala 200:30]
  reg [63:0] excep2_r_pc; // @[playground/src/noop/memory.scala 200:30]
  reg [1:0] excep2_r_etype; // @[playground/src/noop/memory.scala 200:30]
  reg [63:0] mem_data2_r; // @[playground/src/noop/memory.scala 202:30]
  reg [4:0] dst2_r; // @[playground/src/noop/memory.scala 203:30]
  reg [63:0] dst_d2_r; // @[playground/src/noop/memory.scala 204:30]
  reg  dst_en2_r; // @[playground/src/noop/memory.scala 205:30]
  reg [11:0] csr_id2_r; // @[playground/src/noop/memory.scala 206:30]
  reg [63:0] csr_d2_r; // @[playground/src/noop/memory.scala 207:30]
  reg  csr_en2_r; // @[playground/src/noop/memory.scala 208:30]
  reg [11:0] rcsr_id2_r; // @[playground/src/noop/memory.scala 209:30]
  reg [1:0] special2_r; // @[playground/src/noop/memory.scala 210:30]
  reg [31:0] paddr2_r; // @[playground/src/noop/memory.scala 211:30]
  reg  recov2_r; // @[playground/src/noop/memory.scala 213:30]
  reg  dc_hs_r; // @[playground/src/noop/memory.scala 215:30]
  reg [31:0] lr_addr_r; // @[playground/src/noop/memory.scala 217:30]
  reg  lr_valid_r; // @[playground/src/noop/memory.scala 218:30]
  wire  stage2_is_excep = excep1_r_en | io_va2pa_tlb_excep_en; // @[playground/src/noop/memory.scala 227:39]
  wire  _GEN_41 = indi1_r[0] & ~stage2_is_excep | lr_valid_r; // @[playground/src/noop/memory.scala 245:55 246:25 218:30]
  wire [63:0] _GEN_46 = hs1 ? excep1_r_cause : excep2_r_cause; // @[playground/src/noop/memory.scala 228:14 231:21 200:30]
  wire [63:0] _GEN_47 = hs1 ? excep1_r_tval : excep2_r_tval; // @[playground/src/noop/memory.scala 228:14 231:21 200:30]
  wire  _GEN_48 = hs1 ? excep1_r_en : excep2_r_en; // @[playground/src/noop/memory.scala 228:14 231:21 200:30]
  wire [63:0] _GEN_49 = hs1 ? excep1_r_pc : excep2_r_pc; // @[playground/src/noop/memory.scala 228:14 231:21 200:30]
  wire [1:0] _GEN_50 = hs1 ? excep1_r_etype : excep2_r_etype; // @[playground/src/noop/memory.scala 228:14 231:21 200:30]
  wire [4:0] _GEN_54 = hs1 ? ctrl1_r_dcMode : ctrl2_r_dcMode; // @[playground/src/noop/memory.scala 228:14 233:21 201:30]
  wire [63:0] _GEN_59 = hs1 ? dst_d1_r : dst_d2_r; // @[playground/src/noop/memory.scala 228:14 235:21 204:30]
  wire  _GEN_60 = hs1 ? dst_en1_r : dst_en2_r; // @[playground/src/noop/memory.scala 228:14 236:21 205:30]
  wire  _GEN_63 = hs1 ? csr_en1_r : csr_en2_r; // @[playground/src/noop/memory.scala 228:14 239:21 208:30]
  wire  _GEN_67 = hs1 ? recov1_r : recov2_r; // @[playground/src/noop/memory.scala 228:14 243:21 213:30]
  wire  sc_valid = io_va2pa_paddr == lr_addr_r & lr_valid_r; // @[playground/src/noop/memory.scala 261:52]
  wire [4:0] _GEN_71 = indi1_r[1] ? 5'h0 : ctrl1_r_dcMode; // @[playground/src/noop/memory.scala 270:41 271:31 276:31]
  wire [4:0] _GEN_72 = indi1_r[1] ? 5'h0 : _GEN_54; // @[playground/src/noop/memory.scala 270:41 272:29]
  wire  _GEN_73 = indi1_r[1] | _GEN_60; // @[playground/src/noop/memory.scala 270:41 273:25]
  wire [63:0] _GEN_74 = indi1_r[1] ? 64'h1 : _GEN_59; // @[playground/src/noop/memory.scala 270:41 274:25]
  wire [4:0] _GEN_75 = indi1_r[1] & sc_valid ? ctrl1_r_dcMode : _GEN_71; // @[playground/src/noop/memory.scala 266:53 267:31]
  wire  _GEN_76 = indi1_r[1] & sc_valid | _GEN_73; // @[playground/src/noop/memory.scala 266:53 268:25]
  wire [4:0] _GEN_78 = indi1_r[1] & sc_valid ? _GEN_54 : _GEN_72; // @[playground/src/noop/memory.scala 266:53]
  wire [4:0] _GEN_79 = stage2_is_excep ? 5'h0 : _GEN_75; // @[playground/src/noop/memory.scala 263:30 264:31]
  wire [4:0] _GEN_80 = stage2_is_excep ? 5'h0 : _GEN_78; // @[playground/src/noop/memory.scala 263:30 265:29]
  wire  _GEN_81 = stage2_is_excep ? _GEN_60 : _GEN_76; // @[playground/src/noop/memory.scala 263:30]
  wire [4:0] _io_dataRW_dc_mode_T_2 = valid2_r & ~dc_hs_r ? ctrl2_r_dcMode : 5'h0; // @[playground/src/noop/memory.scala 279:33]
  wire [4:0] _GEN_84 = hs1 ? _GEN_80 : _GEN_54; // @[playground/src/noop/memory.scala 262:14]
  wire  _GEN_85 = hs1 ? _GEN_81 : _GEN_60; // @[playground/src/noop/memory.scala 262:14]
  wire  dc_hs = io_dataRW_dc_mode != 5'h0 & io_dataRW_ready; // @[playground/src/noop/memory.scala 283:48]
  wire  _GEN_87 = dc_hs | dc_hs_r; // @[playground/src/noop/memory.scala 284:16 285:17 215:30]
  wire  _T_26 = io_va2pa_tlb_excep_en & _tlb_valid2_T_1; // @[playground/src/noop/memory.scala 296:40]
  wire  _GEN_91 = ctrl1_r_dcMode != 5'h0 ? dc_hs : _GEN_87; // @[playground/src/noop/memory.scala 306:52 307:25]
  wire  _GEN_94 = io_va2pa_tlb_excep_en & _tlb_valid2_T_1 | _GEN_48; // @[playground/src/noop/memory.scala 296:53 299:33]
  wire  _GEN_106 = io_va2pa_tlb_excep_en & _tlb_valid2_T_1 | _GEN_67; // @[playground/src/noop/memory.scala 296:53 221:57]
  wire  _GEN_108 = hs2 ? 1'h0 : valid2_r; // @[playground/src/noop/memory.scala 309:24 310:22 214:30]
  wire  _GEN_110 = hs1 | _GEN_108; // @[playground/src/noop/memory.scala 294:18 295:22]
  wire  _GEN_124 = hs1 & _T_26; // @[playground/src/noop/memory.scala 100:13 294:18]
  wire  _GEN_127 = _stall3_in_T & _GEN_110; // @[playground/src/noop/memory.scala 293:20 314:18]
  wire  _GEN_141 = _stall3_in_T & _GEN_124; // @[playground/src/noop/memory.scala 100:13 293:20]
  wire [1:0] _GEN_145 = valid2_r ? 2'h2 : 2'h0; // @[playground/src/noop/memory.scala 324:25 325:25 327:25]
  wire [1:0] _GEN_146 = valid2_r & _dc_valid3_T ? 2'h1 : _GEN_145; // @[playground/src/noop/memory.scala 322:37 323:25]
  reg [31:0] inst3_r; // @[playground/src/noop/memory.scala 330:30]
  reg [63:0] pc3_r; // @[playground/src/noop/memory.scala 331:30]
  reg [63:0] excep3_r_cause; // @[playground/src/noop/memory.scala 332:30]
  reg [63:0] excep3_r_tval; // @[playground/src/noop/memory.scala 332:30]
  reg  excep3_r_en; // @[playground/src/noop/memory.scala 332:30]
  reg [63:0] excep3_r_pc; // @[playground/src/noop/memory.scala 332:30]
  reg [1:0] excep3_r_etype; // @[playground/src/noop/memory.scala 332:30]
  reg [4:0] dst3_r; // @[playground/src/noop/memory.scala 333:30]
  reg [63:0] dst_d3_r; // @[playground/src/noop/memory.scala 334:30]
  reg  dst_en3_r; // @[playground/src/noop/memory.scala 335:30]
  reg [11:0] csr_id3_r; // @[playground/src/noop/memory.scala 336:30]
  reg [63:0] csr_d3_r; // @[playground/src/noop/memory.scala 337:30]
  reg  csr_en3_r; // @[playground/src/noop/memory.scala 338:30]
  reg [11:0] rcsr_id3_r; // @[playground/src/noop/memory.scala 339:30]
  reg [1:0] special3_r; // @[playground/src/noop/memory.scala 340:30]
  reg  is_mmio_r; // @[playground/src/noop/memory.scala 341:30]
  reg  recov3_r; // @[playground/src/noop/memory.scala 342:30]
  wire [63:0] _GEN_156 = hs2 ? dst_d2_r : dst_d3_r; // @[playground/src/noop/memory.scala 349:14 354:21 334:30]
  wire  _GEN_170 = io_mem2rb_ready ? 1'h0 : valid3_r; // @[playground/src/noop/memory.scala 380:27 381:22 343:30]
  wire  _GEN_171 = hs2 | _GEN_170; // @[playground/src/noop/memory.scala 375:19 376:22]
  wire  _GEN_173 = _stall3_in_T & _GEN_171; // @[playground/src/noop/memory.scala 374:26 384:18]
  assign io_ex2mem_drop = drop2_r | io_mem2rb_drop; // @[playground/src/noop/memory.scala 103:31]
  assign io_ex2mem_stall = stall2_r & _stall3_in_T | io_mem2rb_stall; // @[playground/src/noop/memory.scala 106:45]
  assign io_ex2mem_ready = _stall1_in_T & _GEN_26; // @[playground/src/noop/memory.scala 166:20 165:21]
  assign io_mem2rb_inst = inst3_r; // @[playground/src/noop/memory.scala 386:25]
  assign io_mem2rb_pc = pc3_r; // @[playground/src/noop/memory.scala 387:25]
  assign io_mem2rb_excep_cause = excep3_r_cause; // @[playground/src/noop/memory.scala 388:25]
  assign io_mem2rb_excep_tval = excep3_r_tval; // @[playground/src/noop/memory.scala 388:25]
  assign io_mem2rb_excep_en = excep3_r_en; // @[playground/src/noop/memory.scala 388:25]
  assign io_mem2rb_excep_pc = excep3_r_pc; // @[playground/src/noop/memory.scala 388:25]
  assign io_mem2rb_excep_etype = excep3_r_etype; // @[playground/src/noop/memory.scala 388:25]
  assign io_mem2rb_csr_id = csr_id3_r; // @[playground/src/noop/memory.scala 389:25]
  assign io_mem2rb_csr_d = csr_d3_r; // @[playground/src/noop/memory.scala 390:25]
  assign io_mem2rb_csr_en = csr_en3_r; // @[playground/src/noop/memory.scala 391:25]
  assign io_mem2rb_dst = dst3_r; // @[playground/src/noop/memory.scala 392:25]
  assign io_mem2rb_dst_d = dst_d3_r; // @[playground/src/noop/memory.scala 393:25]
  assign io_mem2rb_dst_en = dst_en3_r; // @[playground/src/noop/memory.scala 394:25]
  assign io_mem2rb_rcsr_id = rcsr_id3_r; // @[playground/src/noop/memory.scala 395:25]
  assign io_mem2rb_special = special3_r; // @[playground/src/noop/memory.scala 396:25]
  assign io_mem2rb_is_mmio = is_mmio_r; // @[playground/src/noop/memory.scala 397:25]
  assign io_mem2rb_recov = recov3_r; // @[playground/src/noop/memory.scala 398:25]
  assign io_mem2rb_valid = valid3_r; // @[playground/src/noop/memory.scala 399:25]
  assign io_dataRW_addr = hs1 ? io_va2pa_paddr : paddr2_r; // @[playground/src/noop/memory.scala 257:29]
  assign io_dataRW_wdata = hs1 ? mem_data1_r : mem_data2_r; // @[playground/src/noop/memory.scala 258:29]
  assign io_dataRW_dc_mode = hs1 ? _GEN_79 : _io_dataRW_dc_mode_T_2; // @[playground/src/noop/memory.scala 262:14 279:27]
  assign io_dataRW_amo = hs1 ? inst1_r[31:27] : inst2_r[31:27]; // @[playground/src/noop/memory.scala 259:29]
  assign io_va2pa_vaddr = hs_in ? io_ex2mem_mem_addr : mem_addr1_r; // @[playground/src/noop/memory.scala 161:27]
  assign io_va2pa_vvalid = _stall1_in_T ? _GEN_32 : _stall1_in_T & is_tlb_r & ~hs1; // @[playground/src/noop/memory.scala 172:20 162:21]
  assign io_va2pa_m_type = _GEN_9[3] ? 2'h3 : 2'h2; // @[playground/src/noop/memory.scala 164:27]
  assign io_d_mem1_id = dst1_r; // @[playground/src/noop/memory.scala 186:20]
  assign io_d_mem1_data = dst_d1_r; // @[playground/src/noop/memory.scala 187:20]
  assign io_d_mem1_state = ~dst_en1_r ? 2'h0 : _GEN_38; // @[playground/src/noop/memory.scala 188:21 189:25]
  assign io_d_mem2_id = dst2_r; // @[playground/src/noop/memory.scala 318:20]
  assign io_d_mem2_data = dst_d2_r; // @[playground/src/noop/memory.scala 319:20]
  assign io_d_mem2_state = ~dst_en2_r ? 2'h0 : _GEN_146; // @[playground/src/noop/memory.scala 320:21 321:25]
  assign io_d_mem3_id = dst3_r; // @[playground/src/noop/memory.scala 401:20]
  assign io_d_mem3_data = dst_d3_r; // @[playground/src/noop/memory.scala 402:20]
  assign io_d_mem3_state = valid3_r & dst_en3_r ? 2'h1 : 2'h0; // @[playground/src/noop/memory.scala 403:32 404:25 406:25]
  always @(posedge clock) begin
    if (reset) begin // @[playground/src/noop/memory.scala 95:26]
      drop2_r <= 1'h0; // @[playground/src/noop/memory.scala 95:26]
    end else begin
      drop2_r <= _GEN_141;
    end
    if (reset) begin // @[playground/src/noop/memory.scala 98:27]
      stall2_r <= 1'h0; // @[playground/src/noop/memory.scala 98:27]
    end else begin
      stall2_r <= _GEN_141;
    end
    if (reset) begin // @[playground/src/noop/memory.scala 111:30]
      inst1_r <= 32'h0; // @[playground/src/noop/memory.scala 111:30]
    end else if (hs_in) begin // @[playground/src/noop/memory.scala 142:16]
      inst1_r <= io_ex2mem_inst; // @[playground/src/noop/memory.scala 143:21]
    end
    if (reset) begin // @[playground/src/noop/memory.scala 112:30]
      pc1_r <= 64'h0; // @[playground/src/noop/memory.scala 112:30]
    end else if (hs_in) begin // @[playground/src/noop/memory.scala 142:16]
      pc1_r <= io_ex2mem_pc; // @[playground/src/noop/memory.scala 144:21]
    end
    if (reset) begin // @[playground/src/noop/memory.scala 113:30]
      excep1_r_cause <= 64'h0; // @[playground/src/noop/memory.scala 113:30]
    end else if (hs_in) begin // @[playground/src/noop/memory.scala 142:16]
      excep1_r_cause <= io_ex2mem_excep_cause; // @[playground/src/noop/memory.scala 145:21]
    end
    if (reset) begin // @[playground/src/noop/memory.scala 113:30]
      excep1_r_tval <= 64'h0; // @[playground/src/noop/memory.scala 113:30]
    end else if (hs_in) begin // @[playground/src/noop/memory.scala 142:16]
      excep1_r_tval <= io_ex2mem_excep_tval; // @[playground/src/noop/memory.scala 145:21]
    end
    if (reset) begin // @[playground/src/noop/memory.scala 113:30]
      excep1_r_en <= 1'h0; // @[playground/src/noop/memory.scala 113:30]
    end else if (hs_in) begin // @[playground/src/noop/memory.scala 142:16]
      excep1_r_en <= io_ex2mem_excep_en; // @[playground/src/noop/memory.scala 145:21]
    end
    if (reset) begin // @[playground/src/noop/memory.scala 113:30]
      excep1_r_pc <= 64'h0; // @[playground/src/noop/memory.scala 113:30]
    end else if (hs_in) begin // @[playground/src/noop/memory.scala 142:16]
      excep1_r_pc <= io_ex2mem_excep_pc; // @[playground/src/noop/memory.scala 145:21]
    end
    if (reset) begin // @[playground/src/noop/memory.scala 113:30]
      excep1_r_etype <= 2'h0; // @[playground/src/noop/memory.scala 113:30]
    end else if (hs_in) begin // @[playground/src/noop/memory.scala 142:16]
      excep1_r_etype <= io_ex2mem_excep_etype; // @[playground/src/noop/memory.scala 145:21]
    end
    if (reset) begin // @[playground/src/noop/memory.scala 114:30]
      ctrl1_r_dcMode <= 5'h0; // @[playground/src/noop/memory.scala 114:30]
    end else if (hs_in) begin // @[playground/src/noop/memory.scala 142:16]
      ctrl1_r_dcMode <= io_ex2mem_ctrl_dcMode; // @[playground/src/noop/memory.scala 146:21]
    end
    if (reset) begin // @[playground/src/noop/memory.scala 115:30]
      mem_addr1_r <= 64'h0; // @[playground/src/noop/memory.scala 115:30]
    end else if (hs_in) begin // @[playground/src/noop/memory.scala 142:16]
      mem_addr1_r <= io_ex2mem_mem_addr; // @[playground/src/noop/memory.scala 147:21]
    end
    if (reset) begin // @[playground/src/noop/memory.scala 116:30]
      mem_data1_r <= 64'h0; // @[playground/src/noop/memory.scala 116:30]
    end else if (hs_in) begin // @[playground/src/noop/memory.scala 142:16]
      mem_data1_r <= io_ex2mem_mem_data; // @[playground/src/noop/memory.scala 148:21]
    end
    if (reset) begin // @[playground/src/noop/memory.scala 117:30]
      dst1_r <= 5'h0; // @[playground/src/noop/memory.scala 117:30]
    end else if (hs_in) begin // @[playground/src/noop/memory.scala 142:16]
      dst1_r <= io_ex2mem_dst; // @[playground/src/noop/memory.scala 149:21]
    end
    if (reset) begin // @[playground/src/noop/memory.scala 118:30]
      dst_d1_r <= 64'h0; // @[playground/src/noop/memory.scala 118:30]
    end else if (hs_in) begin // @[playground/src/noop/memory.scala 142:16]
      dst_d1_r <= io_ex2mem_dst_d; // @[playground/src/noop/memory.scala 150:21]
    end
    if (reset) begin // @[playground/src/noop/memory.scala 119:30]
      dst_en1_r <= 1'h0; // @[playground/src/noop/memory.scala 119:30]
    end else if (hs_in) begin // @[playground/src/noop/memory.scala 142:16]
      dst_en1_r <= io_ex2mem_ctrl_writeRegEn; // @[playground/src/noop/memory.scala 151:21]
    end
    if (reset) begin // @[playground/src/noop/memory.scala 120:30]
      csr_id1_r <= 12'h0; // @[playground/src/noop/memory.scala 120:30]
    end else if (hs_in) begin // @[playground/src/noop/memory.scala 142:16]
      csr_id1_r <= io_ex2mem_csr_id; // @[playground/src/noop/memory.scala 152:21]
    end
    if (reset) begin // @[playground/src/noop/memory.scala 121:30]
      csr_d1_r <= 64'h0; // @[playground/src/noop/memory.scala 121:30]
    end else if (hs_in) begin // @[playground/src/noop/memory.scala 142:16]
      csr_d1_r <= io_ex2mem_csr_d; // @[playground/src/noop/memory.scala 153:21]
    end
    if (reset) begin // @[playground/src/noop/memory.scala 122:30]
      csr_en1_r <= 1'h0; // @[playground/src/noop/memory.scala 122:30]
    end else if (hs_in) begin // @[playground/src/noop/memory.scala 142:16]
      csr_en1_r <= io_ex2mem_ctrl_writeCSREn; // @[playground/src/noop/memory.scala 154:21]
    end
    if (reset) begin // @[playground/src/noop/memory.scala 123:30]
      rcsr_id1_r <= 12'h0; // @[playground/src/noop/memory.scala 123:30]
    end else if (hs_in) begin // @[playground/src/noop/memory.scala 142:16]
      rcsr_id1_r <= io_ex2mem_rcsr_id; // @[playground/src/noop/memory.scala 155:21]
    end
    if (reset) begin // @[playground/src/noop/memory.scala 124:30]
      special1_r <= 2'h0; // @[playground/src/noop/memory.scala 124:30]
    end else if (hs_in) begin // @[playground/src/noop/memory.scala 142:16]
      special1_r <= io_ex2mem_special; // @[playground/src/noop/memory.scala 157:21]
    end
    if (reset) begin // @[playground/src/noop/memory.scala 125:30]
      indi1_r <= 2'h0; // @[playground/src/noop/memory.scala 125:30]
    end else if (hs_in) begin // @[playground/src/noop/memory.scala 142:16]
      indi1_r <= io_ex2mem_indi; // @[playground/src/noop/memory.scala 156:21]
    end
    if (reset) begin // @[playground/src/noop/memory.scala 126:30]
      recov1_r <= 1'h0; // @[playground/src/noop/memory.scala 126:30]
    end else if (hs_in) begin // @[playground/src/noop/memory.scala 142:16]
      recov1_r <= io_ex2mem_recov; // @[playground/src/noop/memory.scala 158:21]
    end
    if (reset) begin // @[playground/src/noop/memory.scala 128:30]
      valid1_r <= 1'h0; // @[playground/src/noop/memory.scala 128:30]
    end else begin
      valid1_r <= _GEN_33;
    end
    if (reset) begin // @[playground/src/noop/memory.scala 134:30]
      is_tlb_r <= 1'h0; // @[playground/src/noop/memory.scala 134:30]
    end else begin
      is_tlb_r <= _GEN_34;
    end
    if (reset) begin // @[playground/src/noop/memory.scala 135:30]
      drop_tlb <= 1'h0; // @[playground/src/noop/memory.scala 135:30]
    end else if (inp_tlb_valid2 & drop_tlb) begin // @[playground/src/noop/memory.scala 224:65]
      drop_tlb <= 1'h0; // @[playground/src/noop/memory.scala 225:18]
    end else if (!(_stall1_in_T)) begin // @[playground/src/noop/memory.scala 172:20]
      drop_tlb <= is_tlb_r & ~io_va2pa_pvalid; // @[playground/src/noop/memory.scala 183:18]
    end
    if (reset) begin // @[playground/src/noop/memory.scala 214:30]
      valid2_r <= 1'h0; // @[playground/src/noop/memory.scala 214:30]
    end else begin
      valid2_r <= _GEN_127;
    end
    if (reset) begin // @[playground/src/noop/memory.scala 343:30]
      valid3_r <= 1'h0; // @[playground/src/noop/memory.scala 343:30]
    end else begin
      valid3_r <= _GEN_173;
    end
    if (reset) begin // @[playground/src/noop/memory.scala 201:30]
      ctrl2_r_dcMode <= 5'h0; // @[playground/src/noop/memory.scala 201:30]
    end else if (_stall3_in_T) begin // @[playground/src/noop/memory.scala 293:20]
      if (hs1) begin // @[playground/src/noop/memory.scala 294:18]
        if (io_va2pa_tlb_excep_en & _tlb_valid2_T_1) begin // @[playground/src/noop/memory.scala 296:53]
          ctrl2_r_dcMode <= 5'h0; // @[playground/src/noop/memory.scala 302:29]
        end else begin
          ctrl2_r_dcMode <= _GEN_84;
        end
      end else begin
        ctrl2_r_dcMode <= _GEN_84;
      end
    end else begin
      ctrl2_r_dcMode <= _GEN_84;
    end
    if (reset) begin // @[playground/src/noop/memory.scala 255:30]
      drop_dc <= 1'h0; // @[playground/src/noop/memory.scala 255:30]
    end else if (io_dataRW_rvalid) begin // @[playground/src/noop/memory.scala 364:27]
      drop_dc <= 1'h0; // @[playground/src/noop/memory.scala 365:17]
    end else if (!(_stall3_in_T)) begin // @[playground/src/noop/memory.scala 293:20]
      drop_dc <= is_dc_r & ~io_dataRW_rvalid; // @[playground/src/noop/memory.scala 315:18]
    end
    if (reset) begin // @[playground/src/noop/memory.scala 198:30]
      inst2_r <= 32'h0; // @[playground/src/noop/memory.scala 198:30]
    end else if (hs1) begin // @[playground/src/noop/memory.scala 228:14]
      inst2_r <= inst1_r; // @[playground/src/noop/memory.scala 229:21]
    end
    if (reset) begin // @[playground/src/noop/memory.scala 199:30]
      pc2_r <= 64'h0; // @[playground/src/noop/memory.scala 199:30]
    end else if (hs1) begin // @[playground/src/noop/memory.scala 228:14]
      pc2_r <= pc1_r; // @[playground/src/noop/memory.scala 230:21]
    end
    if (reset) begin // @[playground/src/noop/memory.scala 200:30]
      excep2_r_cause <= 64'h0; // @[playground/src/noop/memory.scala 200:30]
    end else if (_stall3_in_T) begin // @[playground/src/noop/memory.scala 293:20]
      if (hs1) begin // @[playground/src/noop/memory.scala 294:18]
        if (io_va2pa_tlb_excep_en & _tlb_valid2_T_1) begin // @[playground/src/noop/memory.scala 296:53]
          excep2_r_cause <= io_va2pa_tlb_excep_cause; // @[playground/src/noop/memory.scala 297:33]
        end else begin
          excep2_r_cause <= _GEN_46;
        end
      end else begin
        excep2_r_cause <= _GEN_46;
      end
    end else begin
      excep2_r_cause <= _GEN_46;
    end
    if (reset) begin // @[playground/src/noop/memory.scala 200:30]
      excep2_r_tval <= 64'h0; // @[playground/src/noop/memory.scala 200:30]
    end else if (_stall3_in_T) begin // @[playground/src/noop/memory.scala 293:20]
      if (hs1) begin // @[playground/src/noop/memory.scala 294:18]
        if (io_va2pa_tlb_excep_en & _tlb_valid2_T_1) begin // @[playground/src/noop/memory.scala 296:53]
          excep2_r_tval <= io_va2pa_tlb_excep_tval; // @[playground/src/noop/memory.scala 298:33]
        end else begin
          excep2_r_tval <= _GEN_47;
        end
      end else begin
        excep2_r_tval <= _GEN_47;
      end
    end else begin
      excep2_r_tval <= _GEN_47;
    end
    if (reset) begin // @[playground/src/noop/memory.scala 200:30]
      excep2_r_en <= 1'h0; // @[playground/src/noop/memory.scala 200:30]
    end else if (_stall3_in_T) begin // @[playground/src/noop/memory.scala 293:20]
      if (hs1) begin // @[playground/src/noop/memory.scala 294:18]
        excep2_r_en <= _GEN_94;
      end else begin
        excep2_r_en <= _GEN_48;
      end
    end else begin
      excep2_r_en <= _GEN_48;
    end
    if (reset) begin // @[playground/src/noop/memory.scala 200:30]
      excep2_r_pc <= 64'h0; // @[playground/src/noop/memory.scala 200:30]
    end else if (_stall3_in_T) begin // @[playground/src/noop/memory.scala 293:20]
      if (hs1) begin // @[playground/src/noop/memory.scala 294:18]
        if (io_va2pa_tlb_excep_en & _tlb_valid2_T_1) begin // @[playground/src/noop/memory.scala 296:53]
          excep2_r_pc <= pc1_r; // @[playground/src/noop/memory.scala 300:33]
        end else begin
          excep2_r_pc <= _GEN_49;
        end
      end else begin
        excep2_r_pc <= _GEN_49;
      end
    end else begin
      excep2_r_pc <= _GEN_49;
    end
    if (reset) begin // @[playground/src/noop/memory.scala 200:30]
      excep2_r_etype <= 2'h0; // @[playground/src/noop/memory.scala 200:30]
    end else if (_stall3_in_T) begin // @[playground/src/noop/memory.scala 293:20]
      if (hs1) begin // @[playground/src/noop/memory.scala 294:18]
        if (io_va2pa_tlb_excep_en & _tlb_valid2_T_1) begin // @[playground/src/noop/memory.scala 296:53]
          excep2_r_etype <= 2'h0; // @[playground/src/noop/memory.scala 301:33]
        end else begin
          excep2_r_etype <= _GEN_50;
        end
      end else begin
        excep2_r_etype <= _GEN_50;
      end
    end else begin
      excep2_r_etype <= _GEN_50;
    end
    if (reset) begin // @[playground/src/noop/memory.scala 202:30]
      mem_data2_r <= 64'h0; // @[playground/src/noop/memory.scala 202:30]
    end else if (hs1) begin // @[playground/src/noop/memory.scala 228:14]
      mem_data2_r <= mem_data1_r; // @[playground/src/noop/memory.scala 232:21]
    end
    if (reset) begin // @[playground/src/noop/memory.scala 203:30]
      dst2_r <= 5'h0; // @[playground/src/noop/memory.scala 203:30]
    end else if (hs1) begin // @[playground/src/noop/memory.scala 228:14]
      dst2_r <= dst1_r; // @[playground/src/noop/memory.scala 234:21]
    end
    if (reset) begin // @[playground/src/noop/memory.scala 204:30]
      dst_d2_r <= 64'h0; // @[playground/src/noop/memory.scala 204:30]
    end else if (hs1) begin // @[playground/src/noop/memory.scala 262:14]
      if (stage2_is_excep) begin // @[playground/src/noop/memory.scala 263:30]
        dst_d2_r <= _GEN_59;
      end else if (indi1_r[1] & sc_valid) begin // @[playground/src/noop/memory.scala 266:53]
        dst_d2_r <= 64'h0; // @[playground/src/noop/memory.scala 269:25]
      end else begin
        dst_d2_r <= _GEN_74;
      end
    end else begin
      dst_d2_r <= _GEN_59;
    end
    if (reset) begin // @[playground/src/noop/memory.scala 205:30]
      dst_en2_r <= 1'h0; // @[playground/src/noop/memory.scala 205:30]
    end else if (_stall3_in_T) begin // @[playground/src/noop/memory.scala 293:20]
      if (hs1) begin // @[playground/src/noop/memory.scala 294:18]
        if (io_va2pa_tlb_excep_en & _tlb_valid2_T_1) begin // @[playground/src/noop/memory.scala 296:53]
          dst_en2_r <= 1'h0; // @[playground/src/noop/memory.scala 303:29]
        end else begin
          dst_en2_r <= _GEN_85;
        end
      end else begin
        dst_en2_r <= _GEN_85;
      end
    end else begin
      dst_en2_r <= _GEN_85;
    end
    if (reset) begin // @[playground/src/noop/memory.scala 206:30]
      csr_id2_r <= 12'h0; // @[playground/src/noop/memory.scala 206:30]
    end else if (hs1) begin // @[playground/src/noop/memory.scala 228:14]
      csr_id2_r <= csr_id1_r; // @[playground/src/noop/memory.scala 237:21]
    end
    if (reset) begin // @[playground/src/noop/memory.scala 207:30]
      csr_d2_r <= 64'h0; // @[playground/src/noop/memory.scala 207:30]
    end else if (hs1) begin // @[playground/src/noop/memory.scala 228:14]
      csr_d2_r <= csr_d1_r; // @[playground/src/noop/memory.scala 238:21]
    end
    if (reset) begin // @[playground/src/noop/memory.scala 208:30]
      csr_en2_r <= 1'h0; // @[playground/src/noop/memory.scala 208:30]
    end else if (_stall3_in_T) begin // @[playground/src/noop/memory.scala 293:20]
      if (hs1) begin // @[playground/src/noop/memory.scala 294:18]
        if (io_va2pa_tlb_excep_en & _tlb_valid2_T_1) begin // @[playground/src/noop/memory.scala 296:53]
          csr_en2_r <= 1'h0; // @[playground/src/noop/memory.scala 304:29]
        end else begin
          csr_en2_r <= _GEN_63;
        end
      end else begin
        csr_en2_r <= _GEN_63;
      end
    end else begin
      csr_en2_r <= _GEN_63;
    end
    if (reset) begin // @[playground/src/noop/memory.scala 209:30]
      rcsr_id2_r <= 12'h0; // @[playground/src/noop/memory.scala 209:30]
    end else if (hs1) begin // @[playground/src/noop/memory.scala 228:14]
      rcsr_id2_r <= rcsr_id1_r; // @[playground/src/noop/memory.scala 240:21]
    end
    if (reset) begin // @[playground/src/noop/memory.scala 210:30]
      special2_r <= 2'h0; // @[playground/src/noop/memory.scala 210:30]
    end else if (hs1) begin // @[playground/src/noop/memory.scala 228:14]
      special2_r <= special1_r; // @[playground/src/noop/memory.scala 241:21]
    end
    if (reset) begin // @[playground/src/noop/memory.scala 211:30]
      paddr2_r <= 32'h0; // @[playground/src/noop/memory.scala 211:30]
    end else if (hs1) begin // @[playground/src/noop/memory.scala 228:14]
      paddr2_r <= io_va2pa_paddr; // @[playground/src/noop/memory.scala 244:21]
    end
    if (reset) begin // @[playground/src/noop/memory.scala 213:30]
      recov2_r <= 1'h0; // @[playground/src/noop/memory.scala 213:30]
    end else if (_stall3_in_T) begin // @[playground/src/noop/memory.scala 293:20]
      if (hs1) begin // @[playground/src/noop/memory.scala 294:18]
        recov2_r <= _GEN_106;
      end else begin
        recov2_r <= _GEN_67;
      end
    end else begin
      recov2_r <= _GEN_67;
    end
    if (reset) begin // @[playground/src/noop/memory.scala 215:30]
      dc_hs_r <= 1'h0; // @[playground/src/noop/memory.scala 215:30]
    end else if (_stall3_in_T) begin // @[playground/src/noop/memory.scala 293:20]
      if (hs1) begin // @[playground/src/noop/memory.scala 294:18]
        if (io_va2pa_tlb_excep_en & _tlb_valid2_T_1) begin // @[playground/src/noop/memory.scala 296:53]
          dc_hs_r <= _GEN_87;
        end else begin
          dc_hs_r <= _GEN_91;
        end
      end else if (hs2) begin // @[playground/src/noop/memory.scala 309:24]
        dc_hs_r <= 1'h0; // @[playground/src/noop/memory.scala 311:22]
      end else begin
        dc_hs_r <= _GEN_87;
      end
    end else begin
      dc_hs_r <= _GEN_87;
    end
    if (reset) begin // @[playground/src/noop/memory.scala 217:30]
      lr_addr_r <= 32'h0; // @[playground/src/noop/memory.scala 217:30]
    end else if (hs1) begin // @[playground/src/noop/memory.scala 228:14]
      if (indi1_r[0] & ~stage2_is_excep) begin // @[playground/src/noop/memory.scala 245:55]
        lr_addr_r <= io_va2pa_paddr; // @[playground/src/noop/memory.scala 247:25]
      end
    end
    if (reset) begin // @[playground/src/noop/memory.scala 218:30]
      lr_valid_r <= 1'h0; // @[playground/src/noop/memory.scala 218:30]
    end else if (hs1) begin // @[playground/src/noop/memory.scala 228:14]
      if (excep1_r_en & excep1_r_cause[63]) begin // @[playground/src/noop/memory.scala 249:48]
        lr_valid_r <= 1'h0; // @[playground/src/noop/memory.scala 250:25]
      end else begin
        lr_valid_r <= _GEN_41;
      end
    end
    if (reset) begin // @[playground/src/noop/memory.scala 330:30]
      inst3_r <= 32'h0; // @[playground/src/noop/memory.scala 330:30]
    end else if (hs2) begin // @[playground/src/noop/memory.scala 349:14]
      inst3_r <= inst2_r; // @[playground/src/noop/memory.scala 350:21]
    end
    if (reset) begin // @[playground/src/noop/memory.scala 331:30]
      pc3_r <= 64'h0; // @[playground/src/noop/memory.scala 331:30]
    end else if (hs2) begin // @[playground/src/noop/memory.scala 349:14]
      pc3_r <= pc2_r; // @[playground/src/noop/memory.scala 351:21]
    end
    if (reset) begin // @[playground/src/noop/memory.scala 332:30]
      excep3_r_cause <= 64'h0; // @[playground/src/noop/memory.scala 332:30]
    end else if (hs2) begin // @[playground/src/noop/memory.scala 349:14]
      excep3_r_cause <= excep2_r_cause; // @[playground/src/noop/memory.scala 352:21]
    end
    if (reset) begin // @[playground/src/noop/memory.scala 332:30]
      excep3_r_tval <= 64'h0; // @[playground/src/noop/memory.scala 332:30]
    end else if (hs2) begin // @[playground/src/noop/memory.scala 349:14]
      excep3_r_tval <= excep2_r_tval; // @[playground/src/noop/memory.scala 352:21]
    end
    if (reset) begin // @[playground/src/noop/memory.scala 332:30]
      excep3_r_en <= 1'h0; // @[playground/src/noop/memory.scala 332:30]
    end else if (hs2) begin // @[playground/src/noop/memory.scala 349:14]
      excep3_r_en <= excep2_r_en; // @[playground/src/noop/memory.scala 352:21]
    end
    if (reset) begin // @[playground/src/noop/memory.scala 332:30]
      excep3_r_pc <= 64'h0; // @[playground/src/noop/memory.scala 332:30]
    end else if (hs2) begin // @[playground/src/noop/memory.scala 349:14]
      excep3_r_pc <= excep2_r_pc; // @[playground/src/noop/memory.scala 352:21]
    end
    if (reset) begin // @[playground/src/noop/memory.scala 332:30]
      excep3_r_etype <= 2'h0; // @[playground/src/noop/memory.scala 332:30]
    end else if (hs2) begin // @[playground/src/noop/memory.scala 349:14]
      excep3_r_etype <= excep2_r_etype; // @[playground/src/noop/memory.scala 352:21]
    end
    if (reset) begin // @[playground/src/noop/memory.scala 333:30]
      dst3_r <= 5'h0; // @[playground/src/noop/memory.scala 333:30]
    end else if (hs2) begin // @[playground/src/noop/memory.scala 349:14]
      dst3_r <= dst2_r; // @[playground/src/noop/memory.scala 353:21]
    end
    if (reset) begin // @[playground/src/noop/memory.scala 334:30]
      dst_d3_r <= 64'h0; // @[playground/src/noop/memory.scala 334:30]
    end else if (_stall3_in_T) begin // @[playground/src/noop/memory.scala 374:26]
      if (hs2) begin // @[playground/src/noop/memory.scala 375:19]
        if (is_dc_r) begin // @[playground/src/noop/memory.scala 377:26]
          dst_d3_r <= io_dataRW_rdata; // @[playground/src/noop/memory.scala 378:26]
        end else begin
          dst_d3_r <= _GEN_156;
        end
      end else begin
        dst_d3_r <= _GEN_156;
      end
    end else begin
      dst_d3_r <= _GEN_156;
    end
    if (reset) begin // @[playground/src/noop/memory.scala 335:30]
      dst_en3_r <= 1'h0; // @[playground/src/noop/memory.scala 335:30]
    end else if (hs2) begin // @[playground/src/noop/memory.scala 349:14]
      dst_en3_r <= dst_en2_r; // @[playground/src/noop/memory.scala 355:21]
    end
    if (reset) begin // @[playground/src/noop/memory.scala 336:30]
      csr_id3_r <= 12'h0; // @[playground/src/noop/memory.scala 336:30]
    end else if (hs2) begin // @[playground/src/noop/memory.scala 349:14]
      csr_id3_r <= csr_id2_r; // @[playground/src/noop/memory.scala 356:21]
    end
    if (reset) begin // @[playground/src/noop/memory.scala 337:30]
      csr_d3_r <= 64'h0; // @[playground/src/noop/memory.scala 337:30]
    end else if (hs2) begin // @[playground/src/noop/memory.scala 349:14]
      csr_d3_r <= csr_d2_r; // @[playground/src/noop/memory.scala 357:21]
    end
    if (reset) begin // @[playground/src/noop/memory.scala 338:30]
      csr_en3_r <= 1'h0; // @[playground/src/noop/memory.scala 338:30]
    end else if (hs2) begin // @[playground/src/noop/memory.scala 349:14]
      csr_en3_r <= csr_en2_r; // @[playground/src/noop/memory.scala 358:21]
    end
    if (reset) begin // @[playground/src/noop/memory.scala 339:30]
      rcsr_id3_r <= 12'h0; // @[playground/src/noop/memory.scala 339:30]
    end else if (hs2) begin // @[playground/src/noop/memory.scala 349:14]
      rcsr_id3_r <= rcsr_id2_r; // @[playground/src/noop/memory.scala 359:21]
    end
    if (reset) begin // @[playground/src/noop/memory.scala 340:30]
      special3_r <= 2'h0; // @[playground/src/noop/memory.scala 340:30]
    end else if (hs2) begin // @[playground/src/noop/memory.scala 349:14]
      special3_r <= special2_r; // @[playground/src/noop/memory.scala 360:21]
    end
    if (reset) begin // @[playground/src/noop/memory.scala 341:30]
      is_mmio_r <= 1'h0; // @[playground/src/noop/memory.scala 341:30]
    end else if (hs2) begin // @[playground/src/noop/memory.scala 349:14]
      is_mmio_r <= is_dc_r & paddr2_r < 32'h80000000; // @[playground/src/noop/memory.scala 362:21]
    end
    if (reset) begin // @[playground/src/noop/memory.scala 342:30]
      recov3_r <= 1'h0; // @[playground/src/noop/memory.scala 342:30]
    end else if (hs2) begin // @[playground/src/noop/memory.scala 349:14]
      recov3_r <= recov2_r; // @[playground/src/noop/memory.scala 361:21]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  drop2_r = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  stall2_r = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  inst1_r = _RAND_2[31:0];
  _RAND_3 = {2{`RANDOM}};
  pc1_r = _RAND_3[63:0];
  _RAND_4 = {2{`RANDOM}};
  excep1_r_cause = _RAND_4[63:0];
  _RAND_5 = {2{`RANDOM}};
  excep1_r_tval = _RAND_5[63:0];
  _RAND_6 = {1{`RANDOM}};
  excep1_r_en = _RAND_6[0:0];
  _RAND_7 = {2{`RANDOM}};
  excep1_r_pc = _RAND_7[63:0];
  _RAND_8 = {1{`RANDOM}};
  excep1_r_etype = _RAND_8[1:0];
  _RAND_9 = {1{`RANDOM}};
  ctrl1_r_dcMode = _RAND_9[4:0];
  _RAND_10 = {2{`RANDOM}};
  mem_addr1_r = _RAND_10[63:0];
  _RAND_11 = {2{`RANDOM}};
  mem_data1_r = _RAND_11[63:0];
  _RAND_12 = {1{`RANDOM}};
  dst1_r = _RAND_12[4:0];
  _RAND_13 = {2{`RANDOM}};
  dst_d1_r = _RAND_13[63:0];
  _RAND_14 = {1{`RANDOM}};
  dst_en1_r = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  csr_id1_r = _RAND_15[11:0];
  _RAND_16 = {2{`RANDOM}};
  csr_d1_r = _RAND_16[63:0];
  _RAND_17 = {1{`RANDOM}};
  csr_en1_r = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  rcsr_id1_r = _RAND_18[11:0];
  _RAND_19 = {1{`RANDOM}};
  special1_r = _RAND_19[1:0];
  _RAND_20 = {1{`RANDOM}};
  indi1_r = _RAND_20[1:0];
  _RAND_21 = {1{`RANDOM}};
  recov1_r = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  valid1_r = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  is_tlb_r = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  drop_tlb = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  valid2_r = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  valid3_r = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  ctrl2_r_dcMode = _RAND_27[4:0];
  _RAND_28 = {1{`RANDOM}};
  drop_dc = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  inst2_r = _RAND_29[31:0];
  _RAND_30 = {2{`RANDOM}};
  pc2_r = _RAND_30[63:0];
  _RAND_31 = {2{`RANDOM}};
  excep2_r_cause = _RAND_31[63:0];
  _RAND_32 = {2{`RANDOM}};
  excep2_r_tval = _RAND_32[63:0];
  _RAND_33 = {1{`RANDOM}};
  excep2_r_en = _RAND_33[0:0];
  _RAND_34 = {2{`RANDOM}};
  excep2_r_pc = _RAND_34[63:0];
  _RAND_35 = {1{`RANDOM}};
  excep2_r_etype = _RAND_35[1:0];
  _RAND_36 = {2{`RANDOM}};
  mem_data2_r = _RAND_36[63:0];
  _RAND_37 = {1{`RANDOM}};
  dst2_r = _RAND_37[4:0];
  _RAND_38 = {2{`RANDOM}};
  dst_d2_r = _RAND_38[63:0];
  _RAND_39 = {1{`RANDOM}};
  dst_en2_r = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  csr_id2_r = _RAND_40[11:0];
  _RAND_41 = {2{`RANDOM}};
  csr_d2_r = _RAND_41[63:0];
  _RAND_42 = {1{`RANDOM}};
  csr_en2_r = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  rcsr_id2_r = _RAND_43[11:0];
  _RAND_44 = {1{`RANDOM}};
  special2_r = _RAND_44[1:0];
  _RAND_45 = {1{`RANDOM}};
  paddr2_r = _RAND_45[31:0];
  _RAND_46 = {1{`RANDOM}};
  recov2_r = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  dc_hs_r = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  lr_addr_r = _RAND_48[31:0];
  _RAND_49 = {1{`RANDOM}};
  lr_valid_r = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  inst3_r = _RAND_50[31:0];
  _RAND_51 = {2{`RANDOM}};
  pc3_r = _RAND_51[63:0];
  _RAND_52 = {2{`RANDOM}};
  excep3_r_cause = _RAND_52[63:0];
  _RAND_53 = {2{`RANDOM}};
  excep3_r_tval = _RAND_53[63:0];
  _RAND_54 = {1{`RANDOM}};
  excep3_r_en = _RAND_54[0:0];
  _RAND_55 = {2{`RANDOM}};
  excep3_r_pc = _RAND_55[63:0];
  _RAND_56 = {1{`RANDOM}};
  excep3_r_etype = _RAND_56[1:0];
  _RAND_57 = {1{`RANDOM}};
  dst3_r = _RAND_57[4:0];
  _RAND_58 = {2{`RANDOM}};
  dst_d3_r = _RAND_58[63:0];
  _RAND_59 = {1{`RANDOM}};
  dst_en3_r = _RAND_59[0:0];
  _RAND_60 = {1{`RANDOM}};
  csr_id3_r = _RAND_60[11:0];
  _RAND_61 = {2{`RANDOM}};
  csr_d3_r = _RAND_61[63:0];
  _RAND_62 = {1{`RANDOM}};
  csr_en3_r = _RAND_62[0:0];
  _RAND_63 = {1{`RANDOM}};
  rcsr_id3_r = _RAND_63[11:0];
  _RAND_64 = {1{`RANDOM}};
  special3_r = _RAND_64[1:0];
  _RAND_65 = {1{`RANDOM}};
  is_mmio_r = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  recov3_r = _RAND_66[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Writeback(
  input         clock,
  input         reset,
  input  [31:0] io_mem2rb_inst, // @[playground/src/noop/writeback.scala 10:16]
  input  [63:0] io_mem2rb_pc, // @[playground/src/noop/writeback.scala 10:16]
  input  [63:0] io_mem2rb_excep_cause, // @[playground/src/noop/writeback.scala 10:16]
  input  [63:0] io_mem2rb_excep_tval, // @[playground/src/noop/writeback.scala 10:16]
  input         io_mem2rb_excep_en, // @[playground/src/noop/writeback.scala 10:16]
  input  [63:0] io_mem2rb_excep_pc, // @[playground/src/noop/writeback.scala 10:16]
  input  [1:0]  io_mem2rb_excep_etype, // @[playground/src/noop/writeback.scala 10:16]
  input  [11:0] io_mem2rb_csr_id, // @[playground/src/noop/writeback.scala 10:16]
  input  [63:0] io_mem2rb_csr_d, // @[playground/src/noop/writeback.scala 10:16]
  input         io_mem2rb_csr_en, // @[playground/src/noop/writeback.scala 10:16]
  input  [4:0]  io_mem2rb_dst, // @[playground/src/noop/writeback.scala 10:16]
  input  [63:0] io_mem2rb_dst_d, // @[playground/src/noop/writeback.scala 10:16]
  input         io_mem2rb_dst_en, // @[playground/src/noop/writeback.scala 10:16]
  input  [11:0] io_mem2rb_rcsr_id, // @[playground/src/noop/writeback.scala 10:16]
  input  [1:0]  io_mem2rb_special, // @[playground/src/noop/writeback.scala 10:16]
  input         io_mem2rb_is_mmio, // @[playground/src/noop/writeback.scala 10:16]
  output        io_mem2rb_drop, // @[playground/src/noop/writeback.scala 10:16]
  output        io_mem2rb_stall, // @[playground/src/noop/writeback.scala 10:16]
  input         io_mem2rb_recov, // @[playground/src/noop/writeback.scala 10:16]
  input         io_mem2rb_valid, // @[playground/src/noop/writeback.scala 10:16]
  output        io_mem2rb_ready, // @[playground/src/noop/writeback.scala 10:16]
  output [4:0]  io_wReg_id, // @[playground/src/noop/writeback.scala 10:16]
  output [63:0] io_wReg_data, // @[playground/src/noop/writeback.scala 10:16]
  output        io_wReg_en, // @[playground/src/noop/writeback.scala 10:16]
  output [11:0] io_wCsr_id, // @[playground/src/noop/writeback.scala 10:16]
  output [63:0] io_wCsr_data, // @[playground/src/noop/writeback.scala 10:16]
  output        io_wCsr_en, // @[playground/src/noop/writeback.scala 10:16]
  output [63:0] io_excep_cause, // @[playground/src/noop/writeback.scala 10:16]
  output [63:0] io_excep_tval, // @[playground/src/noop/writeback.scala 10:16]
  output        io_excep_en, // @[playground/src/noop/writeback.scala 10:16]
  output [63:0] io_excep_pc, // @[playground/src/noop/writeback.scala 10:16]
  output [1:0]  io_excep_etype, // @[playground/src/noop/writeback.scala 10:16]
  output [63:0] io_wb2if_seq_pc, // @[playground/src/noop/writeback.scala 10:16]
  output        io_wb2if_valid, // @[playground/src/noop/writeback.scala 10:16]
  output        io_recov, // @[playground/src/noop/writeback.scala 10:16]
  output        io_flush_tlb, // @[playground/src/noop/writeback.scala 10:16]
  output        io_flush_cache // @[playground/src/noop/writeback.scala 10:16]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [63:0] _RAND_12;
  reg [31:0] _RAND_13;
`endif // RANDOMIZE_REG_INIT
  wire  instFinish_clock; // @[playground/src/noop/writeback.scala 79:28]
  wire  instFinish_is_mmio; // @[playground/src/noop/writeback.scala 79:28]
  wire  instFinish_valid; // @[playground/src/noop/writeback.scala 79:28]
  wire [63:0] instFinish_pc; // @[playground/src/noop/writeback.scala 79:28]
  wire [31:0] instFinish_inst; // @[playground/src/noop/writeback.scala 79:28]
  wire [11:0] instFinish_rcsr_id; // @[playground/src/noop/writeback.scala 79:28]
  wire  transExcep_clock; // @[playground/src/noop/writeback.scala 87:28]
  wire  transExcep_intr; // @[playground/src/noop/writeback.scala 87:28]
  wire [63:0] transExcep_cause; // @[playground/src/noop/writeback.scala 87:28]
  wire [63:0] transExcep_pc; // @[playground/src/noop/writeback.scala 87:28]
  reg  recov_r; // @[playground/src/noop/writeback.scala 22:30]
  reg [63:0] forceJmp_seq_pc; // @[playground/src/noop/writeback.scala 25:30]
  reg  forceJmp_valid; // @[playground/src/noop/writeback.scala 25:30]
  reg  tlb_r; // @[playground/src/noop/writeback.scala 26:30]
  reg  cache_r; // @[playground/src/noop/writeback.scala 27:30]
  reg  valid_r; // @[playground/src/noop/writeback.scala 28:30]
  reg [63:0] excep_r_cause; // @[playground/src/noop/writeback.scala 29:30]
  reg  excep_r_en; // @[playground/src/noop/writeback.scala 29:30]
  reg [63:0] excep_r_pc; // @[playground/src/noop/writeback.scala 29:30]
  reg [1:0] excep_r_etype; // @[playground/src/noop/writeback.scala 29:30]
  reg [11:0] rcsr_id_r; // @[playground/src/noop/writeback.scala 30:30]
  reg [31:0] inst_r; // @[playground/src/noop/writeback.scala 40:30]
  reg [63:0] pc_r; // @[playground/src/noop/writeback.scala 41:30]
  wire  _T_4 = io_mem2rb_special != 2'h0 | io_mem2rb_recov & ~io_mem2rb_excep_en; // @[playground/src/noop/writeback.scala 67:44]
  wire [63:0] _forceJmp_seq_pc_T_1 = io_mem2rb_pc + 64'h4; // @[playground/src/noop/writeback.scala 69:49]
  wire  _T_5 = io_mem2rb_special == 2'h1; // @[playground/src/noop/writeback.scala 70:40]
  wire  _T_6 = io_mem2rb_special == 2'h2; // @[playground/src/noop/writeback.scala 72:46]
  wire  _GEN_2 = io_mem2rb_special == 2'h1 ? 1'h0 : _T_6; // @[playground/src/noop/writeback.scala 32:21 70:60]
  wire  _GEN_5 = (io_mem2rb_special != 2'h0 | io_mem2rb_recov & ~io_mem2rb_excep_en) & _T_5; // @[playground/src/noop/writeback.scala 33:21 67:88]
  wire  _GEN_6 = (io_mem2rb_special != 2'h0 | io_mem2rb_recov & ~io_mem2rb_excep_en) & _GEN_2; // @[playground/src/noop/writeback.scala 32:21 67:88]
  wire  _GEN_10 = io_mem2rb_valid & io_mem2rb_excep_en; // @[playground/src/noop/writeback.scala 49:21 56:30 60:29]
  wire  _GEN_13 = io_mem2rb_valid & io_mem2rb_recov; // @[playground/src/noop/writeback.scala 56:30 64:21 24:32]
  wire  _GEN_19 = io_mem2rb_valid & _T_4; // @[playground/src/noop/writeback.scala 34:21 56:30]
  wire  _GEN_21 = io_mem2rb_valid & _GEN_5; // @[playground/src/noop/writeback.scala 33:21 56:30]
  wire  _GEN_22 = io_mem2rb_valid & _GEN_6; // @[playground/src/noop/writeback.scala 32:21 56:30]
  reg  is_mmio_r; // @[playground/src/noop/writeback.scala 78:30]
  InstFinish instFinish ( // @[playground/src/noop/writeback.scala 79:28]
    .clock(instFinish_clock),
    .is_mmio(instFinish_is_mmio),
    .valid(instFinish_valid),
    .pc(instFinish_pc),
    .inst(instFinish_inst),
    .rcsr_id(instFinish_rcsr_id)
  );
  TransExcep transExcep ( // @[playground/src/noop/writeback.scala 87:28]
    .clock(transExcep_clock),
    .intr(transExcep_intr),
    .cause(transExcep_cause),
    .pc(transExcep_pc)
  );
  assign io_mem2rb_drop = 1'h0; // @[playground/src/noop/writeback.scala 38:21]
  assign io_mem2rb_stall = 1'h0; // @[playground/src/noop/writeback.scala 54:21]
  assign io_mem2rb_ready = io_mem2rb_valid; // @[playground/src/noop/writeback.scala 55:18 53:21]
  assign io_wReg_id = io_mem2rb_dst; // @[playground/src/noop/writeback.scala 42:21]
  assign io_wReg_data = io_mem2rb_dst_d; // @[playground/src/noop/writeback.scala 43:21]
  assign io_wReg_en = io_mem2rb_valid & io_mem2rb_dst_en; // @[playground/src/noop/writeback.scala 44:21 56:30 58:29]
  assign io_wCsr_id = io_mem2rb_csr_id; // @[playground/src/noop/writeback.scala 45:21]
  assign io_wCsr_data = io_mem2rb_csr_d; // @[playground/src/noop/writeback.scala 46:21]
  assign io_wCsr_en = io_mem2rb_valid & io_mem2rb_csr_en; // @[playground/src/noop/writeback.scala 47:21 56:30 59:29]
  assign io_excep_cause = io_mem2rb_excep_cause; // @[playground/src/noop/writeback.scala 48:21]
  assign io_excep_tval = io_mem2rb_excep_tval; // @[playground/src/noop/writeback.scala 48:21]
  assign io_excep_en = io_mem2rb_valid & io_mem2rb_excep_en; // @[playground/src/noop/writeback.scala 49:21 56:30 60:29]
  assign io_excep_pc = io_mem2rb_excep_pc; // @[playground/src/noop/writeback.scala 48:21]
  assign io_excep_etype = io_mem2rb_excep_etype; // @[playground/src/noop/writeback.scala 48:21]
  assign io_wb2if_seq_pc = forceJmp_seq_pc; // @[playground/src/noop/writeback.scala 52:21]
  assign io_wb2if_valid = forceJmp_valid; // @[playground/src/noop/writeback.scala 52:21]
  assign io_recov = recov_r; // @[playground/src/noop/writeback.scala 39:21]
  assign io_flush_tlb = tlb_r; // @[playground/src/noop/writeback.scala 50:21]
  assign io_flush_cache = cache_r; // @[playground/src/noop/writeback.scala 51:21]
  assign instFinish_clock = clock; // @[playground/src/noop/writeback.scala 80:29]
  assign instFinish_is_mmio = is_mmio_r; // @[playground/src/noop/writeback.scala 81:29]
  assign instFinish_valid = valid_r; // @[playground/src/noop/writeback.scala 82:29]
  assign instFinish_pc = pc_r; // @[playground/src/noop/writeback.scala 83:29]
  assign instFinish_inst = inst_r; // @[playground/src/noop/writeback.scala 84:29]
  assign instFinish_rcsr_id = rcsr_id_r; // @[playground/src/noop/writeback.scala 85:29]
  assign transExcep_clock = clock; // @[playground/src/noop/writeback.scala 88:29]
  assign transExcep_intr = excep_r_en & excep_r_etype == 2'h0; // @[playground/src/noop/writeback.scala 89:43]
  assign transExcep_cause = excep_r_cause; // @[playground/src/noop/writeback.scala 90:29]
  assign transExcep_pc = excep_r_pc; // @[playground/src/noop/writeback.scala 91:29]
  always @(posedge clock) begin
    if (reset) begin // @[playground/src/noop/writeback.scala 22:30]
      recov_r <= 1'h0; // @[playground/src/noop/writeback.scala 22:30]
    end else begin
      recov_r <= _GEN_13;
    end
    if (reset) begin // @[playground/src/noop/writeback.scala 25:30]
      forceJmp_seq_pc <= 64'h0; // @[playground/src/noop/writeback.scala 25:30]
    end else if (io_mem2rb_valid) begin // @[playground/src/noop/writeback.scala 56:30]
      if (io_mem2rb_special != 2'h0 | io_mem2rb_recov & ~io_mem2rb_excep_en) begin // @[playground/src/noop/writeback.scala 67:88]
        forceJmp_seq_pc <= _forceJmp_seq_pc_T_1; // @[playground/src/noop/writeback.scala 69:33]
      end
    end
    if (reset) begin // @[playground/src/noop/writeback.scala 25:30]
      forceJmp_valid <= 1'h0; // @[playground/src/noop/writeback.scala 25:30]
    end else begin
      forceJmp_valid <= _GEN_19;
    end
    if (reset) begin // @[playground/src/noop/writeback.scala 26:30]
      tlb_r <= 1'h0; // @[playground/src/noop/writeback.scala 26:30]
    end else begin
      tlb_r <= _GEN_22;
    end
    if (reset) begin // @[playground/src/noop/writeback.scala 27:30]
      cache_r <= 1'h0; // @[playground/src/noop/writeback.scala 27:30]
    end else begin
      cache_r <= _GEN_21;
    end
    if (reset) begin // @[playground/src/noop/writeback.scala 28:30]
      valid_r <= 1'h0; // @[playground/src/noop/writeback.scala 28:30]
    end else begin
      valid_r <= io_mem2rb_valid;
    end
    if (reset) begin // @[playground/src/noop/writeback.scala 29:30]
      excep_r_cause <= 64'h0; // @[playground/src/noop/writeback.scala 29:30]
    end else if (io_mem2rb_valid) begin // @[playground/src/noop/writeback.scala 56:30]
      excep_r_cause <= io_mem2rb_excep_cause; // @[playground/src/noop/writeback.scala 65:21]
    end
    if (reset) begin // @[playground/src/noop/writeback.scala 29:30]
      excep_r_en <= 1'h0; // @[playground/src/noop/writeback.scala 29:30]
    end else begin
      excep_r_en <= _GEN_10;
    end
    if (reset) begin // @[playground/src/noop/writeback.scala 29:30]
      excep_r_pc <= 64'h0; // @[playground/src/noop/writeback.scala 29:30]
    end else if (io_mem2rb_valid) begin // @[playground/src/noop/writeback.scala 56:30]
      excep_r_pc <= io_mem2rb_excep_pc; // @[playground/src/noop/writeback.scala 65:21]
    end
    if (reset) begin // @[playground/src/noop/writeback.scala 29:30]
      excep_r_etype <= 2'h0; // @[playground/src/noop/writeback.scala 29:30]
    end else if (io_mem2rb_valid) begin // @[playground/src/noop/writeback.scala 56:30]
      excep_r_etype <= io_mem2rb_excep_etype; // @[playground/src/noop/writeback.scala 65:21]
    end
    if (reset) begin // @[playground/src/noop/writeback.scala 30:30]
      rcsr_id_r <= 12'h0; // @[playground/src/noop/writeback.scala 30:30]
    end else if (io_mem2rb_valid) begin // @[playground/src/noop/writeback.scala 56:30]
      rcsr_id_r <= io_mem2rb_rcsr_id; // @[playground/src/noop/writeback.scala 66:25]
    end else begin
      rcsr_id_r <= 12'h0; // @[playground/src/noop/writeback.scala 36:21]
    end
    if (reset) begin // @[playground/src/noop/writeback.scala 40:30]
      inst_r <= 32'h0; // @[playground/src/noop/writeback.scala 40:30]
    end else if (io_mem2rb_valid) begin // @[playground/src/noop/writeback.scala 56:30]
      inst_r <= io_mem2rb_inst; // @[playground/src/noop/writeback.scala 62:21]
    end
    if (reset) begin // @[playground/src/noop/writeback.scala 41:30]
      pc_r <= 64'h0; // @[playground/src/noop/writeback.scala 41:30]
    end else if (io_mem2rb_valid) begin // @[playground/src/noop/writeback.scala 56:30]
      pc_r <= io_mem2rb_pc; // @[playground/src/noop/writeback.scala 63:21]
    end
    is_mmio_r <= io_mem2rb_is_mmio; // @[playground/src/noop/writeback.scala 78:30]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  recov_r = _RAND_0[0:0];
  _RAND_1 = {2{`RANDOM}};
  forceJmp_seq_pc = _RAND_1[63:0];
  _RAND_2 = {1{`RANDOM}};
  forceJmp_valid = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  tlb_r = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  cache_r = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  valid_r = _RAND_5[0:0];
  _RAND_6 = {2{`RANDOM}};
  excep_r_cause = _RAND_6[63:0];
  _RAND_7 = {1{`RANDOM}};
  excep_r_en = _RAND_7[0:0];
  _RAND_8 = {2{`RANDOM}};
  excep_r_pc = _RAND_8[63:0];
  _RAND_9 = {1{`RANDOM}};
  excep_r_etype = _RAND_9[1:0];
  _RAND_10 = {1{`RANDOM}};
  rcsr_id_r = _RAND_10[11:0];
  _RAND_11 = {1{`RANDOM}};
  inst_r = _RAND_11[31:0];
  _RAND_12 = {2{`RANDOM}};
  pc_r = _RAND_12[63:0];
  _RAND_13 = {1{`RANDOM}};
  is_mmio_r = _RAND_13[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Regs(
  input         clock,
  input         reset,
  input  [4:0]  io_rs1_id, // @[playground/src/noop/regs.scala 10:16]
  output [63:0] io_rs1_data, // @[playground/src/noop/regs.scala 10:16]
  input  [4:0]  io_rs2_id, // @[playground/src/noop/regs.scala 10:16]
  output [63:0] io_rs2_data, // @[playground/src/noop/regs.scala 10:16]
  input  [4:0]  io_dst_id, // @[playground/src/noop/regs.scala 10:16]
  input  [63:0] io_dst_data, // @[playground/src/noop/regs.scala 10:16]
  input         io_dst_en // @[playground/src/noop/regs.scala 10:16]
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [63:0] _RAND_12;
  reg [63:0] _RAND_13;
  reg [63:0] _RAND_14;
  reg [63:0] _RAND_15;
  reg [63:0] _RAND_16;
  reg [63:0] _RAND_17;
  reg [63:0] _RAND_18;
  reg [63:0] _RAND_19;
  reg [63:0] _RAND_20;
  reg [63:0] _RAND_21;
  reg [63:0] _RAND_22;
  reg [63:0] _RAND_23;
  reg [63:0] _RAND_24;
  reg [63:0] _RAND_25;
  reg [63:0] _RAND_26;
  reg [63:0] _RAND_27;
  reg [63:0] _RAND_28;
  reg [63:0] _RAND_29;
  reg [63:0] _RAND_30;
  reg [63:0] _RAND_31;
`endif // RANDOMIZE_REG_INIT
  wire [2047:0] updateRegs_regs_data; // @[playground/src/noop/regs.scala 21:28]
  wire  updateRegs_clock; // @[playground/src/noop/regs.scala 21:28]
  reg [63:0] regs_0; // @[playground/src/noop/regs.scala 15:23]
  reg [63:0] regs_1; // @[playground/src/noop/regs.scala 15:23]
  reg [63:0] regs_2; // @[playground/src/noop/regs.scala 15:23]
  reg [63:0] regs_3; // @[playground/src/noop/regs.scala 15:23]
  reg [63:0] regs_4; // @[playground/src/noop/regs.scala 15:23]
  reg [63:0] regs_5; // @[playground/src/noop/regs.scala 15:23]
  reg [63:0] regs_6; // @[playground/src/noop/regs.scala 15:23]
  reg [63:0] regs_7; // @[playground/src/noop/regs.scala 15:23]
  reg [63:0] regs_8; // @[playground/src/noop/regs.scala 15:23]
  reg [63:0] regs_9; // @[playground/src/noop/regs.scala 15:23]
  reg [63:0] regs_10; // @[playground/src/noop/regs.scala 15:23]
  reg [63:0] regs_11; // @[playground/src/noop/regs.scala 15:23]
  reg [63:0] regs_12; // @[playground/src/noop/regs.scala 15:23]
  reg [63:0] regs_13; // @[playground/src/noop/regs.scala 15:23]
  reg [63:0] regs_14; // @[playground/src/noop/regs.scala 15:23]
  reg [63:0] regs_15; // @[playground/src/noop/regs.scala 15:23]
  reg [63:0] regs_16; // @[playground/src/noop/regs.scala 15:23]
  reg [63:0] regs_17; // @[playground/src/noop/regs.scala 15:23]
  reg [63:0] regs_18; // @[playground/src/noop/regs.scala 15:23]
  reg [63:0] regs_19; // @[playground/src/noop/regs.scala 15:23]
  reg [63:0] regs_20; // @[playground/src/noop/regs.scala 15:23]
  reg [63:0] regs_21; // @[playground/src/noop/regs.scala 15:23]
  reg [63:0] regs_22; // @[playground/src/noop/regs.scala 15:23]
  reg [63:0] regs_23; // @[playground/src/noop/regs.scala 15:23]
  reg [63:0] regs_24; // @[playground/src/noop/regs.scala 15:23]
  reg [63:0] regs_25; // @[playground/src/noop/regs.scala 15:23]
  reg [63:0] regs_26; // @[playground/src/noop/regs.scala 15:23]
  reg [63:0] regs_27; // @[playground/src/noop/regs.scala 15:23]
  reg [63:0] regs_28; // @[playground/src/noop/regs.scala 15:23]
  reg [63:0] regs_29; // @[playground/src/noop/regs.scala 15:23]
  reg [63:0] regs_30; // @[playground/src/noop/regs.scala 15:23]
  reg [63:0] regs_31; // @[playground/src/noop/regs.scala 15:23]
  wire [63:0] _GEN_1 = 5'h1 == io_rs1_id ? regs_1 : regs_0; // @[playground/src/noop/regs.scala 16:{17,17}]
  wire [63:0] _GEN_2 = 5'h2 == io_rs1_id ? regs_2 : _GEN_1; // @[playground/src/noop/regs.scala 16:{17,17}]
  wire [63:0] _GEN_3 = 5'h3 == io_rs1_id ? regs_3 : _GEN_2; // @[playground/src/noop/regs.scala 16:{17,17}]
  wire [63:0] _GEN_4 = 5'h4 == io_rs1_id ? regs_4 : _GEN_3; // @[playground/src/noop/regs.scala 16:{17,17}]
  wire [63:0] _GEN_5 = 5'h5 == io_rs1_id ? regs_5 : _GEN_4; // @[playground/src/noop/regs.scala 16:{17,17}]
  wire [63:0] _GEN_6 = 5'h6 == io_rs1_id ? regs_6 : _GEN_5; // @[playground/src/noop/regs.scala 16:{17,17}]
  wire [63:0] _GEN_7 = 5'h7 == io_rs1_id ? regs_7 : _GEN_6; // @[playground/src/noop/regs.scala 16:{17,17}]
  wire [63:0] _GEN_8 = 5'h8 == io_rs1_id ? regs_8 : _GEN_7; // @[playground/src/noop/regs.scala 16:{17,17}]
  wire [63:0] _GEN_9 = 5'h9 == io_rs1_id ? regs_9 : _GEN_8; // @[playground/src/noop/regs.scala 16:{17,17}]
  wire [63:0] _GEN_10 = 5'ha == io_rs1_id ? regs_10 : _GEN_9; // @[playground/src/noop/regs.scala 16:{17,17}]
  wire [63:0] _GEN_11 = 5'hb == io_rs1_id ? regs_11 : _GEN_10; // @[playground/src/noop/regs.scala 16:{17,17}]
  wire [63:0] _GEN_12 = 5'hc == io_rs1_id ? regs_12 : _GEN_11; // @[playground/src/noop/regs.scala 16:{17,17}]
  wire [63:0] _GEN_13 = 5'hd == io_rs1_id ? regs_13 : _GEN_12; // @[playground/src/noop/regs.scala 16:{17,17}]
  wire [63:0] _GEN_14 = 5'he == io_rs1_id ? regs_14 : _GEN_13; // @[playground/src/noop/regs.scala 16:{17,17}]
  wire [63:0] _GEN_15 = 5'hf == io_rs1_id ? regs_15 : _GEN_14; // @[playground/src/noop/regs.scala 16:{17,17}]
  wire [63:0] _GEN_16 = 5'h10 == io_rs1_id ? regs_16 : _GEN_15; // @[playground/src/noop/regs.scala 16:{17,17}]
  wire [63:0] _GEN_17 = 5'h11 == io_rs1_id ? regs_17 : _GEN_16; // @[playground/src/noop/regs.scala 16:{17,17}]
  wire [63:0] _GEN_18 = 5'h12 == io_rs1_id ? regs_18 : _GEN_17; // @[playground/src/noop/regs.scala 16:{17,17}]
  wire [63:0] _GEN_19 = 5'h13 == io_rs1_id ? regs_19 : _GEN_18; // @[playground/src/noop/regs.scala 16:{17,17}]
  wire [63:0] _GEN_20 = 5'h14 == io_rs1_id ? regs_20 : _GEN_19; // @[playground/src/noop/regs.scala 16:{17,17}]
  wire [63:0] _GEN_21 = 5'h15 == io_rs1_id ? regs_21 : _GEN_20; // @[playground/src/noop/regs.scala 16:{17,17}]
  wire [63:0] _GEN_22 = 5'h16 == io_rs1_id ? regs_22 : _GEN_21; // @[playground/src/noop/regs.scala 16:{17,17}]
  wire [63:0] _GEN_23 = 5'h17 == io_rs1_id ? regs_23 : _GEN_22; // @[playground/src/noop/regs.scala 16:{17,17}]
  wire [63:0] _GEN_24 = 5'h18 == io_rs1_id ? regs_24 : _GEN_23; // @[playground/src/noop/regs.scala 16:{17,17}]
  wire [63:0] _GEN_25 = 5'h19 == io_rs1_id ? regs_25 : _GEN_24; // @[playground/src/noop/regs.scala 16:{17,17}]
  wire [63:0] _GEN_26 = 5'h1a == io_rs1_id ? regs_26 : _GEN_25; // @[playground/src/noop/regs.scala 16:{17,17}]
  wire [63:0] _GEN_27 = 5'h1b == io_rs1_id ? regs_27 : _GEN_26; // @[playground/src/noop/regs.scala 16:{17,17}]
  wire [63:0] _GEN_28 = 5'h1c == io_rs1_id ? regs_28 : _GEN_27; // @[playground/src/noop/regs.scala 16:{17,17}]
  wire [63:0] _GEN_29 = 5'h1d == io_rs1_id ? regs_29 : _GEN_28; // @[playground/src/noop/regs.scala 16:{17,17}]
  wire [63:0] _GEN_30 = 5'h1e == io_rs1_id ? regs_30 : _GEN_29; // @[playground/src/noop/regs.scala 16:{17,17}]
  wire [63:0] _GEN_33 = 5'h1 == io_rs2_id ? regs_1 : regs_0; // @[playground/src/noop/regs.scala 17:{17,17}]
  wire [63:0] _GEN_34 = 5'h2 == io_rs2_id ? regs_2 : _GEN_33; // @[playground/src/noop/regs.scala 17:{17,17}]
  wire [63:0] _GEN_35 = 5'h3 == io_rs2_id ? regs_3 : _GEN_34; // @[playground/src/noop/regs.scala 17:{17,17}]
  wire [63:0] _GEN_36 = 5'h4 == io_rs2_id ? regs_4 : _GEN_35; // @[playground/src/noop/regs.scala 17:{17,17}]
  wire [63:0] _GEN_37 = 5'h5 == io_rs2_id ? regs_5 : _GEN_36; // @[playground/src/noop/regs.scala 17:{17,17}]
  wire [63:0] _GEN_38 = 5'h6 == io_rs2_id ? regs_6 : _GEN_37; // @[playground/src/noop/regs.scala 17:{17,17}]
  wire [63:0] _GEN_39 = 5'h7 == io_rs2_id ? regs_7 : _GEN_38; // @[playground/src/noop/regs.scala 17:{17,17}]
  wire [63:0] _GEN_40 = 5'h8 == io_rs2_id ? regs_8 : _GEN_39; // @[playground/src/noop/regs.scala 17:{17,17}]
  wire [63:0] _GEN_41 = 5'h9 == io_rs2_id ? regs_9 : _GEN_40; // @[playground/src/noop/regs.scala 17:{17,17}]
  wire [63:0] _GEN_42 = 5'ha == io_rs2_id ? regs_10 : _GEN_41; // @[playground/src/noop/regs.scala 17:{17,17}]
  wire [63:0] _GEN_43 = 5'hb == io_rs2_id ? regs_11 : _GEN_42; // @[playground/src/noop/regs.scala 17:{17,17}]
  wire [63:0] _GEN_44 = 5'hc == io_rs2_id ? regs_12 : _GEN_43; // @[playground/src/noop/regs.scala 17:{17,17}]
  wire [63:0] _GEN_45 = 5'hd == io_rs2_id ? regs_13 : _GEN_44; // @[playground/src/noop/regs.scala 17:{17,17}]
  wire [63:0] _GEN_46 = 5'he == io_rs2_id ? regs_14 : _GEN_45; // @[playground/src/noop/regs.scala 17:{17,17}]
  wire [63:0] _GEN_47 = 5'hf == io_rs2_id ? regs_15 : _GEN_46; // @[playground/src/noop/regs.scala 17:{17,17}]
  wire [63:0] _GEN_48 = 5'h10 == io_rs2_id ? regs_16 : _GEN_47; // @[playground/src/noop/regs.scala 17:{17,17}]
  wire [63:0] _GEN_49 = 5'h11 == io_rs2_id ? regs_17 : _GEN_48; // @[playground/src/noop/regs.scala 17:{17,17}]
  wire [63:0] _GEN_50 = 5'h12 == io_rs2_id ? regs_18 : _GEN_49; // @[playground/src/noop/regs.scala 17:{17,17}]
  wire [63:0] _GEN_51 = 5'h13 == io_rs2_id ? regs_19 : _GEN_50; // @[playground/src/noop/regs.scala 17:{17,17}]
  wire [63:0] _GEN_52 = 5'h14 == io_rs2_id ? regs_20 : _GEN_51; // @[playground/src/noop/regs.scala 17:{17,17}]
  wire [63:0] _GEN_53 = 5'h15 == io_rs2_id ? regs_21 : _GEN_52; // @[playground/src/noop/regs.scala 17:{17,17}]
  wire [63:0] _GEN_54 = 5'h16 == io_rs2_id ? regs_22 : _GEN_53; // @[playground/src/noop/regs.scala 17:{17,17}]
  wire [63:0] _GEN_55 = 5'h17 == io_rs2_id ? regs_23 : _GEN_54; // @[playground/src/noop/regs.scala 17:{17,17}]
  wire [63:0] _GEN_56 = 5'h18 == io_rs2_id ? regs_24 : _GEN_55; // @[playground/src/noop/regs.scala 17:{17,17}]
  wire [63:0] _GEN_57 = 5'h19 == io_rs2_id ? regs_25 : _GEN_56; // @[playground/src/noop/regs.scala 17:{17,17}]
  wire [63:0] _GEN_58 = 5'h1a == io_rs2_id ? regs_26 : _GEN_57; // @[playground/src/noop/regs.scala 17:{17,17}]
  wire [63:0] _GEN_59 = 5'h1b == io_rs2_id ? regs_27 : _GEN_58; // @[playground/src/noop/regs.scala 17:{17,17}]
  wire [63:0] _GEN_60 = 5'h1c == io_rs2_id ? regs_28 : _GEN_59; // @[playground/src/noop/regs.scala 17:{17,17}]
  wire [63:0] _GEN_61 = 5'h1d == io_rs2_id ? regs_29 : _GEN_60; // @[playground/src/noop/regs.scala 17:{17,17}]
  wire [63:0] _GEN_62 = 5'h1e == io_rs2_id ? regs_30 : _GEN_61; // @[playground/src/noop/regs.scala 17:{17,17}]
  wire [511:0] updateRegs_io_regs_data_lo_lo = {regs_7,regs_6,regs_5,regs_4,regs_3,regs_2,regs_1,regs_0}; // @[playground/src/noop/regs.scala 22:37]
  wire [1023:0] updateRegs_io_regs_data_lo = {regs_15,regs_14,regs_13,regs_12,regs_11,regs_10,regs_9,regs_8,
    updateRegs_io_regs_data_lo_lo}; // @[playground/src/noop/regs.scala 22:37]
  wire [511:0] updateRegs_io_regs_data_hi_lo = {regs_23,regs_22,regs_21,regs_20,regs_19,regs_18,regs_17,regs_16}; // @[playground/src/noop/regs.scala 22:37]
  wire [1023:0] updateRegs_io_regs_data_hi = {regs_31,regs_30,regs_29,regs_28,regs_27,regs_26,regs_25,regs_24,
    updateRegs_io_regs_data_hi_lo}; // @[playground/src/noop/regs.scala 22:37]
  UpdateRegs updateRegs ( // @[playground/src/noop/regs.scala 21:28]
    .regs_data(updateRegs_regs_data),
    .clock(updateRegs_clock)
  );
  assign io_rs1_data = 5'h1f == io_rs1_id ? regs_31 : _GEN_30; // @[playground/src/noop/regs.scala 16:{17,17}]
  assign io_rs2_data = 5'h1f == io_rs2_id ? regs_31 : _GEN_62; // @[playground/src/noop/regs.scala 17:{17,17}]
  assign updateRegs_regs_data = {updateRegs_io_regs_data_hi,updateRegs_io_regs_data_lo}; // @[playground/src/noop/regs.scala 22:37]
  assign updateRegs_clock = clock; // @[playground/src/noop/regs.scala 23:25]
  always @(posedge clock) begin
    if (reset) begin // @[playground/src/noop/regs.scala 15:23]
      regs_0 <= 64'h0; // @[playground/src/noop/regs.scala 15:23]
    end else if (io_dst_en & io_dst_id != 5'h0) begin // @[playground/src/noop/regs.scala 18:41]
      if (5'h0 == io_dst_id) begin // @[playground/src/noop/regs.scala 19:25]
        regs_0 <= io_dst_data; // @[playground/src/noop/regs.scala 19:25]
      end
    end
    if (reset) begin // @[playground/src/noop/regs.scala 15:23]
      regs_1 <= 64'h0; // @[playground/src/noop/regs.scala 15:23]
    end else if (io_dst_en & io_dst_id != 5'h0) begin // @[playground/src/noop/regs.scala 18:41]
      if (5'h1 == io_dst_id) begin // @[playground/src/noop/regs.scala 19:25]
        regs_1 <= io_dst_data; // @[playground/src/noop/regs.scala 19:25]
      end
    end
    if (reset) begin // @[playground/src/noop/regs.scala 15:23]
      regs_2 <= 64'h0; // @[playground/src/noop/regs.scala 15:23]
    end else if (io_dst_en & io_dst_id != 5'h0) begin // @[playground/src/noop/regs.scala 18:41]
      if (5'h2 == io_dst_id) begin // @[playground/src/noop/regs.scala 19:25]
        regs_2 <= io_dst_data; // @[playground/src/noop/regs.scala 19:25]
      end
    end
    if (reset) begin // @[playground/src/noop/regs.scala 15:23]
      regs_3 <= 64'h0; // @[playground/src/noop/regs.scala 15:23]
    end else if (io_dst_en & io_dst_id != 5'h0) begin // @[playground/src/noop/regs.scala 18:41]
      if (5'h3 == io_dst_id) begin // @[playground/src/noop/regs.scala 19:25]
        regs_3 <= io_dst_data; // @[playground/src/noop/regs.scala 19:25]
      end
    end
    if (reset) begin // @[playground/src/noop/regs.scala 15:23]
      regs_4 <= 64'h0; // @[playground/src/noop/regs.scala 15:23]
    end else if (io_dst_en & io_dst_id != 5'h0) begin // @[playground/src/noop/regs.scala 18:41]
      if (5'h4 == io_dst_id) begin // @[playground/src/noop/regs.scala 19:25]
        regs_4 <= io_dst_data; // @[playground/src/noop/regs.scala 19:25]
      end
    end
    if (reset) begin // @[playground/src/noop/regs.scala 15:23]
      regs_5 <= 64'h0; // @[playground/src/noop/regs.scala 15:23]
    end else if (io_dst_en & io_dst_id != 5'h0) begin // @[playground/src/noop/regs.scala 18:41]
      if (5'h5 == io_dst_id) begin // @[playground/src/noop/regs.scala 19:25]
        regs_5 <= io_dst_data; // @[playground/src/noop/regs.scala 19:25]
      end
    end
    if (reset) begin // @[playground/src/noop/regs.scala 15:23]
      regs_6 <= 64'h0; // @[playground/src/noop/regs.scala 15:23]
    end else if (io_dst_en & io_dst_id != 5'h0) begin // @[playground/src/noop/regs.scala 18:41]
      if (5'h6 == io_dst_id) begin // @[playground/src/noop/regs.scala 19:25]
        regs_6 <= io_dst_data; // @[playground/src/noop/regs.scala 19:25]
      end
    end
    if (reset) begin // @[playground/src/noop/regs.scala 15:23]
      regs_7 <= 64'h0; // @[playground/src/noop/regs.scala 15:23]
    end else if (io_dst_en & io_dst_id != 5'h0) begin // @[playground/src/noop/regs.scala 18:41]
      if (5'h7 == io_dst_id) begin // @[playground/src/noop/regs.scala 19:25]
        regs_7 <= io_dst_data; // @[playground/src/noop/regs.scala 19:25]
      end
    end
    if (reset) begin // @[playground/src/noop/regs.scala 15:23]
      regs_8 <= 64'h0; // @[playground/src/noop/regs.scala 15:23]
    end else if (io_dst_en & io_dst_id != 5'h0) begin // @[playground/src/noop/regs.scala 18:41]
      if (5'h8 == io_dst_id) begin // @[playground/src/noop/regs.scala 19:25]
        regs_8 <= io_dst_data; // @[playground/src/noop/regs.scala 19:25]
      end
    end
    if (reset) begin // @[playground/src/noop/regs.scala 15:23]
      regs_9 <= 64'h0; // @[playground/src/noop/regs.scala 15:23]
    end else if (io_dst_en & io_dst_id != 5'h0) begin // @[playground/src/noop/regs.scala 18:41]
      if (5'h9 == io_dst_id) begin // @[playground/src/noop/regs.scala 19:25]
        regs_9 <= io_dst_data; // @[playground/src/noop/regs.scala 19:25]
      end
    end
    if (reset) begin // @[playground/src/noop/regs.scala 15:23]
      regs_10 <= 64'h0; // @[playground/src/noop/regs.scala 15:23]
    end else if (io_dst_en & io_dst_id != 5'h0) begin // @[playground/src/noop/regs.scala 18:41]
      if (5'ha == io_dst_id) begin // @[playground/src/noop/regs.scala 19:25]
        regs_10 <= io_dst_data; // @[playground/src/noop/regs.scala 19:25]
      end
    end
    if (reset) begin // @[playground/src/noop/regs.scala 15:23]
      regs_11 <= 64'h0; // @[playground/src/noop/regs.scala 15:23]
    end else if (io_dst_en & io_dst_id != 5'h0) begin // @[playground/src/noop/regs.scala 18:41]
      if (5'hb == io_dst_id) begin // @[playground/src/noop/regs.scala 19:25]
        regs_11 <= io_dst_data; // @[playground/src/noop/regs.scala 19:25]
      end
    end
    if (reset) begin // @[playground/src/noop/regs.scala 15:23]
      regs_12 <= 64'h0; // @[playground/src/noop/regs.scala 15:23]
    end else if (io_dst_en & io_dst_id != 5'h0) begin // @[playground/src/noop/regs.scala 18:41]
      if (5'hc == io_dst_id) begin // @[playground/src/noop/regs.scala 19:25]
        regs_12 <= io_dst_data; // @[playground/src/noop/regs.scala 19:25]
      end
    end
    if (reset) begin // @[playground/src/noop/regs.scala 15:23]
      regs_13 <= 64'h0; // @[playground/src/noop/regs.scala 15:23]
    end else if (io_dst_en & io_dst_id != 5'h0) begin // @[playground/src/noop/regs.scala 18:41]
      if (5'hd == io_dst_id) begin // @[playground/src/noop/regs.scala 19:25]
        regs_13 <= io_dst_data; // @[playground/src/noop/regs.scala 19:25]
      end
    end
    if (reset) begin // @[playground/src/noop/regs.scala 15:23]
      regs_14 <= 64'h0; // @[playground/src/noop/regs.scala 15:23]
    end else if (io_dst_en & io_dst_id != 5'h0) begin // @[playground/src/noop/regs.scala 18:41]
      if (5'he == io_dst_id) begin // @[playground/src/noop/regs.scala 19:25]
        regs_14 <= io_dst_data; // @[playground/src/noop/regs.scala 19:25]
      end
    end
    if (reset) begin // @[playground/src/noop/regs.scala 15:23]
      regs_15 <= 64'h0; // @[playground/src/noop/regs.scala 15:23]
    end else if (io_dst_en & io_dst_id != 5'h0) begin // @[playground/src/noop/regs.scala 18:41]
      if (5'hf == io_dst_id) begin // @[playground/src/noop/regs.scala 19:25]
        regs_15 <= io_dst_data; // @[playground/src/noop/regs.scala 19:25]
      end
    end
    if (reset) begin // @[playground/src/noop/regs.scala 15:23]
      regs_16 <= 64'h0; // @[playground/src/noop/regs.scala 15:23]
    end else if (io_dst_en & io_dst_id != 5'h0) begin // @[playground/src/noop/regs.scala 18:41]
      if (5'h10 == io_dst_id) begin // @[playground/src/noop/regs.scala 19:25]
        regs_16 <= io_dst_data; // @[playground/src/noop/regs.scala 19:25]
      end
    end
    if (reset) begin // @[playground/src/noop/regs.scala 15:23]
      regs_17 <= 64'h0; // @[playground/src/noop/regs.scala 15:23]
    end else if (io_dst_en & io_dst_id != 5'h0) begin // @[playground/src/noop/regs.scala 18:41]
      if (5'h11 == io_dst_id) begin // @[playground/src/noop/regs.scala 19:25]
        regs_17 <= io_dst_data; // @[playground/src/noop/regs.scala 19:25]
      end
    end
    if (reset) begin // @[playground/src/noop/regs.scala 15:23]
      regs_18 <= 64'h0; // @[playground/src/noop/regs.scala 15:23]
    end else if (io_dst_en & io_dst_id != 5'h0) begin // @[playground/src/noop/regs.scala 18:41]
      if (5'h12 == io_dst_id) begin // @[playground/src/noop/regs.scala 19:25]
        regs_18 <= io_dst_data; // @[playground/src/noop/regs.scala 19:25]
      end
    end
    if (reset) begin // @[playground/src/noop/regs.scala 15:23]
      regs_19 <= 64'h0; // @[playground/src/noop/regs.scala 15:23]
    end else if (io_dst_en & io_dst_id != 5'h0) begin // @[playground/src/noop/regs.scala 18:41]
      if (5'h13 == io_dst_id) begin // @[playground/src/noop/regs.scala 19:25]
        regs_19 <= io_dst_data; // @[playground/src/noop/regs.scala 19:25]
      end
    end
    if (reset) begin // @[playground/src/noop/regs.scala 15:23]
      regs_20 <= 64'h0; // @[playground/src/noop/regs.scala 15:23]
    end else if (io_dst_en & io_dst_id != 5'h0) begin // @[playground/src/noop/regs.scala 18:41]
      if (5'h14 == io_dst_id) begin // @[playground/src/noop/regs.scala 19:25]
        regs_20 <= io_dst_data; // @[playground/src/noop/regs.scala 19:25]
      end
    end
    if (reset) begin // @[playground/src/noop/regs.scala 15:23]
      regs_21 <= 64'h0; // @[playground/src/noop/regs.scala 15:23]
    end else if (io_dst_en & io_dst_id != 5'h0) begin // @[playground/src/noop/regs.scala 18:41]
      if (5'h15 == io_dst_id) begin // @[playground/src/noop/regs.scala 19:25]
        regs_21 <= io_dst_data; // @[playground/src/noop/regs.scala 19:25]
      end
    end
    if (reset) begin // @[playground/src/noop/regs.scala 15:23]
      regs_22 <= 64'h0; // @[playground/src/noop/regs.scala 15:23]
    end else if (io_dst_en & io_dst_id != 5'h0) begin // @[playground/src/noop/regs.scala 18:41]
      if (5'h16 == io_dst_id) begin // @[playground/src/noop/regs.scala 19:25]
        regs_22 <= io_dst_data; // @[playground/src/noop/regs.scala 19:25]
      end
    end
    if (reset) begin // @[playground/src/noop/regs.scala 15:23]
      regs_23 <= 64'h0; // @[playground/src/noop/regs.scala 15:23]
    end else if (io_dst_en & io_dst_id != 5'h0) begin // @[playground/src/noop/regs.scala 18:41]
      if (5'h17 == io_dst_id) begin // @[playground/src/noop/regs.scala 19:25]
        regs_23 <= io_dst_data; // @[playground/src/noop/regs.scala 19:25]
      end
    end
    if (reset) begin // @[playground/src/noop/regs.scala 15:23]
      regs_24 <= 64'h0; // @[playground/src/noop/regs.scala 15:23]
    end else if (io_dst_en & io_dst_id != 5'h0) begin // @[playground/src/noop/regs.scala 18:41]
      if (5'h18 == io_dst_id) begin // @[playground/src/noop/regs.scala 19:25]
        regs_24 <= io_dst_data; // @[playground/src/noop/regs.scala 19:25]
      end
    end
    if (reset) begin // @[playground/src/noop/regs.scala 15:23]
      regs_25 <= 64'h0; // @[playground/src/noop/regs.scala 15:23]
    end else if (io_dst_en & io_dst_id != 5'h0) begin // @[playground/src/noop/regs.scala 18:41]
      if (5'h19 == io_dst_id) begin // @[playground/src/noop/regs.scala 19:25]
        regs_25 <= io_dst_data; // @[playground/src/noop/regs.scala 19:25]
      end
    end
    if (reset) begin // @[playground/src/noop/regs.scala 15:23]
      regs_26 <= 64'h0; // @[playground/src/noop/regs.scala 15:23]
    end else if (io_dst_en & io_dst_id != 5'h0) begin // @[playground/src/noop/regs.scala 18:41]
      if (5'h1a == io_dst_id) begin // @[playground/src/noop/regs.scala 19:25]
        regs_26 <= io_dst_data; // @[playground/src/noop/regs.scala 19:25]
      end
    end
    if (reset) begin // @[playground/src/noop/regs.scala 15:23]
      regs_27 <= 64'h0; // @[playground/src/noop/regs.scala 15:23]
    end else if (io_dst_en & io_dst_id != 5'h0) begin // @[playground/src/noop/regs.scala 18:41]
      if (5'h1b == io_dst_id) begin // @[playground/src/noop/regs.scala 19:25]
        regs_27 <= io_dst_data; // @[playground/src/noop/regs.scala 19:25]
      end
    end
    if (reset) begin // @[playground/src/noop/regs.scala 15:23]
      regs_28 <= 64'h0; // @[playground/src/noop/regs.scala 15:23]
    end else if (io_dst_en & io_dst_id != 5'h0) begin // @[playground/src/noop/regs.scala 18:41]
      if (5'h1c == io_dst_id) begin // @[playground/src/noop/regs.scala 19:25]
        regs_28 <= io_dst_data; // @[playground/src/noop/regs.scala 19:25]
      end
    end
    if (reset) begin // @[playground/src/noop/regs.scala 15:23]
      regs_29 <= 64'h0; // @[playground/src/noop/regs.scala 15:23]
    end else if (io_dst_en & io_dst_id != 5'h0) begin // @[playground/src/noop/regs.scala 18:41]
      if (5'h1d == io_dst_id) begin // @[playground/src/noop/regs.scala 19:25]
        regs_29 <= io_dst_data; // @[playground/src/noop/regs.scala 19:25]
      end
    end
    if (reset) begin // @[playground/src/noop/regs.scala 15:23]
      regs_30 <= 64'h0; // @[playground/src/noop/regs.scala 15:23]
    end else if (io_dst_en & io_dst_id != 5'h0) begin // @[playground/src/noop/regs.scala 18:41]
      if (5'h1e == io_dst_id) begin // @[playground/src/noop/regs.scala 19:25]
        regs_30 <= io_dst_data; // @[playground/src/noop/regs.scala 19:25]
      end
    end
    if (reset) begin // @[playground/src/noop/regs.scala 15:23]
      regs_31 <= 64'h0; // @[playground/src/noop/regs.scala 15:23]
    end else if (io_dst_en & io_dst_id != 5'h0) begin // @[playground/src/noop/regs.scala 18:41]
      if (5'h1f == io_dst_id) begin // @[playground/src/noop/regs.scala 19:25]
        regs_31 <= io_dst_data; // @[playground/src/noop/regs.scala 19:25]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  regs_0 = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  regs_1 = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  regs_2 = _RAND_2[63:0];
  _RAND_3 = {2{`RANDOM}};
  regs_3 = _RAND_3[63:0];
  _RAND_4 = {2{`RANDOM}};
  regs_4 = _RAND_4[63:0];
  _RAND_5 = {2{`RANDOM}};
  regs_5 = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  regs_6 = _RAND_6[63:0];
  _RAND_7 = {2{`RANDOM}};
  regs_7 = _RAND_7[63:0];
  _RAND_8 = {2{`RANDOM}};
  regs_8 = _RAND_8[63:0];
  _RAND_9 = {2{`RANDOM}};
  regs_9 = _RAND_9[63:0];
  _RAND_10 = {2{`RANDOM}};
  regs_10 = _RAND_10[63:0];
  _RAND_11 = {2{`RANDOM}};
  regs_11 = _RAND_11[63:0];
  _RAND_12 = {2{`RANDOM}};
  regs_12 = _RAND_12[63:0];
  _RAND_13 = {2{`RANDOM}};
  regs_13 = _RAND_13[63:0];
  _RAND_14 = {2{`RANDOM}};
  regs_14 = _RAND_14[63:0];
  _RAND_15 = {2{`RANDOM}};
  regs_15 = _RAND_15[63:0];
  _RAND_16 = {2{`RANDOM}};
  regs_16 = _RAND_16[63:0];
  _RAND_17 = {2{`RANDOM}};
  regs_17 = _RAND_17[63:0];
  _RAND_18 = {2{`RANDOM}};
  regs_18 = _RAND_18[63:0];
  _RAND_19 = {2{`RANDOM}};
  regs_19 = _RAND_19[63:0];
  _RAND_20 = {2{`RANDOM}};
  regs_20 = _RAND_20[63:0];
  _RAND_21 = {2{`RANDOM}};
  regs_21 = _RAND_21[63:0];
  _RAND_22 = {2{`RANDOM}};
  regs_22 = _RAND_22[63:0];
  _RAND_23 = {2{`RANDOM}};
  regs_23 = _RAND_23[63:0];
  _RAND_24 = {2{`RANDOM}};
  regs_24 = _RAND_24[63:0];
  _RAND_25 = {2{`RANDOM}};
  regs_25 = _RAND_25[63:0];
  _RAND_26 = {2{`RANDOM}};
  regs_26 = _RAND_26[63:0];
  _RAND_27 = {2{`RANDOM}};
  regs_27 = _RAND_27[63:0];
  _RAND_28 = {2{`RANDOM}};
  regs_28 = _RAND_28[63:0];
  _RAND_29 = {2{`RANDOM}};
  regs_29 = _RAND_29[63:0];
  _RAND_30 = {2{`RANDOM}};
  regs_30 = _RAND_30[63:0];
  _RAND_31 = {2{`RANDOM}};
  regs_31 = _RAND_31[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Csrs(
  input         clock,
  input         reset,
  input  [11:0] io_rs_id, // @[playground/src/noop/regs.scala 27:16]
  output [63:0] io_rs_data, // @[playground/src/noop/regs.scala 27:16]
  output        io_rs_is_err, // @[playground/src/noop/regs.scala 27:16]
  input  [11:0] io_rd_id, // @[playground/src/noop/regs.scala 27:16]
  input  [63:0] io_rd_data, // @[playground/src/noop/regs.scala 27:16]
  input         io_rd_en, // @[playground/src/noop/regs.scala 27:16]
  input  [63:0] io_excep_cause, // @[playground/src/noop/regs.scala 27:16]
  input  [63:0] io_excep_tval, // @[playground/src/noop/regs.scala 27:16]
  input         io_excep_en, // @[playground/src/noop/regs.scala 27:16]
  input  [63:0] io_excep_pc, // @[playground/src/noop/regs.scala 27:16]
  input  [1:0]  io_excep_etype, // @[playground/src/noop/regs.scala 27:16]
  output [1:0]  io_mmuState_priv, // @[playground/src/noop/regs.scala 27:16]
  output [63:0] io_mmuState_mstatus, // @[playground/src/noop/regs.scala 27:16]
  output [63:0] io_mmuState_satp, // @[playground/src/noop/regs.scala 27:16]
  output [1:0]  io_idState_priv, // @[playground/src/noop/regs.scala 27:16]
  output [63:0] io_reg2if_seq_pc, // @[playground/src/noop/regs.scala 27:16]
  output        io_reg2if_valid, // @[playground/src/noop/regs.scala 27:16]
  output        io_intr_out_en, // @[playground/src/noop/regs.scala 27:16]
  output [63:0] io_intr_out_cause, // @[playground/src/noop/regs.scala 27:16]
  input         io_clint_raise, // @[playground/src/noop/regs.scala 27:16]
  input         io_clint_clear, // @[playground/src/noop/regs.scala 27:16]
  input         io_plic_m_raise, // @[playground/src/noop/regs.scala 27:16]
  input         io_plic_m_clear, // @[playground/src/noop/regs.scala 27:16]
  input         io_plic_s_raise, // @[playground/src/noop/regs.scala 27:16]
  input         io_plic_s_clear, // @[playground/src/noop/regs.scala 27:16]
  output [63:0] io_updateNextPc_seq_pc, // @[playground/src/noop/regs.scala 27:16]
  output        io_updateNextPc_valid, // @[playground/src/noop/regs.scala 27:16]
  input         io_intr_msip_raise, // @[playground/src/noop/regs.scala 27:16]
  input         io_intr_msip_clear // @[playground/src/noop/regs.scala 27:16]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [63:0] _RAND_14;
  reg [63:0] _RAND_15;
  reg [63:0] _RAND_16;
  reg [63:0] _RAND_17;
  reg [63:0] _RAND_18;
  reg [63:0] _RAND_19;
  reg [63:0] _RAND_20;
  reg [63:0] _RAND_21;
  reg [63:0] _RAND_22;
  reg [63:0] _RAND_23;
  reg [63:0] _RAND_24;
  reg [63:0] _RAND_25;
  reg [63:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [63:0] _RAND_29;
  reg [31:0] _RAND_30;
`endif // RANDOMIZE_REG_INIT
  wire [1:0] updateCsrs_priv; // @[playground/src/noop/regs.scala 298:28]
  wire [75:0] updateCsrs_mstatus; // @[playground/src/noop/regs.scala 298:28]
  wire [75:0] updateCsrs_mepc; // @[playground/src/noop/regs.scala 298:28]
  wire [75:0] updateCsrs_mtval; // @[playground/src/noop/regs.scala 298:28]
  wire [75:0] updateCsrs_mscratch; // @[playground/src/noop/regs.scala 298:28]
  wire [75:0] updateCsrs_mcause; // @[playground/src/noop/regs.scala 298:28]
  wire [75:0] updateCsrs_mtvec; // @[playground/src/noop/regs.scala 298:28]
  wire [75:0] updateCsrs_mie; // @[playground/src/noop/regs.scala 298:28]
  wire [75:0] updateCsrs_mip; // @[playground/src/noop/regs.scala 298:28]
  wire [75:0] updateCsrs_medeleg; // @[playground/src/noop/regs.scala 298:28]
  wire [75:0] updateCsrs_mideleg; // @[playground/src/noop/regs.scala 298:28]
  wire [75:0] updateCsrs_sepc; // @[playground/src/noop/regs.scala 298:28]
  wire [75:0] updateCsrs_stval; // @[playground/src/noop/regs.scala 298:28]
  wire [75:0] updateCsrs_sscratch; // @[playground/src/noop/regs.scala 298:28]
  wire [75:0] updateCsrs_stvec; // @[playground/src/noop/regs.scala 298:28]
  wire [75:0] updateCsrs_satp; // @[playground/src/noop/regs.scala 298:28]
  wire [75:0] updateCsrs_scause; // @[playground/src/noop/regs.scala 298:28]
  wire  updateCsrs_clock; // @[playground/src/noop/regs.scala 298:28]
  reg [1:0] priv; // @[playground/src/noop/regs.scala 41:30]
  reg [63:0] misa; // @[playground/src/noop/regs.scala 42:30]
  reg [63:0] mstatus; // @[playground/src/noop/regs.scala 43:30]
  reg [63:0] mepc; // @[playground/src/noop/regs.scala 44:30]
  reg [63:0] mtval; // @[playground/src/noop/regs.scala 45:30]
  reg [63:0] mscratch; // @[playground/src/noop/regs.scala 46:30]
  reg [63:0] mcause; // @[playground/src/noop/regs.scala 47:30]
  reg [63:0] mtvec; // @[playground/src/noop/regs.scala 48:30]
  reg [63:0] mie; // @[playground/src/noop/regs.scala 49:30]
  reg [63:0] mip; // @[playground/src/noop/regs.scala 50:30]
  reg [63:0] medeleg; // @[playground/src/noop/regs.scala 51:30]
  reg [63:0] mideleg; // @[playground/src/noop/regs.scala 52:30]
  reg [31:0] mcounteren; // @[playground/src/noop/regs.scala 53:30]
  reg [31:0] scounteren; // @[playground/src/noop/regs.scala 54:30]
  reg [63:0] sepc; // @[playground/src/noop/regs.scala 55:30]
  reg [63:0] stval; // @[playground/src/noop/regs.scala 56:30]
  reg [63:0] sscratch; // @[playground/src/noop/regs.scala 57:30]
  reg [63:0] stvec; // @[playground/src/noop/regs.scala 58:30]
  reg [63:0] satp; // @[playground/src/noop/regs.scala 59:30]
  reg [63:0] scause; // @[playground/src/noop/regs.scala 60:30]
  reg [63:0] pmpaddr0; // @[playground/src/noop/regs.scala 61:30]
  reg [63:0] pmpaddr1; // @[playground/src/noop/regs.scala 62:30]
  reg [63:0] pmpaddr2; // @[playground/src/noop/regs.scala 63:30]
  reg [63:0] pmpaddr3; // @[playground/src/noop/regs.scala 64:30]
  reg [63:0] uscratch; // @[playground/src/noop/regs.scala 65:30]
  reg [63:0] mhartid; // @[playground/src/noop/regs.scala 67:30]
  wire [63:0] sstatus = mstatus & 64'h80000003000de122; // @[playground/src/noop/regs.scala 68:31]
  reg [63:0] forceJmp_seq_pc; // @[playground/src/noop/regs.scala 74:34]
  reg  forceJmp_valid; // @[playground/src/noop/regs.scala 74:34]
  wire [1:0] _priv_T_1 = {1'h0,sstatus[8]}; // @[playground/src/noop/regs.scala 84:35]
  wire [63:0] new_sstatus = {sstatus[63:9],1'h0,sstatus[7:6],1'h1,sstatus[4:2],sstatus[5],sstatus[0]}; // @[playground/src/noop/regs.scala 85:34]
  wire [63:0] _mstatus_T_1 = mstatus & 64'hfffffffffff21edd; // @[playground/src/noop/common.scala 201:17]
  wire [63:0] _mstatus_T_2 = new_sstatus & 64'hde122; // @[playground/src/noop/common.scala 201:36]
  wire [63:0] _mstatus_T_3 = _mstatus_T_1 | _mstatus_T_2; // @[playground/src/noop/common.scala 201:26]
  wire [63:0] new_mstatus = {mstatus[63:13],2'h0,mstatus[10:8],1'h1,mstatus[6:4],mstatus[7],mstatus[2:0]}; // @[playground/src/noop/regs.scala 92:34]
  wire [63:0] deleg = io_excep_cause[63] ? mideleg : medeleg; // @[playground/src/noop/regs.scala 96:28]
  wire  _T_2 = priv <= 2'h1; // @[playground/src/noop/regs.scala 97:23]
  wire [63:0] _T_4 = deleg >> io_excep_cause[62:0]; // @[playground/src/noop/regs.scala 97:40]
  wire [65:0] _GEN_109 = {io_excep_cause, 2'h0}; // @[playground/src/noop/regs.scala 98:66]
  wire [66:0] _seq_pc_T_2 = {{1'd0}, _GEN_109}; // @[playground/src/noop/regs.scala 98:66]
  wire [66:0] _seq_pc_T_3 = stvec[1] ? _seq_pc_T_2 : 67'h0; // @[playground/src/noop/regs.scala 98:41]
  wire [66:0] _GEN_113 = {{3'd0}, stvec}; // @[playground/src/noop/regs.scala 98:36]
  wire [66:0] seq_pc = _GEN_113 + _seq_pc_T_3; // @[playground/src/noop/regs.scala 98:36]
  wire [63:0] new_sstatus_1 = {sstatus[63:9],priv[0],sstatus[7:6],sstatus[1],sstatus[4:2],1'h0,sstatus[0]}; // @[playground/src/noop/regs.scala 104:38]
  wire [63:0] _mstatus_T_6 = new_sstatus_1 & 64'hde122; // @[playground/src/noop/common.scala 201:36]
  wire [63:0] _mstatus_T_7 = _mstatus_T_1 | _mstatus_T_6; // @[playground/src/noop/common.scala 201:26]
  wire [66:0] _seq_pc_T_7 = mtvec[1] ? _seq_pc_T_2 : 67'h0; // @[playground/src/noop/regs.scala 109:46]
  wire [66:0] _GEN_124 = {{3'd0}, mtvec}; // @[playground/src/noop/regs.scala 109:41]
  wire [66:0] seq_pc_1 = _GEN_124 + _seq_pc_T_7; // @[playground/src/noop/regs.scala 109:41]
  wire [63:0] new_mstatus_1 = {mstatus[63:13],priv,mstatus[10:8],mstatus[3],mstatus[6:4],1'h0,mstatus[2:0]}; // @[playground/src/noop/regs.scala 115:38]
  wire [66:0] _GEN_0 = priv <= 2'h1 & _T_4[0] ? seq_pc : seq_pc_1; // @[playground/src/noop/regs.scala 110:33 97:54 99:33]
  wire [63:0] _GEN_2 = priv <= 2'h1 & _T_4[0] ? io_excep_cause : scause; // @[playground/src/noop/regs.scala 101:33 60:30 97:54]
  wire [63:0] _GEN_3 = priv <= 2'h1 & _T_4[0] ? io_excep_pc : sepc; // @[playground/src/noop/regs.scala 102:33 55:30 97:54]
  wire [63:0] _GEN_4 = priv <= 2'h1 & _T_4[0] ? _mstatus_T_7 : new_mstatus_1; // @[playground/src/noop/regs.scala 105:33 116:33 97:54]
  wire [63:0] _GEN_5 = priv <= 2'h1 & _T_4[0] ? io_excep_tval : stval; // @[playground/src/noop/regs.scala 106:33 56:30 97:54]
  wire [1:0] _GEN_6 = priv <= 2'h1 & _T_4[0] ? 2'h1 : 2'h3; // @[playground/src/noop/regs.scala 107:33 118:33 97:54]
  wire [63:0] _GEN_7 = priv <= 2'h1 & _T_4[0] ? mcause : io_excep_cause; // @[playground/src/noop/regs.scala 47:30 112:33 97:54]
  wire [63:0] _GEN_8 = priv <= 2'h1 & _T_4[0] ? mepc : io_excep_pc; // @[playground/src/noop/regs.scala 44:30 113:33 97:54]
  wire [63:0] _GEN_9 = priv <= 2'h1 & _T_4[0] ? mtval : io_excep_tval; // @[playground/src/noop/regs.scala 45:30 117:33 97:54]
  wire [66:0] _GEN_10 = io_excep_etype == 2'h3 ? {{3'd0}, mepc} : _GEN_0; // @[playground/src/noop/regs.scala 87:50 88:29]
  wire [63:0] _GEN_13 = io_excep_etype == 2'h3 ? new_mstatus : _GEN_4; // @[playground/src/noop/regs.scala 87:50 93:29]
  wire [63:0] _GEN_14 = io_excep_etype == 2'h3 ? scause : _GEN_2; // @[playground/src/noop/regs.scala 60:30 87:50]
  wire [63:0] _GEN_15 = io_excep_etype == 2'h3 ? sepc : _GEN_3; // @[playground/src/noop/regs.scala 55:30 87:50]
  wire [63:0] _GEN_16 = io_excep_etype == 2'h3 ? stval : _GEN_5; // @[playground/src/noop/regs.scala 56:30 87:50]
  wire [63:0] _GEN_17 = io_excep_etype == 2'h3 ? mcause : _GEN_7; // @[playground/src/noop/regs.scala 47:30 87:50]
  wire [63:0] _GEN_18 = io_excep_etype == 2'h3 ? mepc : _GEN_8; // @[playground/src/noop/regs.scala 44:30 87:50]
  wire [63:0] _GEN_19 = io_excep_etype == 2'h3 ? mtval : _GEN_9; // @[playground/src/noop/regs.scala 45:30 87:50]
  wire [66:0] _GEN_20 = io_excep_etype == 2'h2 ? {{3'd0}, sepc} : _GEN_10; // @[playground/src/noop/regs.scala 80:44 81:29]
  wire [63:0] _GEN_23 = io_excep_etype == 2'h2 ? _mstatus_T_3 : _GEN_13; // @[playground/src/noop/regs.scala 80:44 86:29]
  wire [63:0] _GEN_24 = io_excep_etype == 2'h2 ? scause : _GEN_14; // @[playground/src/noop/regs.scala 60:30 80:44]
  wire [63:0] _GEN_25 = io_excep_etype == 2'h2 ? sepc : _GEN_15; // @[playground/src/noop/regs.scala 55:30 80:44]
  wire [63:0] _GEN_26 = io_excep_etype == 2'h2 ? stval : _GEN_16; // @[playground/src/noop/regs.scala 56:30 80:44]
  wire [63:0] _GEN_27 = io_excep_etype == 2'h2 ? mcause : _GEN_17; // @[playground/src/noop/regs.scala 47:30 80:44]
  wire [63:0] _GEN_28 = io_excep_etype == 2'h2 ? mepc : _GEN_18; // @[playground/src/noop/regs.scala 44:30 80:44]
  wire [63:0] _GEN_29 = io_excep_etype == 2'h2 ? mtval : _GEN_19; // @[playground/src/noop/regs.scala 45:30 80:44]
  wire [66:0] _GEN_30 = io_excep_en ? _GEN_20 : {{3'd0}, forceJmp_seq_pc}; // @[playground/src/noop/regs.scala 79:22 74:34]
  wire [63:0] _GEN_33 = io_excep_en ? _GEN_23 : mstatus; // @[playground/src/noop/regs.scala 79:22 43:30]
  wire [63:0] _GEN_34 = io_excep_en ? _GEN_24 : scause; // @[playground/src/noop/regs.scala 79:22 60:30]
  wire [63:0] _GEN_35 = io_excep_en ? _GEN_25 : sepc; // @[playground/src/noop/regs.scala 79:22 55:30]
  wire [63:0] _GEN_36 = io_excep_en ? _GEN_26 : stval; // @[playground/src/noop/regs.scala 79:22 56:30]
  wire [63:0] _GEN_37 = io_excep_en ? _GEN_27 : mcause; // @[playground/src/noop/regs.scala 79:22 47:30]
  wire [63:0] _GEN_38 = io_excep_en ? _GEN_28 : mepc; // @[playground/src/noop/regs.scala 79:22 44:30]
  wire [63:0] _GEN_39 = io_excep_en ? _GEN_29 : mtval; // @[playground/src/noop/regs.scala 79:22 45:30]
  reg  intr_out_r_en; // @[playground/src/noop/regs.scala 123:29]
  reg [63:0] intr_out_r_cause; // @[playground/src/noop/regs.scala 123:29]
  reg  intr_seip; // @[playground/src/noop/regs.scala 125:28]
  wire [63:0] _mip_T_2 = mip & 64'hffffffffffffff7f; // @[playground/src/noop/common.scala 201:17]
  wire [63:0] _mip_T_4 = _mip_T_2 | 64'h80; // @[playground/src/noop/common.scala 201:26]
  wire [63:0] _GEN_40 = io_clint_raise ? _mip_T_4 : mip; // @[playground/src/noop/regs.scala 126:25 127:13 50:30]
  wire [63:0] _GEN_41 = io_clint_clear ? _mip_T_2 : _GEN_40; // @[playground/src/noop/regs.scala 129:25 130:13]
  wire [63:0] _mip_T_11 = mip & 64'hfffffffffffff7ff; // @[playground/src/noop/common.scala 201:17]
  wire [63:0] _mip_T_13 = _mip_T_11 | 64'h800; // @[playground/src/noop/common.scala 201:26]
  wire [63:0] _GEN_42 = io_plic_m_raise ? _mip_T_13 : _GEN_41; // @[playground/src/noop/regs.scala 132:26 133:13]
  wire [63:0] _GEN_43 = io_plic_m_clear ? _mip_T_11 : _GEN_42; // @[playground/src/noop/regs.scala 135:26 136:13]
  wire  _GEN_44 = io_plic_s_raise | intr_seip; // @[playground/src/noop/regs.scala 138:26 139:19 125:28]
  wire [63:0] _mip_T_20 = mip & 64'hfffffffffffffff7; // @[playground/src/noop/common.scala 201:17]
  wire [63:0] _mip_T_22 = _mip_T_20 | 64'h8; // @[playground/src/noop/common.scala 201:26]
  wire [63:0] _GEN_46 = io_intr_msip_raise ? _mip_T_22 : _GEN_43; // @[playground/src/noop/regs.scala 144:29 145:13]
  wire [63:0] _GEN_47 = io_intr_msip_clear ? _mip_T_20 : _GEN_46; // @[playground/src/noop/regs.scala 147:29 148:13]
  wire [9:0] _GEN_131 = {intr_seip, 9'h0}; // @[playground/src/noop/regs.scala 150:42]
  wire [15:0] _pending_int_T = {{6'd0}, _GEN_131}; // @[playground/src/noop/regs.scala 150:42]
  wire [63:0] _GEN_139 = {{48'd0}, _pending_int_T}; // @[playground/src/noop/regs.scala 150:29]
  wire [63:0] _pending_int_T_1 = mip | _GEN_139; // @[playground/src/noop/regs.scala 150:29]
  wire [63:0] pending_int = _pending_int_T_1 & mie; // @[playground/src/noop/regs.scala 150:59]
  wire  m_enable = priv < 2'h3 | priv == 2'h3 & mstatus[3]; // @[playground/src/noop/regs.scala 151:35]
  wire [63:0] _enable_int_m_T = ~mideleg; // @[playground/src/noop/regs.scala 152:38]
  wire [63:0] _enable_int_m_T_1 = pending_int & _enable_int_m_T; // @[playground/src/noop/regs.scala 152:36]
  wire [63:0] _enable_int_m_T_4 = m_enable ? 64'hffffffffffffffff : 64'h0; // @[playground/src/noop/regs.scala 152:53]
  wire [63:0] enable_int_m = _enable_int_m_T_1 & _enable_int_m_T_4; // @[playground/src/noop/regs.scala 152:47]
  wire  s_enable = _T_2 & mstatus[1]; // @[playground/src/noop/regs.scala 153:36]
  wire [63:0] _enable_int_s_T = pending_int & mideleg; // @[playground/src/noop/regs.scala 154:36]
  wire [63:0] _enable_int_s_T_3 = s_enable ? 64'hffffffffffffffff : 64'h0; // @[playground/src/noop/regs.scala 154:52]
  wire [63:0] enable_int_s = _enable_int_s_T & _enable_int_s_T_3; // @[playground/src/noop/regs.scala 154:46]
  wire [63:0] enable_int = enable_int_m != 64'h0 ? enable_int_m : enable_int_s; // @[playground/src/noop/regs.scala 155:25]
  wire [5:0] _intr_out_r_cause_T_6 = enable_int[5] ? 6'h5 : 6'h3f; // @[src/main/scala/chisel3/util/Mux.scala 47:70]
  wire [5:0] _intr_out_r_cause_T_7 = enable_int[1] ? 6'h1 : _intr_out_r_cause_T_6; // @[src/main/scala/chisel3/util/Mux.scala 47:70]
  wire [5:0] _intr_out_r_cause_T_8 = enable_int[9] ? 6'h9 : _intr_out_r_cause_T_7; // @[src/main/scala/chisel3/util/Mux.scala 47:70]
  wire [5:0] _intr_out_r_cause_T_9 = enable_int[7] ? 6'h7 : _intr_out_r_cause_T_8; // @[src/main/scala/chisel3/util/Mux.scala 47:70]
  wire [5:0] _intr_out_r_cause_T_10 = enable_int[3] ? 6'h3 : _intr_out_r_cause_T_9; // @[src/main/scala/chisel3/util/Mux.scala 47:70]
  wire [5:0] _intr_out_r_cause_T_11 = enable_int[11] ? 6'hb : _intr_out_r_cause_T_10; // @[src/main/scala/chisel3/util/Mux.scala 47:70]
  wire [63:0] _GEN_148 = {{58'd0}, _intr_out_r_cause_T_11}; // @[playground/src/noop/regs.scala 167:8]
  wire [63:0] _intr_out_r_cause_T_13 = _GEN_148 | 64'h8000000000000000; // @[playground/src/noop/regs.scala 167:8]
  wire [63:0] _io_rs_data_T = mie & mideleg; // @[playground/src/noop/regs.scala 211:27]
  wire [63:0] _io_rs_data_T_1 = mip & 64'h222; // @[playground/src/noop/regs.scala 213:27]
  wire [63:0] _GEN_48 = io_rs_id == 12'hf14 ? mhartid : 64'h0; // @[playground/src/noop/regs.scala 226:41 227:20 229:25]
  wire  _GEN_49 = io_rs_id == 12'hf14 ? 1'h0 : 1'h1; // @[playground/src/noop/regs.scala 169:21 226:41 230:25]
  wire [63:0] _GEN_50 = io_rs_id == 12'h40 ? uscratch : _GEN_48; // @[playground/src/noop/regs.scala 224:42 225:20]
  wire  _GEN_51 = io_rs_id == 12'h40 ? 1'h0 : _GEN_49; // @[playground/src/noop/regs.scala 169:21 224:42]
  wire [63:0] _GEN_52 = io_rs_id == 12'h3a0 ? pmpaddr3 : _GEN_50; // @[playground/src/noop/regs.scala 222:41 223:20]
  wire  _GEN_53 = io_rs_id == 12'h3a0 ? 1'h0 : _GEN_51; // @[playground/src/noop/regs.scala 169:21 222:41]
  wire [63:0] _GEN_54 = io_rs_id == 12'h3b3 ? pmpaddr3 : _GEN_52; // @[playground/src/noop/regs.scala 220:42 221:20]
  wire  _GEN_55 = io_rs_id == 12'h3b3 ? 1'h0 : _GEN_53; // @[playground/src/noop/regs.scala 169:21 220:42]
  wire [63:0] _GEN_56 = io_rs_id == 12'h3b2 ? pmpaddr2 : _GEN_54; // @[playground/src/noop/regs.scala 218:42 219:20]
  wire  _GEN_57 = io_rs_id == 12'h3b2 ? 1'h0 : _GEN_55; // @[playground/src/noop/regs.scala 169:21 218:42]
  wire [63:0] _GEN_58 = io_rs_id == 12'h3b1 ? pmpaddr1 : _GEN_56; // @[playground/src/noop/regs.scala 216:42 217:20]
  wire  _GEN_59 = io_rs_id == 12'h3b1 ? 1'h0 : _GEN_57; // @[playground/src/noop/regs.scala 169:21 216:42]
  wire [63:0] _GEN_60 = io_rs_id == 12'h3b0 ? pmpaddr0 : _GEN_58; // @[playground/src/noop/regs.scala 214:42 215:20]
  wire  _GEN_61 = io_rs_id == 12'h3b0 ? 1'h0 : _GEN_59; // @[playground/src/noop/regs.scala 169:21 214:42]
  wire [63:0] _GEN_62 = io_rs_id == 12'h144 ? _io_rs_data_T_1 : _GEN_60; // @[playground/src/noop/regs.scala 212:37 213:20]
  wire  _GEN_63 = io_rs_id == 12'h144 ? 1'h0 : _GEN_61; // @[playground/src/noop/regs.scala 169:21 212:37]
  wire [63:0] _GEN_64 = io_rs_id == 12'h104 ? _io_rs_data_T : _GEN_62; // @[playground/src/noop/regs.scala 210:37 211:20]
  wire  _GEN_65 = io_rs_id == 12'h104 ? 1'h0 : _GEN_63; // @[playground/src/noop/regs.scala 169:21 210:37]
  wire [63:0] _GEN_66 = io_rs_id == 12'h100 ? sstatus : _GEN_64; // @[playground/src/noop/regs.scala 208:41 209:20]
  wire  _GEN_67 = io_rs_id == 12'h100 ? 1'h0 : _GEN_65; // @[playground/src/noop/regs.scala 169:21 208:41]
  wire [63:0] _GEN_68 = io_rs_id == 12'h142 ? scause : _GEN_66; // @[playground/src/noop/regs.scala 206:40 207:20]
  wire  _GEN_69 = io_rs_id == 12'h142 ? 1'h0 : _GEN_67; // @[playground/src/noop/regs.scala 169:21 206:40]
  wire [63:0] _GEN_70 = io_rs_id == 12'h180 ? satp : _GEN_68; // @[playground/src/noop/regs.scala 204:38 205:20]
  wire  _GEN_71 = io_rs_id == 12'h180 ? 1'h0 : _GEN_69; // @[playground/src/noop/regs.scala 169:21 204:38]
  wire [63:0] _GEN_72 = io_rs_id == 12'h105 ? stvec : _GEN_70; // @[playground/src/noop/regs.scala 202:39 203:20]
  wire  _GEN_73 = io_rs_id == 12'h105 ? 1'h0 : _GEN_71; // @[playground/src/noop/regs.scala 169:21 202:39]
  wire [63:0] _GEN_74 = io_rs_id == 12'h140 ? sscratch : _GEN_72; // @[playground/src/noop/regs.scala 200:42 201:20]
  wire  _GEN_75 = io_rs_id == 12'h140 ? 1'h0 : _GEN_73; // @[playground/src/noop/regs.scala 169:21 200:42]
  wire [63:0] _GEN_76 = io_rs_id == 12'h143 ? stval : _GEN_74; // @[playground/src/noop/regs.scala 198:39 199:20]
  wire  _GEN_77 = io_rs_id == 12'h143 ? 1'h0 : _GEN_75; // @[playground/src/noop/regs.scala 169:21 198:39]
  wire [63:0] _GEN_78 = io_rs_id == 12'h141 ? sepc : _GEN_76; // @[playground/src/noop/regs.scala 196:38 197:20]
  wire  _GEN_79 = io_rs_id == 12'h141 ? 1'h0 : _GEN_77; // @[playground/src/noop/regs.scala 169:21 196:38]
  wire [63:0] _GEN_80 = io_rs_id == 12'h106 ? {{32'd0}, scounteren} : _GEN_78; // @[playground/src/noop/regs.scala 194:44 195:20]
  wire  _GEN_81 = io_rs_id == 12'h106 ? 1'h0 : _GEN_79; // @[playground/src/noop/regs.scala 169:21 194:44]
  wire [63:0] _GEN_82 = io_rs_id == 12'h306 ? {{32'd0}, mcounteren} : _GEN_80; // @[playground/src/noop/regs.scala 192:44 193:20]
  wire  _GEN_83 = io_rs_id == 12'h306 ? 1'h0 : _GEN_81; // @[playground/src/noop/regs.scala 169:21 192:44]
  wire [63:0] _GEN_84 = io_rs_id == 12'h303 ? mideleg : _GEN_82; // @[playground/src/noop/regs.scala 190:41 191:20]
  wire  _GEN_85 = io_rs_id == 12'h303 ? 1'h0 : _GEN_83; // @[playground/src/noop/regs.scala 169:21 190:41]
  wire [63:0] _GEN_86 = io_rs_id == 12'h302 ? medeleg : _GEN_84; // @[playground/src/noop/regs.scala 188:41 189:20]
  wire  _GEN_87 = io_rs_id == 12'h302 ? 1'h0 : _GEN_85; // @[playground/src/noop/regs.scala 169:21 188:41]
  wire [63:0] _GEN_88 = io_rs_id == 12'h342 ? mcause : _GEN_86; // @[playground/src/noop/regs.scala 186:40 187:20]
  wire  _GEN_89 = io_rs_id == 12'h342 ? 1'h0 : _GEN_87; // @[playground/src/noop/regs.scala 169:21 186:40]
  wire [63:0] _GEN_90 = io_rs_id == 12'h344 ? mip : _GEN_88; // @[playground/src/noop/regs.scala 184:37 185:20]
  wire  _GEN_91 = io_rs_id == 12'h344 ? 1'h0 : _GEN_89; // @[playground/src/noop/regs.scala 169:21 184:37]
  wire [63:0] _GEN_92 = io_rs_id == 12'h304 ? mie : _GEN_90; // @[playground/src/noop/regs.scala 182:37 183:20]
  wire  _GEN_93 = io_rs_id == 12'h304 ? 1'h0 : _GEN_91; // @[playground/src/noop/regs.scala 169:21 182:37]
  wire [63:0] _GEN_94 = io_rs_id == 12'h305 ? mtvec : _GEN_92; // @[playground/src/noop/regs.scala 180:39 181:20]
  wire  _GEN_95 = io_rs_id == 12'h305 ? 1'h0 : _GEN_93; // @[playground/src/noop/regs.scala 169:21 180:39]
  wire [63:0] _GEN_96 = io_rs_id == 12'h340 ? mscratch : _GEN_94; // @[playground/src/noop/regs.scala 178:42 179:20]
  wire  _GEN_97 = io_rs_id == 12'h340 ? 1'h0 : _GEN_95; // @[playground/src/noop/regs.scala 169:21 178:42]
  wire [63:0] _GEN_98 = io_rs_id == 12'h343 ? mtval : _GEN_96; // @[playground/src/noop/regs.scala 176:39 177:20]
  wire  _GEN_99 = io_rs_id == 12'h343 ? 1'h0 : _GEN_97; // @[playground/src/noop/regs.scala 169:21 176:39]
  wire [63:0] _GEN_100 = io_rs_id == 12'h341 ? mepc : _GEN_98; // @[playground/src/noop/regs.scala 174:38 175:20]
  wire  _GEN_101 = io_rs_id == 12'h341 ? 1'h0 : _GEN_99; // @[playground/src/noop/regs.scala 169:21 174:38]
  wire [63:0] _GEN_102 = io_rs_id == 12'h300 ? mstatus : _GEN_100; // @[playground/src/noop/regs.scala 172:41 173:20]
  wire  _GEN_103 = io_rs_id == 12'h300 ? 1'h0 : _GEN_101; // @[playground/src/noop/regs.scala 169:21 172:41]
  wire [63:0] new_mstatus_2 = io_rd_data & 64'h7e7faa; // @[playground/src/noop/regs.scala 236:38]
  wire [63:0] sd = io_rd_data[14:13] == 2'h3 | io_rd_data[16:15] == 2'h3 ? 64'h8000000000000000 : 64'h0; // @[playground/src/noop/regs.scala 237:30]
  wire [63:0] _mstatus_T_9 = new_mstatus_2 | sd; // @[playground/src/noop/regs.scala 238:86]
  wire [63:0] _mstatus_T_11 = mstatus & 64'h7fffffffff818055; // @[playground/src/noop/common.scala 201:17]
  wire [63:0] _mstatus_T_12 = _mstatus_T_9 & 64'h80000000007e7faa; // @[playground/src/noop/common.scala 201:36]
  wire [63:0] _mstatus_T_13 = _mstatus_T_11 | _mstatus_T_12; // @[playground/src/noop/common.scala 201:26]
  wire [63:0] _mip_T_28 = mip & 64'hffffffffffffffdd; // @[playground/src/noop/common.scala 201:17]
  wire [63:0] _mip_T_29 = io_rd_data & 64'h22; // @[playground/src/noop/common.scala 201:36]
  wire [63:0] _mip_T_30 = _mip_T_28 | _mip_T_29; // @[playground/src/noop/common.scala 201:26]
  wire [63:0] _mip_T_32 = _mip_T_30 | _GEN_139; // @[playground/src/noop/regs.scala 250:61]
  wire [63:0] _medeleg_T = io_rd_data & 64'hb309; // @[playground/src/noop/regs.scala 254:31]
  wire [63:0] _mideleg_T = io_rd_data & 64'h222; // @[playground/src/noop/regs.scala 256:31]
  wire [63:0] _satp_T_1 = satp & 64'hffff00000000000; // @[playground/src/noop/common.scala 201:17]
  wire [63:0] _satp_T_2 = io_rd_data & 64'hf0000fffffffffff; // @[playground/src/noop/common.scala 201:36]
  wire [63:0] _satp_T_3 = _satp_T_1 | _satp_T_2; // @[playground/src/noop/common.scala 201:26]
  wire [63:0] _new_mstatus_T_13 = io_rd_data & 64'hde122; // @[playground/src/noop/common.scala 201:36]
  wire [63:0] new_mstatus_3 = _mstatus_T_1 | _new_mstatus_T_13; // @[playground/src/noop/common.scala 201:26]
  wire [63:0] _mstatus_T_16 = {sd[63:62],new_mstatus_3[61:0]}; // @[playground/src/noop/regs.scala 276:23]
  wire [63:0] _mie_T_1 = mie & _enable_int_m_T; // @[playground/src/noop/common.scala 201:17]
  wire [63:0] _mie_T_2 = io_rd_data & mideleg; // @[playground/src/noop/common.scala 201:36]
  wire [63:0] _mie_T_3 = _mie_T_1 | _mie_T_2; // @[playground/src/noop/common.scala 201:26]
  wire [63:0] _mip_T_34 = mip & 64'hfffffffffffffddd; // @[playground/src/noop/common.scala 201:17]
  wire [63:0] _mip_T_36 = _mip_T_34 | _mideleg_T; // @[playground/src/noop/common.scala 201:26]
  wire [63:0] _pmpaddr0_T = io_rd_data & 64'h3fffffffffffff; // @[playground/src/noop/regs.scala 282:32]
  wire [63:0] _GEN_106 = io_rd_id == 12'hf14 ? io_rd_data : mhartid; // @[playground/src/noop/regs.scala 293:41 294:17 67:30]
  wire [63:0] _GEN_107 = io_rd_id == 12'h40 ? io_rd_data : uscratch; // @[playground/src/noop/regs.scala 291:42 292:18 65:30]
  wire [63:0] _GEN_108 = io_rd_id == 12'h40 ? mhartid : _GEN_106; // @[playground/src/noop/regs.scala 291:42 67:30]
  wire [63:0] _GEN_110 = io_rd_id == 12'h3a0 ? uscratch : _GEN_107; // @[playground/src/noop/regs.scala 289:41 65:30]
  wire [63:0] _GEN_111 = io_rd_id == 12'h3a0 ? mhartid : _GEN_108; // @[playground/src/noop/regs.scala 289:41 67:30]
  wire [63:0] _GEN_112 = io_rd_id == 12'h3b3 ? _pmpaddr0_T : pmpaddr3; // @[playground/src/noop/regs.scala 287:42 288:18 64:30]
  wire [63:0] _GEN_114 = io_rd_id == 12'h3b3 ? uscratch : _GEN_110; // @[playground/src/noop/regs.scala 287:42 65:30]
  wire [63:0] _GEN_115 = io_rd_id == 12'h3b3 ? mhartid : _GEN_111; // @[playground/src/noop/regs.scala 287:42 67:30]
  wire [63:0] _GEN_116 = io_rd_id == 12'h3b2 ? _pmpaddr0_T : pmpaddr2; // @[playground/src/noop/regs.scala 285:42 286:18 63:30]
  wire [63:0] _GEN_117 = io_rd_id == 12'h3b2 ? pmpaddr3 : _GEN_112; // @[playground/src/noop/regs.scala 285:42 64:30]
  wire [63:0] _GEN_119 = io_rd_id == 12'h3b2 ? uscratch : _GEN_114; // @[playground/src/noop/regs.scala 285:42 65:30]
  wire [63:0] _GEN_120 = io_rd_id == 12'h3b2 ? mhartid : _GEN_115; // @[playground/src/noop/regs.scala 285:42 67:30]
  wire [63:0] _GEN_121 = io_rd_id == 12'h3b1 ? _pmpaddr0_T : pmpaddr1; // @[playground/src/noop/regs.scala 283:42 284:18 62:30]
  wire [63:0] _GEN_122 = io_rd_id == 12'h3b1 ? pmpaddr2 : _GEN_116; // @[playground/src/noop/regs.scala 283:42 63:30]
  wire [63:0] _GEN_123 = io_rd_id == 12'h3b1 ? pmpaddr3 : _GEN_117; // @[playground/src/noop/regs.scala 283:42 64:30]
  wire [63:0] _GEN_125 = io_rd_id == 12'h3b1 ? uscratch : _GEN_119; // @[playground/src/noop/regs.scala 283:42 65:30]
  wire [63:0] _GEN_126 = io_rd_id == 12'h3b1 ? mhartid : _GEN_120; // @[playground/src/noop/regs.scala 283:42 67:30]
  wire [63:0] _GEN_127 = io_rd_id == 12'h3b0 ? _pmpaddr0_T : pmpaddr0; // @[playground/src/noop/regs.scala 281:42 282:18 61:30]
  wire [63:0] _GEN_128 = io_rd_id == 12'h3b0 ? pmpaddr1 : _GEN_121; // @[playground/src/noop/regs.scala 281:42 62:30]
  wire [63:0] _GEN_129 = io_rd_id == 12'h3b0 ? pmpaddr2 : _GEN_122; // @[playground/src/noop/regs.scala 281:42 63:30]
  wire [63:0] _GEN_130 = io_rd_id == 12'h3b0 ? pmpaddr3 : _GEN_123; // @[playground/src/noop/regs.scala 281:42 64:30]
  wire [63:0] _GEN_132 = io_rd_id == 12'h3b0 ? uscratch : _GEN_125; // @[playground/src/noop/regs.scala 281:42 65:30]
  wire [63:0] _GEN_133 = io_rd_id == 12'h3b0 ? mhartid : _GEN_126; // @[playground/src/noop/regs.scala 281:42 67:30]
  wire [63:0] _GEN_134 = io_rd_id == 12'h144 ? _mip_T_36 : _GEN_47; // @[playground/src/noop/regs.scala 279:37 280:13]
  wire [63:0] _GEN_135 = io_rd_id == 12'h144 ? pmpaddr0 : _GEN_127; // @[playground/src/noop/regs.scala 279:37 61:30]
  wire [63:0] _GEN_136 = io_rd_id == 12'h144 ? pmpaddr1 : _GEN_128; // @[playground/src/noop/regs.scala 279:37 62:30]
  wire [63:0] _GEN_137 = io_rd_id == 12'h144 ? pmpaddr2 : _GEN_129; // @[playground/src/noop/regs.scala 279:37 63:30]
  wire [63:0] _GEN_138 = io_rd_id == 12'h144 ? pmpaddr3 : _GEN_130; // @[playground/src/noop/regs.scala 279:37 64:30]
  wire [63:0] _GEN_140 = io_rd_id == 12'h144 ? uscratch : _GEN_132; // @[playground/src/noop/regs.scala 279:37 65:30]
  wire [63:0] _GEN_141 = io_rd_id == 12'h144 ? mhartid : _GEN_133; // @[playground/src/noop/regs.scala 279:37 67:30]
  wire [63:0] _GEN_142 = io_rd_id == 12'h104 ? _mie_T_3 : mie; // @[playground/src/noop/regs.scala 277:37 278:13 49:30]
  wire [63:0] _GEN_143 = io_rd_id == 12'h104 ? _GEN_47 : _GEN_134; // @[playground/src/noop/regs.scala 277:37]
  wire [63:0] _GEN_144 = io_rd_id == 12'h104 ? pmpaddr0 : _GEN_135; // @[playground/src/noop/regs.scala 277:37 61:30]
  wire [63:0] _GEN_145 = io_rd_id == 12'h104 ? pmpaddr1 : _GEN_136; // @[playground/src/noop/regs.scala 277:37 62:30]
  wire [63:0] _GEN_146 = io_rd_id == 12'h104 ? pmpaddr2 : _GEN_137; // @[playground/src/noop/regs.scala 277:37 63:30]
  wire [63:0] _GEN_147 = io_rd_id == 12'h104 ? pmpaddr3 : _GEN_138; // @[playground/src/noop/regs.scala 277:37 64:30]
  wire [63:0] _GEN_149 = io_rd_id == 12'h104 ? uscratch : _GEN_140; // @[playground/src/noop/regs.scala 277:37 65:30]
  wire [63:0] _GEN_150 = io_rd_id == 12'h104 ? mhartid : _GEN_141; // @[playground/src/noop/regs.scala 277:37 67:30]
  wire [63:0] _GEN_151 = io_rd_id == 12'h100 ? _mstatus_T_16 : _GEN_33; // @[playground/src/noop/regs.scala 273:41 276:17]
  wire [63:0] _GEN_152 = io_rd_id == 12'h100 ? mie : _GEN_142; // @[playground/src/noop/regs.scala 273:41 49:30]
  wire [63:0] _GEN_153 = io_rd_id == 12'h100 ? _GEN_47 : _GEN_143; // @[playground/src/noop/regs.scala 273:41]
  wire [63:0] _GEN_154 = io_rd_id == 12'h100 ? pmpaddr0 : _GEN_144; // @[playground/src/noop/regs.scala 273:41 61:30]
  wire [63:0] _GEN_155 = io_rd_id == 12'h100 ? pmpaddr1 : _GEN_145; // @[playground/src/noop/regs.scala 273:41 62:30]
  wire [63:0] _GEN_156 = io_rd_id == 12'h100 ? pmpaddr2 : _GEN_146; // @[playground/src/noop/regs.scala 273:41 63:30]
  wire [63:0] _GEN_157 = io_rd_id == 12'h100 ? pmpaddr3 : _GEN_147; // @[playground/src/noop/regs.scala 273:41 64:30]
  wire [63:0] _GEN_159 = io_rd_id == 12'h100 ? uscratch : _GEN_149; // @[playground/src/noop/regs.scala 273:41 65:30]
  wire [63:0] _GEN_160 = io_rd_id == 12'h100 ? mhartid : _GEN_150; // @[playground/src/noop/regs.scala 273:41 67:30]
  wire [63:0] _GEN_161 = io_rd_id == 12'h142 ? io_rd_data : _GEN_34; // @[playground/src/noop/regs.scala 271:40 272:16]
  wire [63:0] _GEN_162 = io_rd_id == 12'h142 ? _GEN_33 : _GEN_151; // @[playground/src/noop/regs.scala 271:40]
  wire [63:0] _GEN_163 = io_rd_id == 12'h142 ? mie : _GEN_152; // @[playground/src/noop/regs.scala 271:40 49:30]
  wire [63:0] _GEN_164 = io_rd_id == 12'h142 ? _GEN_47 : _GEN_153; // @[playground/src/noop/regs.scala 271:40]
  wire [63:0] _GEN_165 = io_rd_id == 12'h142 ? pmpaddr0 : _GEN_154; // @[playground/src/noop/regs.scala 271:40 61:30]
  wire [63:0] _GEN_166 = io_rd_id == 12'h142 ? pmpaddr1 : _GEN_155; // @[playground/src/noop/regs.scala 271:40 62:30]
  wire [63:0] _GEN_167 = io_rd_id == 12'h142 ? pmpaddr2 : _GEN_156; // @[playground/src/noop/regs.scala 271:40 63:30]
  wire [63:0] _GEN_168 = io_rd_id == 12'h142 ? pmpaddr3 : _GEN_157; // @[playground/src/noop/regs.scala 271:40 64:30]
  wire [63:0] _GEN_170 = io_rd_id == 12'h142 ? uscratch : _GEN_159; // @[playground/src/noop/regs.scala 271:40 65:30]
  wire [63:0] _GEN_171 = io_rd_id == 12'h142 ? mhartid : _GEN_160; // @[playground/src/noop/regs.scala 271:40 67:30]
  wire [63:0] _GEN_172 = io_rd_id == 12'h180 ? _satp_T_3 : satp; // @[playground/src/noop/regs.scala 269:38 270:14 59:30]
  wire [63:0] _GEN_173 = io_rd_id == 12'h180 ? _GEN_34 : _GEN_161; // @[playground/src/noop/regs.scala 269:38]
  wire [63:0] _GEN_174 = io_rd_id == 12'h180 ? _GEN_33 : _GEN_162; // @[playground/src/noop/regs.scala 269:38]
  wire [63:0] _GEN_175 = io_rd_id == 12'h180 ? mie : _GEN_163; // @[playground/src/noop/regs.scala 269:38 49:30]
  wire [63:0] _GEN_176 = io_rd_id == 12'h180 ? _GEN_47 : _GEN_164; // @[playground/src/noop/regs.scala 269:38]
  wire [63:0] _GEN_177 = io_rd_id == 12'h180 ? pmpaddr0 : _GEN_165; // @[playground/src/noop/regs.scala 269:38 61:30]
  wire [63:0] _GEN_178 = io_rd_id == 12'h180 ? pmpaddr1 : _GEN_166; // @[playground/src/noop/regs.scala 269:38 62:30]
  wire [63:0] _GEN_179 = io_rd_id == 12'h180 ? pmpaddr2 : _GEN_167; // @[playground/src/noop/regs.scala 269:38 63:30]
  wire [63:0] _GEN_180 = io_rd_id == 12'h180 ? pmpaddr3 : _GEN_168; // @[playground/src/noop/regs.scala 269:38 64:30]
  wire [63:0] _GEN_182 = io_rd_id == 12'h180 ? uscratch : _GEN_170; // @[playground/src/noop/regs.scala 269:38 65:30]
  wire [63:0] _GEN_183 = io_rd_id == 12'h180 ? mhartid : _GEN_171; // @[playground/src/noop/regs.scala 269:38 67:30]
  wire [63:0] _GEN_184 = io_rd_id == 12'h105 ? io_rd_data : stvec; // @[playground/src/noop/regs.scala 267:39 268:15 58:30]
  wire [63:0] _GEN_185 = io_rd_id == 12'h105 ? satp : _GEN_172; // @[playground/src/noop/regs.scala 267:39 59:30]
  wire [63:0] _GEN_186 = io_rd_id == 12'h105 ? _GEN_34 : _GEN_173; // @[playground/src/noop/regs.scala 267:39]
  wire [63:0] _GEN_187 = io_rd_id == 12'h105 ? _GEN_33 : _GEN_174; // @[playground/src/noop/regs.scala 267:39]
  wire [63:0] _GEN_188 = io_rd_id == 12'h105 ? mie : _GEN_175; // @[playground/src/noop/regs.scala 267:39 49:30]
  wire [63:0] _GEN_189 = io_rd_id == 12'h105 ? _GEN_47 : _GEN_176; // @[playground/src/noop/regs.scala 267:39]
  wire [63:0] _GEN_190 = io_rd_id == 12'h105 ? pmpaddr0 : _GEN_177; // @[playground/src/noop/regs.scala 267:39 61:30]
  wire [63:0] _GEN_191 = io_rd_id == 12'h105 ? pmpaddr1 : _GEN_178; // @[playground/src/noop/regs.scala 267:39 62:30]
  wire [63:0] _GEN_192 = io_rd_id == 12'h105 ? pmpaddr2 : _GEN_179; // @[playground/src/noop/regs.scala 267:39 63:30]
  wire [63:0] _GEN_193 = io_rd_id == 12'h105 ? pmpaddr3 : _GEN_180; // @[playground/src/noop/regs.scala 267:39 64:30]
  wire [63:0] _GEN_195 = io_rd_id == 12'h105 ? uscratch : _GEN_182; // @[playground/src/noop/regs.scala 267:39 65:30]
  wire [63:0] _GEN_196 = io_rd_id == 12'h105 ? mhartid : _GEN_183; // @[playground/src/noop/regs.scala 267:39 67:30]
  wire [63:0] _GEN_197 = io_rd_id == 12'h140 ? io_rd_data : sscratch; // @[playground/src/noop/regs.scala 265:42 266:18 57:30]
  wire [63:0] _GEN_198 = io_rd_id == 12'h140 ? stvec : _GEN_184; // @[playground/src/noop/regs.scala 265:42 58:30]
  wire [63:0] _GEN_199 = io_rd_id == 12'h140 ? satp : _GEN_185; // @[playground/src/noop/regs.scala 265:42 59:30]
  wire [63:0] _GEN_200 = io_rd_id == 12'h140 ? _GEN_34 : _GEN_186; // @[playground/src/noop/regs.scala 265:42]
  wire [63:0] _GEN_201 = io_rd_id == 12'h140 ? _GEN_33 : _GEN_187; // @[playground/src/noop/regs.scala 265:42]
  wire [63:0] _GEN_202 = io_rd_id == 12'h140 ? mie : _GEN_188; // @[playground/src/noop/regs.scala 265:42 49:30]
  wire [63:0] _GEN_203 = io_rd_id == 12'h140 ? _GEN_47 : _GEN_189; // @[playground/src/noop/regs.scala 265:42]
  wire [63:0] _GEN_204 = io_rd_id == 12'h140 ? pmpaddr0 : _GEN_190; // @[playground/src/noop/regs.scala 265:42 61:30]
  wire [63:0] _GEN_205 = io_rd_id == 12'h140 ? pmpaddr1 : _GEN_191; // @[playground/src/noop/regs.scala 265:42 62:30]
  wire [63:0] _GEN_206 = io_rd_id == 12'h140 ? pmpaddr2 : _GEN_192; // @[playground/src/noop/regs.scala 265:42 63:30]
  wire [63:0] _GEN_207 = io_rd_id == 12'h140 ? pmpaddr3 : _GEN_193; // @[playground/src/noop/regs.scala 265:42 64:30]
  wire [63:0] _GEN_209 = io_rd_id == 12'h140 ? uscratch : _GEN_195; // @[playground/src/noop/regs.scala 265:42 65:30]
  wire [63:0] _GEN_210 = io_rd_id == 12'h140 ? mhartid : _GEN_196; // @[playground/src/noop/regs.scala 265:42 67:30]
  wire [63:0] _GEN_211 = io_rd_id == 12'h143 ? io_rd_data : _GEN_36; // @[playground/src/noop/regs.scala 263:39 264:15]
  wire [63:0] _GEN_212 = io_rd_id == 12'h143 ? sscratch : _GEN_197; // @[playground/src/noop/regs.scala 263:39 57:30]
  wire [63:0] _GEN_213 = io_rd_id == 12'h143 ? stvec : _GEN_198; // @[playground/src/noop/regs.scala 263:39 58:30]
  wire [63:0] _GEN_214 = io_rd_id == 12'h143 ? satp : _GEN_199; // @[playground/src/noop/regs.scala 263:39 59:30]
  wire [63:0] _GEN_215 = io_rd_id == 12'h143 ? _GEN_34 : _GEN_200; // @[playground/src/noop/regs.scala 263:39]
  wire [63:0] _GEN_216 = io_rd_id == 12'h143 ? _GEN_33 : _GEN_201; // @[playground/src/noop/regs.scala 263:39]
  wire [63:0] _GEN_217 = io_rd_id == 12'h143 ? mie : _GEN_202; // @[playground/src/noop/regs.scala 263:39 49:30]
  wire [63:0] _GEN_218 = io_rd_id == 12'h143 ? _GEN_47 : _GEN_203; // @[playground/src/noop/regs.scala 263:39]
  wire [63:0] _GEN_219 = io_rd_id == 12'h143 ? pmpaddr0 : _GEN_204; // @[playground/src/noop/regs.scala 263:39 61:30]
  wire [63:0] _GEN_220 = io_rd_id == 12'h143 ? pmpaddr1 : _GEN_205; // @[playground/src/noop/regs.scala 263:39 62:30]
  wire [63:0] _GEN_221 = io_rd_id == 12'h143 ? pmpaddr2 : _GEN_206; // @[playground/src/noop/regs.scala 263:39 63:30]
  wire [63:0] _GEN_222 = io_rd_id == 12'h143 ? pmpaddr3 : _GEN_207; // @[playground/src/noop/regs.scala 263:39 64:30]
  wire [63:0] _GEN_224 = io_rd_id == 12'h143 ? uscratch : _GEN_209; // @[playground/src/noop/regs.scala 263:39 65:30]
  wire [63:0] _GEN_225 = io_rd_id == 12'h143 ? mhartid : _GEN_210; // @[playground/src/noop/regs.scala 263:39 67:30]
  wire [63:0] _GEN_226 = io_rd_id == 12'h141 ? io_rd_data : _GEN_35; // @[playground/src/noop/regs.scala 261:38 262:14]
  wire [63:0] _GEN_227 = io_rd_id == 12'h141 ? _GEN_36 : _GEN_211; // @[playground/src/noop/regs.scala 261:38]
  wire [63:0] _GEN_228 = io_rd_id == 12'h141 ? sscratch : _GEN_212; // @[playground/src/noop/regs.scala 261:38 57:30]
  wire [63:0] _GEN_229 = io_rd_id == 12'h141 ? stvec : _GEN_213; // @[playground/src/noop/regs.scala 261:38 58:30]
  wire [63:0] _GEN_230 = io_rd_id == 12'h141 ? satp : _GEN_214; // @[playground/src/noop/regs.scala 261:38 59:30]
  wire [63:0] _GEN_231 = io_rd_id == 12'h141 ? _GEN_34 : _GEN_215; // @[playground/src/noop/regs.scala 261:38]
  wire [63:0] _GEN_232 = io_rd_id == 12'h141 ? _GEN_33 : _GEN_216; // @[playground/src/noop/regs.scala 261:38]
  wire [63:0] _GEN_233 = io_rd_id == 12'h141 ? mie : _GEN_217; // @[playground/src/noop/regs.scala 261:38 49:30]
  wire [63:0] _GEN_234 = io_rd_id == 12'h141 ? _GEN_47 : _GEN_218; // @[playground/src/noop/regs.scala 261:38]
  wire [63:0] _GEN_235 = io_rd_id == 12'h141 ? pmpaddr0 : _GEN_219; // @[playground/src/noop/regs.scala 261:38 61:30]
  wire [63:0] _GEN_236 = io_rd_id == 12'h141 ? pmpaddr1 : _GEN_220; // @[playground/src/noop/regs.scala 261:38 62:30]
  wire [63:0] _GEN_237 = io_rd_id == 12'h141 ? pmpaddr2 : _GEN_221; // @[playground/src/noop/regs.scala 261:38 63:30]
  wire [63:0] _GEN_238 = io_rd_id == 12'h141 ? pmpaddr3 : _GEN_222; // @[playground/src/noop/regs.scala 261:38 64:30]
  wire [63:0] _GEN_240 = io_rd_id == 12'h141 ? uscratch : _GEN_224; // @[playground/src/noop/regs.scala 261:38 65:30]
  wire [63:0] _GEN_241 = io_rd_id == 12'h141 ? mhartid : _GEN_225; // @[playground/src/noop/regs.scala 261:38 67:30]
  wire [63:0] _GEN_242 = io_rd_id == 12'h106 ? io_rd_data : {{32'd0}, scounteren}; // @[playground/src/noop/regs.scala 259:44 260:20 54:30]
  wire [63:0] _GEN_243 = io_rd_id == 12'h106 ? _GEN_35 : _GEN_226; // @[playground/src/noop/regs.scala 259:44]
  wire [63:0] _GEN_244 = io_rd_id == 12'h106 ? _GEN_36 : _GEN_227; // @[playground/src/noop/regs.scala 259:44]
  wire [63:0] _GEN_245 = io_rd_id == 12'h106 ? sscratch : _GEN_228; // @[playground/src/noop/regs.scala 259:44 57:30]
  wire [63:0] _GEN_246 = io_rd_id == 12'h106 ? stvec : _GEN_229; // @[playground/src/noop/regs.scala 259:44 58:30]
  wire [63:0] _GEN_247 = io_rd_id == 12'h106 ? satp : _GEN_230; // @[playground/src/noop/regs.scala 259:44 59:30]
  wire [63:0] _GEN_248 = io_rd_id == 12'h106 ? _GEN_34 : _GEN_231; // @[playground/src/noop/regs.scala 259:44]
  wire [63:0] _GEN_249 = io_rd_id == 12'h106 ? _GEN_33 : _GEN_232; // @[playground/src/noop/regs.scala 259:44]
  wire [63:0] _GEN_250 = io_rd_id == 12'h106 ? mie : _GEN_233; // @[playground/src/noop/regs.scala 259:44 49:30]
  wire [63:0] _GEN_251 = io_rd_id == 12'h106 ? _GEN_47 : _GEN_234; // @[playground/src/noop/regs.scala 259:44]
  wire [63:0] _GEN_252 = io_rd_id == 12'h106 ? pmpaddr0 : _GEN_235; // @[playground/src/noop/regs.scala 259:44 61:30]
  wire [63:0] _GEN_253 = io_rd_id == 12'h106 ? pmpaddr1 : _GEN_236; // @[playground/src/noop/regs.scala 259:44 62:30]
  wire [63:0] _GEN_254 = io_rd_id == 12'h106 ? pmpaddr2 : _GEN_237; // @[playground/src/noop/regs.scala 259:44 63:30]
  wire [63:0] _GEN_255 = io_rd_id == 12'h106 ? pmpaddr3 : _GEN_238; // @[playground/src/noop/regs.scala 259:44 64:30]
  wire [63:0] _GEN_257 = io_rd_id == 12'h106 ? uscratch : _GEN_240; // @[playground/src/noop/regs.scala 259:44 65:30]
  wire [63:0] _GEN_258 = io_rd_id == 12'h106 ? mhartid : _GEN_241; // @[playground/src/noop/regs.scala 259:44 67:30]
  wire [63:0] _GEN_259 = io_rd_id == 12'h306 ? io_rd_data : {{32'd0}, mcounteren}; // @[playground/src/noop/regs.scala 257:44 258:20 53:30]
  wire [63:0] _GEN_260 = io_rd_id == 12'h306 ? {{32'd0}, scounteren} : _GEN_242; // @[playground/src/noop/regs.scala 257:44 54:30]
  wire [63:0] _GEN_261 = io_rd_id == 12'h306 ? _GEN_35 : _GEN_243; // @[playground/src/noop/regs.scala 257:44]
  wire [63:0] _GEN_262 = io_rd_id == 12'h306 ? _GEN_36 : _GEN_244; // @[playground/src/noop/regs.scala 257:44]
  wire [63:0] _GEN_263 = io_rd_id == 12'h306 ? sscratch : _GEN_245; // @[playground/src/noop/regs.scala 257:44 57:30]
  wire [63:0] _GEN_264 = io_rd_id == 12'h306 ? stvec : _GEN_246; // @[playground/src/noop/regs.scala 257:44 58:30]
  wire [63:0] _GEN_265 = io_rd_id == 12'h306 ? satp : _GEN_247; // @[playground/src/noop/regs.scala 257:44 59:30]
  wire [63:0] _GEN_266 = io_rd_id == 12'h306 ? _GEN_34 : _GEN_248; // @[playground/src/noop/regs.scala 257:44]
  wire [63:0] _GEN_267 = io_rd_id == 12'h306 ? _GEN_33 : _GEN_249; // @[playground/src/noop/regs.scala 257:44]
  wire [63:0] _GEN_268 = io_rd_id == 12'h306 ? mie : _GEN_250; // @[playground/src/noop/regs.scala 257:44 49:30]
  wire [63:0] _GEN_269 = io_rd_id == 12'h306 ? _GEN_47 : _GEN_251; // @[playground/src/noop/regs.scala 257:44]
  wire [63:0] _GEN_270 = io_rd_id == 12'h306 ? pmpaddr0 : _GEN_252; // @[playground/src/noop/regs.scala 257:44 61:30]
  wire [63:0] _GEN_271 = io_rd_id == 12'h306 ? pmpaddr1 : _GEN_253; // @[playground/src/noop/regs.scala 257:44 62:30]
  wire [63:0] _GEN_272 = io_rd_id == 12'h306 ? pmpaddr2 : _GEN_254; // @[playground/src/noop/regs.scala 257:44 63:30]
  wire [63:0] _GEN_273 = io_rd_id == 12'h306 ? pmpaddr3 : _GEN_255; // @[playground/src/noop/regs.scala 257:44 64:30]
  wire [63:0] _GEN_275 = io_rd_id == 12'h306 ? uscratch : _GEN_257; // @[playground/src/noop/regs.scala 257:44 65:30]
  wire [63:0] _GEN_276 = io_rd_id == 12'h306 ? mhartid : _GEN_258; // @[playground/src/noop/regs.scala 257:44 67:30]
  wire [63:0] _GEN_277 = io_rd_id == 12'h303 ? _mideleg_T : mideleg; // @[playground/src/noop/regs.scala 255:41 256:17 52:30]
  wire [63:0] _GEN_278 = io_rd_id == 12'h303 ? {{32'd0}, mcounteren} : _GEN_259; // @[playground/src/noop/regs.scala 255:41 53:30]
  wire [63:0] _GEN_279 = io_rd_id == 12'h303 ? {{32'd0}, scounteren} : _GEN_260; // @[playground/src/noop/regs.scala 255:41 54:30]
  wire [63:0] _GEN_280 = io_rd_id == 12'h303 ? _GEN_35 : _GEN_261; // @[playground/src/noop/regs.scala 255:41]
  wire [63:0] _GEN_281 = io_rd_id == 12'h303 ? _GEN_36 : _GEN_262; // @[playground/src/noop/regs.scala 255:41]
  wire [63:0] _GEN_282 = io_rd_id == 12'h303 ? sscratch : _GEN_263; // @[playground/src/noop/regs.scala 255:41 57:30]
  wire [63:0] _GEN_283 = io_rd_id == 12'h303 ? stvec : _GEN_264; // @[playground/src/noop/regs.scala 255:41 58:30]
  wire [63:0] _GEN_284 = io_rd_id == 12'h303 ? satp : _GEN_265; // @[playground/src/noop/regs.scala 255:41 59:30]
  wire [63:0] _GEN_285 = io_rd_id == 12'h303 ? _GEN_34 : _GEN_266; // @[playground/src/noop/regs.scala 255:41]
  wire [63:0] _GEN_286 = io_rd_id == 12'h303 ? _GEN_33 : _GEN_267; // @[playground/src/noop/regs.scala 255:41]
  wire [63:0] _GEN_287 = io_rd_id == 12'h303 ? mie : _GEN_268; // @[playground/src/noop/regs.scala 255:41 49:30]
  wire [63:0] _GEN_288 = io_rd_id == 12'h303 ? _GEN_47 : _GEN_269; // @[playground/src/noop/regs.scala 255:41]
  wire [63:0] _GEN_289 = io_rd_id == 12'h303 ? pmpaddr0 : _GEN_270; // @[playground/src/noop/regs.scala 255:41 61:30]
  wire [63:0] _GEN_290 = io_rd_id == 12'h303 ? pmpaddr1 : _GEN_271; // @[playground/src/noop/regs.scala 255:41 62:30]
  wire [63:0] _GEN_291 = io_rd_id == 12'h303 ? pmpaddr2 : _GEN_272; // @[playground/src/noop/regs.scala 255:41 63:30]
  wire [63:0] _GEN_292 = io_rd_id == 12'h303 ? pmpaddr3 : _GEN_273; // @[playground/src/noop/regs.scala 255:41 64:30]
  wire [63:0] _GEN_294 = io_rd_id == 12'h303 ? uscratch : _GEN_275; // @[playground/src/noop/regs.scala 255:41 65:30]
  wire [63:0] _GEN_295 = io_rd_id == 12'h303 ? mhartid : _GEN_276; // @[playground/src/noop/regs.scala 255:41 67:30]
  wire [63:0] _GEN_296 = io_rd_id == 12'h302 ? _medeleg_T : medeleg; // @[playground/src/noop/regs.scala 253:41 254:17 51:30]
  wire [63:0] _GEN_297 = io_rd_id == 12'h302 ? mideleg : _GEN_277; // @[playground/src/noop/regs.scala 253:41 52:30]
  wire [63:0] _GEN_298 = io_rd_id == 12'h302 ? {{32'd0}, mcounteren} : _GEN_278; // @[playground/src/noop/regs.scala 253:41 53:30]
  wire [63:0] _GEN_299 = io_rd_id == 12'h302 ? {{32'd0}, scounteren} : _GEN_279; // @[playground/src/noop/regs.scala 253:41 54:30]
  wire [63:0] _GEN_300 = io_rd_id == 12'h302 ? _GEN_35 : _GEN_280; // @[playground/src/noop/regs.scala 253:41]
  wire [63:0] _GEN_301 = io_rd_id == 12'h302 ? _GEN_36 : _GEN_281; // @[playground/src/noop/regs.scala 253:41]
  wire [63:0] _GEN_302 = io_rd_id == 12'h302 ? sscratch : _GEN_282; // @[playground/src/noop/regs.scala 253:41 57:30]
  wire [63:0] _GEN_303 = io_rd_id == 12'h302 ? stvec : _GEN_283; // @[playground/src/noop/regs.scala 253:41 58:30]
  wire [63:0] _GEN_304 = io_rd_id == 12'h302 ? satp : _GEN_284; // @[playground/src/noop/regs.scala 253:41 59:30]
  wire [63:0] _GEN_305 = io_rd_id == 12'h302 ? _GEN_34 : _GEN_285; // @[playground/src/noop/regs.scala 253:41]
  wire [63:0] _GEN_306 = io_rd_id == 12'h302 ? _GEN_33 : _GEN_286; // @[playground/src/noop/regs.scala 253:41]
  wire [63:0] _GEN_307 = io_rd_id == 12'h302 ? mie : _GEN_287; // @[playground/src/noop/regs.scala 253:41 49:30]
  wire [63:0] _GEN_308 = io_rd_id == 12'h302 ? _GEN_47 : _GEN_288; // @[playground/src/noop/regs.scala 253:41]
  wire [63:0] _GEN_309 = io_rd_id == 12'h302 ? pmpaddr0 : _GEN_289; // @[playground/src/noop/regs.scala 253:41 61:30]
  wire [63:0] _GEN_310 = io_rd_id == 12'h302 ? pmpaddr1 : _GEN_290; // @[playground/src/noop/regs.scala 253:41 62:30]
  wire [63:0] _GEN_311 = io_rd_id == 12'h302 ? pmpaddr2 : _GEN_291; // @[playground/src/noop/regs.scala 253:41 63:30]
  wire [63:0] _GEN_312 = io_rd_id == 12'h302 ? pmpaddr3 : _GEN_292; // @[playground/src/noop/regs.scala 253:41 64:30]
  wire [63:0] _GEN_314 = io_rd_id == 12'h302 ? uscratch : _GEN_294; // @[playground/src/noop/regs.scala 253:41 65:30]
  wire [63:0] _GEN_315 = io_rd_id == 12'h302 ? mhartid : _GEN_295; // @[playground/src/noop/regs.scala 253:41 67:30]
  wire [63:0] _GEN_316 = io_rd_id == 12'h342 ? io_rd_data : _GEN_37; // @[playground/src/noop/regs.scala 251:40 252:16]
  wire [63:0] _GEN_317 = io_rd_id == 12'h342 ? medeleg : _GEN_296; // @[playground/src/noop/regs.scala 251:40 51:30]
  wire [63:0] _GEN_318 = io_rd_id == 12'h342 ? mideleg : _GEN_297; // @[playground/src/noop/regs.scala 251:40 52:30]
  wire [63:0] _GEN_319 = io_rd_id == 12'h342 ? {{32'd0}, mcounteren} : _GEN_298; // @[playground/src/noop/regs.scala 251:40 53:30]
  wire [63:0] _GEN_320 = io_rd_id == 12'h342 ? {{32'd0}, scounteren} : _GEN_299; // @[playground/src/noop/regs.scala 251:40 54:30]
  wire [63:0] _GEN_321 = io_rd_id == 12'h342 ? _GEN_35 : _GEN_300; // @[playground/src/noop/regs.scala 251:40]
  wire [63:0] _GEN_322 = io_rd_id == 12'h342 ? _GEN_36 : _GEN_301; // @[playground/src/noop/regs.scala 251:40]
  wire [63:0] _GEN_323 = io_rd_id == 12'h342 ? sscratch : _GEN_302; // @[playground/src/noop/regs.scala 251:40 57:30]
  wire [63:0] _GEN_324 = io_rd_id == 12'h342 ? stvec : _GEN_303; // @[playground/src/noop/regs.scala 251:40 58:30]
  wire [63:0] _GEN_325 = io_rd_id == 12'h342 ? satp : _GEN_304; // @[playground/src/noop/regs.scala 251:40 59:30]
  wire [63:0] _GEN_326 = io_rd_id == 12'h342 ? _GEN_34 : _GEN_305; // @[playground/src/noop/regs.scala 251:40]
  wire [63:0] _GEN_327 = io_rd_id == 12'h342 ? _GEN_33 : _GEN_306; // @[playground/src/noop/regs.scala 251:40]
  wire [63:0] _GEN_328 = io_rd_id == 12'h342 ? mie : _GEN_307; // @[playground/src/noop/regs.scala 251:40 49:30]
  wire [63:0] _GEN_329 = io_rd_id == 12'h342 ? _GEN_47 : _GEN_308; // @[playground/src/noop/regs.scala 251:40]
  wire [63:0] _GEN_330 = io_rd_id == 12'h342 ? pmpaddr0 : _GEN_309; // @[playground/src/noop/regs.scala 251:40 61:30]
  wire [63:0] _GEN_331 = io_rd_id == 12'h342 ? pmpaddr1 : _GEN_310; // @[playground/src/noop/regs.scala 251:40 62:30]
  wire [63:0] _GEN_332 = io_rd_id == 12'h342 ? pmpaddr2 : _GEN_311; // @[playground/src/noop/regs.scala 251:40 63:30]
  wire [63:0] _GEN_333 = io_rd_id == 12'h342 ? pmpaddr3 : _GEN_312; // @[playground/src/noop/regs.scala 251:40 64:30]
  wire [63:0] _GEN_335 = io_rd_id == 12'h342 ? uscratch : _GEN_314; // @[playground/src/noop/regs.scala 251:40 65:30]
  wire [63:0] _GEN_336 = io_rd_id == 12'h342 ? mhartid : _GEN_315; // @[playground/src/noop/regs.scala 251:40 67:30]
  wire [63:0] _GEN_337 = io_rd_id == 12'h344 ? _mip_T_32 : _GEN_329; // @[playground/src/noop/regs.scala 249:37 250:13]
  wire [63:0] _GEN_338 = io_rd_id == 12'h344 ? _GEN_37 : _GEN_316; // @[playground/src/noop/regs.scala 249:37]
  wire [63:0] _GEN_339 = io_rd_id == 12'h344 ? medeleg : _GEN_317; // @[playground/src/noop/regs.scala 249:37 51:30]
  wire [63:0] _GEN_340 = io_rd_id == 12'h344 ? mideleg : _GEN_318; // @[playground/src/noop/regs.scala 249:37 52:30]
  wire [63:0] _GEN_341 = io_rd_id == 12'h344 ? {{32'd0}, mcounteren} : _GEN_319; // @[playground/src/noop/regs.scala 249:37 53:30]
  wire [63:0] _GEN_342 = io_rd_id == 12'h344 ? {{32'd0}, scounteren} : _GEN_320; // @[playground/src/noop/regs.scala 249:37 54:30]
  wire [63:0] _GEN_343 = io_rd_id == 12'h344 ? _GEN_35 : _GEN_321; // @[playground/src/noop/regs.scala 249:37]
  wire [63:0] _GEN_344 = io_rd_id == 12'h344 ? _GEN_36 : _GEN_322; // @[playground/src/noop/regs.scala 249:37]
  wire [63:0] _GEN_345 = io_rd_id == 12'h344 ? sscratch : _GEN_323; // @[playground/src/noop/regs.scala 249:37 57:30]
  wire [63:0] _GEN_346 = io_rd_id == 12'h344 ? stvec : _GEN_324; // @[playground/src/noop/regs.scala 249:37 58:30]
  wire [63:0] _GEN_347 = io_rd_id == 12'h344 ? satp : _GEN_325; // @[playground/src/noop/regs.scala 249:37 59:30]
  wire [63:0] _GEN_348 = io_rd_id == 12'h344 ? _GEN_34 : _GEN_326; // @[playground/src/noop/regs.scala 249:37]
  wire [63:0] _GEN_349 = io_rd_id == 12'h344 ? _GEN_33 : _GEN_327; // @[playground/src/noop/regs.scala 249:37]
  wire [63:0] _GEN_350 = io_rd_id == 12'h344 ? mie : _GEN_328; // @[playground/src/noop/regs.scala 249:37 49:30]
  wire [63:0] _GEN_351 = io_rd_id == 12'h344 ? pmpaddr0 : _GEN_330; // @[playground/src/noop/regs.scala 249:37 61:30]
  wire [63:0] _GEN_352 = io_rd_id == 12'h344 ? pmpaddr1 : _GEN_331; // @[playground/src/noop/regs.scala 249:37 62:30]
  wire [63:0] _GEN_353 = io_rd_id == 12'h344 ? pmpaddr2 : _GEN_332; // @[playground/src/noop/regs.scala 249:37 63:30]
  wire [63:0] _GEN_354 = io_rd_id == 12'h344 ? pmpaddr3 : _GEN_333; // @[playground/src/noop/regs.scala 249:37 64:30]
  wire [63:0] _GEN_356 = io_rd_id == 12'h344 ? uscratch : _GEN_335; // @[playground/src/noop/regs.scala 249:37 65:30]
  wire [63:0] _GEN_357 = io_rd_id == 12'h344 ? mhartid : _GEN_336; // @[playground/src/noop/regs.scala 249:37 67:30]
  wire [63:0] _GEN_358 = io_rd_id == 12'h304 ? io_rd_data : _GEN_350; // @[playground/src/noop/regs.scala 247:37 248:13]
  wire [63:0] _GEN_359 = io_rd_id == 12'h304 ? _GEN_47 : _GEN_337; // @[playground/src/noop/regs.scala 247:37]
  wire [63:0] _GEN_360 = io_rd_id == 12'h304 ? _GEN_37 : _GEN_338; // @[playground/src/noop/regs.scala 247:37]
  wire [63:0] _GEN_361 = io_rd_id == 12'h304 ? medeleg : _GEN_339; // @[playground/src/noop/regs.scala 247:37 51:30]
  wire [63:0] _GEN_362 = io_rd_id == 12'h304 ? mideleg : _GEN_340; // @[playground/src/noop/regs.scala 247:37 52:30]
  wire [63:0] _GEN_363 = io_rd_id == 12'h304 ? {{32'd0}, mcounteren} : _GEN_341; // @[playground/src/noop/regs.scala 247:37 53:30]
  wire [63:0] _GEN_364 = io_rd_id == 12'h304 ? {{32'd0}, scounteren} : _GEN_342; // @[playground/src/noop/regs.scala 247:37 54:30]
  wire [63:0] _GEN_365 = io_rd_id == 12'h304 ? _GEN_35 : _GEN_343; // @[playground/src/noop/regs.scala 247:37]
  wire [63:0] _GEN_366 = io_rd_id == 12'h304 ? _GEN_36 : _GEN_344; // @[playground/src/noop/regs.scala 247:37]
  wire [63:0] _GEN_367 = io_rd_id == 12'h304 ? sscratch : _GEN_345; // @[playground/src/noop/regs.scala 247:37 57:30]
  wire [63:0] _GEN_368 = io_rd_id == 12'h304 ? stvec : _GEN_346; // @[playground/src/noop/regs.scala 247:37 58:30]
  wire [63:0] _GEN_369 = io_rd_id == 12'h304 ? satp : _GEN_347; // @[playground/src/noop/regs.scala 247:37 59:30]
  wire [63:0] _GEN_370 = io_rd_id == 12'h304 ? _GEN_34 : _GEN_348; // @[playground/src/noop/regs.scala 247:37]
  wire [63:0] _GEN_371 = io_rd_id == 12'h304 ? _GEN_33 : _GEN_349; // @[playground/src/noop/regs.scala 247:37]
  wire [63:0] _GEN_372 = io_rd_id == 12'h304 ? pmpaddr0 : _GEN_351; // @[playground/src/noop/regs.scala 247:37 61:30]
  wire [63:0] _GEN_373 = io_rd_id == 12'h304 ? pmpaddr1 : _GEN_352; // @[playground/src/noop/regs.scala 247:37 62:30]
  wire [63:0] _GEN_374 = io_rd_id == 12'h304 ? pmpaddr2 : _GEN_353; // @[playground/src/noop/regs.scala 247:37 63:30]
  wire [63:0] _GEN_375 = io_rd_id == 12'h304 ? pmpaddr3 : _GEN_354; // @[playground/src/noop/regs.scala 247:37 64:30]
  wire [63:0] _GEN_377 = io_rd_id == 12'h304 ? uscratch : _GEN_356; // @[playground/src/noop/regs.scala 247:37 65:30]
  wire [63:0] _GEN_378 = io_rd_id == 12'h304 ? mhartid : _GEN_357; // @[playground/src/noop/regs.scala 247:37 67:30]
  wire [63:0] _GEN_379 = io_rd_id == 12'h305 ? io_rd_data : mtvec; // @[playground/src/noop/regs.scala 245:39 246:15 48:30]
  wire [63:0] _GEN_380 = io_rd_id == 12'h305 ? mie : _GEN_358; // @[playground/src/noop/regs.scala 245:39 49:30]
  wire [63:0] _GEN_381 = io_rd_id == 12'h305 ? _GEN_47 : _GEN_359; // @[playground/src/noop/regs.scala 245:39]
  wire [63:0] _GEN_382 = io_rd_id == 12'h305 ? _GEN_37 : _GEN_360; // @[playground/src/noop/regs.scala 245:39]
  wire [63:0] _GEN_383 = io_rd_id == 12'h305 ? medeleg : _GEN_361; // @[playground/src/noop/regs.scala 245:39 51:30]
  wire [63:0] _GEN_384 = io_rd_id == 12'h305 ? mideleg : _GEN_362; // @[playground/src/noop/regs.scala 245:39 52:30]
  wire [63:0] _GEN_385 = io_rd_id == 12'h305 ? {{32'd0}, mcounteren} : _GEN_363; // @[playground/src/noop/regs.scala 245:39 53:30]
  wire [63:0] _GEN_386 = io_rd_id == 12'h305 ? {{32'd0}, scounteren} : _GEN_364; // @[playground/src/noop/regs.scala 245:39 54:30]
  wire [63:0] _GEN_387 = io_rd_id == 12'h305 ? _GEN_35 : _GEN_365; // @[playground/src/noop/regs.scala 245:39]
  wire [63:0] _GEN_388 = io_rd_id == 12'h305 ? _GEN_36 : _GEN_366; // @[playground/src/noop/regs.scala 245:39]
  wire [63:0] _GEN_389 = io_rd_id == 12'h305 ? sscratch : _GEN_367; // @[playground/src/noop/regs.scala 245:39 57:30]
  wire [63:0] _GEN_390 = io_rd_id == 12'h305 ? stvec : _GEN_368; // @[playground/src/noop/regs.scala 245:39 58:30]
  wire [63:0] _GEN_391 = io_rd_id == 12'h305 ? satp : _GEN_369; // @[playground/src/noop/regs.scala 245:39 59:30]
  wire [63:0] _GEN_392 = io_rd_id == 12'h305 ? _GEN_34 : _GEN_370; // @[playground/src/noop/regs.scala 245:39]
  wire [63:0] _GEN_393 = io_rd_id == 12'h305 ? _GEN_33 : _GEN_371; // @[playground/src/noop/regs.scala 245:39]
  wire [63:0] _GEN_394 = io_rd_id == 12'h305 ? pmpaddr0 : _GEN_372; // @[playground/src/noop/regs.scala 245:39 61:30]
  wire [63:0] _GEN_395 = io_rd_id == 12'h305 ? pmpaddr1 : _GEN_373; // @[playground/src/noop/regs.scala 245:39 62:30]
  wire [63:0] _GEN_396 = io_rd_id == 12'h305 ? pmpaddr2 : _GEN_374; // @[playground/src/noop/regs.scala 245:39 63:30]
  wire [63:0] _GEN_397 = io_rd_id == 12'h305 ? pmpaddr3 : _GEN_375; // @[playground/src/noop/regs.scala 245:39 64:30]
  wire [63:0] _GEN_399 = io_rd_id == 12'h305 ? uscratch : _GEN_377; // @[playground/src/noop/regs.scala 245:39 65:30]
  wire [63:0] _GEN_400 = io_rd_id == 12'h305 ? mhartid : _GEN_378; // @[playground/src/noop/regs.scala 245:39 67:30]
  wire [63:0] _GEN_401 = io_rd_id == 12'h340 ? io_rd_data : mscratch; // @[playground/src/noop/regs.scala 243:42 244:18 46:30]
  wire [63:0] _GEN_402 = io_rd_id == 12'h340 ? mtvec : _GEN_379; // @[playground/src/noop/regs.scala 243:42 48:30]
  wire [63:0] _GEN_403 = io_rd_id == 12'h340 ? mie : _GEN_380; // @[playground/src/noop/regs.scala 243:42 49:30]
  wire [63:0] _GEN_404 = io_rd_id == 12'h340 ? _GEN_47 : _GEN_381; // @[playground/src/noop/regs.scala 243:42]
  wire [63:0] _GEN_405 = io_rd_id == 12'h340 ? _GEN_37 : _GEN_382; // @[playground/src/noop/regs.scala 243:42]
  wire [63:0] _GEN_406 = io_rd_id == 12'h340 ? medeleg : _GEN_383; // @[playground/src/noop/regs.scala 243:42 51:30]
  wire [63:0] _GEN_407 = io_rd_id == 12'h340 ? mideleg : _GEN_384; // @[playground/src/noop/regs.scala 243:42 52:30]
  wire [63:0] _GEN_408 = io_rd_id == 12'h340 ? {{32'd0}, mcounteren} : _GEN_385; // @[playground/src/noop/regs.scala 243:42 53:30]
  wire [63:0] _GEN_409 = io_rd_id == 12'h340 ? {{32'd0}, scounteren} : _GEN_386; // @[playground/src/noop/regs.scala 243:42 54:30]
  wire [63:0] _GEN_410 = io_rd_id == 12'h340 ? _GEN_35 : _GEN_387; // @[playground/src/noop/regs.scala 243:42]
  wire [63:0] _GEN_411 = io_rd_id == 12'h340 ? _GEN_36 : _GEN_388; // @[playground/src/noop/regs.scala 243:42]
  wire [63:0] _GEN_412 = io_rd_id == 12'h340 ? sscratch : _GEN_389; // @[playground/src/noop/regs.scala 243:42 57:30]
  wire [63:0] _GEN_413 = io_rd_id == 12'h340 ? stvec : _GEN_390; // @[playground/src/noop/regs.scala 243:42 58:30]
  wire [63:0] _GEN_414 = io_rd_id == 12'h340 ? satp : _GEN_391; // @[playground/src/noop/regs.scala 243:42 59:30]
  wire [63:0] _GEN_415 = io_rd_id == 12'h340 ? _GEN_34 : _GEN_392; // @[playground/src/noop/regs.scala 243:42]
  wire [63:0] _GEN_416 = io_rd_id == 12'h340 ? _GEN_33 : _GEN_393; // @[playground/src/noop/regs.scala 243:42]
  wire [63:0] _GEN_417 = io_rd_id == 12'h340 ? pmpaddr0 : _GEN_394; // @[playground/src/noop/regs.scala 243:42 61:30]
  wire [63:0] _GEN_418 = io_rd_id == 12'h340 ? pmpaddr1 : _GEN_395; // @[playground/src/noop/regs.scala 243:42 62:30]
  wire [63:0] _GEN_419 = io_rd_id == 12'h340 ? pmpaddr2 : _GEN_396; // @[playground/src/noop/regs.scala 243:42 63:30]
  wire [63:0] _GEN_420 = io_rd_id == 12'h340 ? pmpaddr3 : _GEN_397; // @[playground/src/noop/regs.scala 243:42 64:30]
  wire [63:0] _GEN_422 = io_rd_id == 12'h340 ? uscratch : _GEN_399; // @[playground/src/noop/regs.scala 243:42 65:30]
  wire [63:0] _GEN_423 = io_rd_id == 12'h340 ? mhartid : _GEN_400; // @[playground/src/noop/regs.scala 243:42 67:30]
  wire [63:0] _GEN_424 = io_rd_id == 12'h343 ? io_rd_data : _GEN_39; // @[playground/src/noop/regs.scala 241:39 242:15]
  wire [63:0] _GEN_425 = io_rd_id == 12'h343 ? mscratch : _GEN_401; // @[playground/src/noop/regs.scala 241:39 46:30]
  wire [63:0] _GEN_426 = io_rd_id == 12'h343 ? mtvec : _GEN_402; // @[playground/src/noop/regs.scala 241:39 48:30]
  wire [63:0] _GEN_427 = io_rd_id == 12'h343 ? mie : _GEN_403; // @[playground/src/noop/regs.scala 241:39 49:30]
  wire [63:0] _GEN_428 = io_rd_id == 12'h343 ? _GEN_47 : _GEN_404; // @[playground/src/noop/regs.scala 241:39]
  wire [63:0] _GEN_429 = io_rd_id == 12'h343 ? _GEN_37 : _GEN_405; // @[playground/src/noop/regs.scala 241:39]
  wire [63:0] _GEN_430 = io_rd_id == 12'h343 ? medeleg : _GEN_406; // @[playground/src/noop/regs.scala 241:39 51:30]
  wire [63:0] _GEN_431 = io_rd_id == 12'h343 ? mideleg : _GEN_407; // @[playground/src/noop/regs.scala 241:39 52:30]
  wire [63:0] _GEN_432 = io_rd_id == 12'h343 ? {{32'd0}, mcounteren} : _GEN_408; // @[playground/src/noop/regs.scala 241:39 53:30]
  wire [63:0] _GEN_433 = io_rd_id == 12'h343 ? {{32'd0}, scounteren} : _GEN_409; // @[playground/src/noop/regs.scala 241:39 54:30]
  wire [63:0] _GEN_434 = io_rd_id == 12'h343 ? _GEN_35 : _GEN_410; // @[playground/src/noop/regs.scala 241:39]
  wire [63:0] _GEN_435 = io_rd_id == 12'h343 ? _GEN_36 : _GEN_411; // @[playground/src/noop/regs.scala 241:39]
  wire [63:0] _GEN_436 = io_rd_id == 12'h343 ? sscratch : _GEN_412; // @[playground/src/noop/regs.scala 241:39 57:30]
  wire [63:0] _GEN_437 = io_rd_id == 12'h343 ? stvec : _GEN_413; // @[playground/src/noop/regs.scala 241:39 58:30]
  wire [63:0] _GEN_438 = io_rd_id == 12'h343 ? satp : _GEN_414; // @[playground/src/noop/regs.scala 241:39 59:30]
  wire [63:0] _GEN_439 = io_rd_id == 12'h343 ? _GEN_34 : _GEN_415; // @[playground/src/noop/regs.scala 241:39]
  wire [63:0] _GEN_440 = io_rd_id == 12'h343 ? _GEN_33 : _GEN_416; // @[playground/src/noop/regs.scala 241:39]
  wire [63:0] _GEN_441 = io_rd_id == 12'h343 ? pmpaddr0 : _GEN_417; // @[playground/src/noop/regs.scala 241:39 61:30]
  wire [63:0] _GEN_442 = io_rd_id == 12'h343 ? pmpaddr1 : _GEN_418; // @[playground/src/noop/regs.scala 241:39 62:30]
  wire [63:0] _GEN_443 = io_rd_id == 12'h343 ? pmpaddr2 : _GEN_419; // @[playground/src/noop/regs.scala 241:39 63:30]
  wire [63:0] _GEN_444 = io_rd_id == 12'h343 ? pmpaddr3 : _GEN_420; // @[playground/src/noop/regs.scala 241:39 64:30]
  wire [63:0] _GEN_446 = io_rd_id == 12'h343 ? uscratch : _GEN_422; // @[playground/src/noop/regs.scala 241:39 65:30]
  wire [63:0] _GEN_447 = io_rd_id == 12'h343 ? mhartid : _GEN_423; // @[playground/src/noop/regs.scala 241:39 67:30]
  wire [63:0] _GEN_448 = io_rd_id == 12'h341 ? io_rd_data : _GEN_38; // @[playground/src/noop/regs.scala 239:38 240:14]
  wire [63:0] _GEN_449 = io_rd_id == 12'h341 ? _GEN_39 : _GEN_424; // @[playground/src/noop/regs.scala 239:38]
  wire [63:0] _GEN_450 = io_rd_id == 12'h341 ? mscratch : _GEN_425; // @[playground/src/noop/regs.scala 239:38 46:30]
  wire [63:0] _GEN_451 = io_rd_id == 12'h341 ? mtvec : _GEN_426; // @[playground/src/noop/regs.scala 239:38 48:30]
  wire [63:0] _GEN_452 = io_rd_id == 12'h341 ? mie : _GEN_427; // @[playground/src/noop/regs.scala 239:38 49:30]
  wire [63:0] _GEN_453 = io_rd_id == 12'h341 ? _GEN_47 : _GEN_428; // @[playground/src/noop/regs.scala 239:38]
  wire [63:0] _GEN_454 = io_rd_id == 12'h341 ? _GEN_37 : _GEN_429; // @[playground/src/noop/regs.scala 239:38]
  wire [63:0] _GEN_455 = io_rd_id == 12'h341 ? medeleg : _GEN_430; // @[playground/src/noop/regs.scala 239:38 51:30]
  wire [63:0] _GEN_456 = io_rd_id == 12'h341 ? mideleg : _GEN_431; // @[playground/src/noop/regs.scala 239:38 52:30]
  wire [63:0] _GEN_457 = io_rd_id == 12'h341 ? {{32'd0}, mcounteren} : _GEN_432; // @[playground/src/noop/regs.scala 239:38 53:30]
  wire [63:0] _GEN_458 = io_rd_id == 12'h341 ? {{32'd0}, scounteren} : _GEN_433; // @[playground/src/noop/regs.scala 239:38 54:30]
  wire [63:0] _GEN_459 = io_rd_id == 12'h341 ? _GEN_35 : _GEN_434; // @[playground/src/noop/regs.scala 239:38]
  wire [63:0] _GEN_460 = io_rd_id == 12'h341 ? _GEN_36 : _GEN_435; // @[playground/src/noop/regs.scala 239:38]
  wire [63:0] _GEN_461 = io_rd_id == 12'h341 ? sscratch : _GEN_436; // @[playground/src/noop/regs.scala 239:38 57:30]
  wire [63:0] _GEN_462 = io_rd_id == 12'h341 ? stvec : _GEN_437; // @[playground/src/noop/regs.scala 239:38 58:30]
  wire [63:0] _GEN_463 = io_rd_id == 12'h341 ? satp : _GEN_438; // @[playground/src/noop/regs.scala 239:38 59:30]
  wire [63:0] _GEN_464 = io_rd_id == 12'h341 ? _GEN_34 : _GEN_439; // @[playground/src/noop/regs.scala 239:38]
  wire [63:0] _GEN_465 = io_rd_id == 12'h341 ? _GEN_33 : _GEN_440; // @[playground/src/noop/regs.scala 239:38]
  wire [63:0] _GEN_466 = io_rd_id == 12'h341 ? pmpaddr0 : _GEN_441; // @[playground/src/noop/regs.scala 239:38 61:30]
  wire [63:0] _GEN_467 = io_rd_id == 12'h341 ? pmpaddr1 : _GEN_442; // @[playground/src/noop/regs.scala 239:38 62:30]
  wire [63:0] _GEN_468 = io_rd_id == 12'h341 ? pmpaddr2 : _GEN_443; // @[playground/src/noop/regs.scala 239:38 63:30]
  wire [63:0] _GEN_469 = io_rd_id == 12'h341 ? pmpaddr3 : _GEN_444; // @[playground/src/noop/regs.scala 239:38 64:30]
  wire [63:0] _GEN_471 = io_rd_id == 12'h341 ? uscratch : _GEN_446; // @[playground/src/noop/regs.scala 239:38 65:30]
  wire [63:0] _GEN_472 = io_rd_id == 12'h341 ? mhartid : _GEN_447; // @[playground/src/noop/regs.scala 239:38 67:30]
  wire [63:0] _GEN_483 = io_rd_id == 12'h300 ? {{32'd0}, mcounteren} : _GEN_457; // @[playground/src/noop/regs.scala 235:41 53:30]
  wire [63:0] _GEN_484 = io_rd_id == 12'h300 ? {{32'd0}, scounteren} : _GEN_458; // @[playground/src/noop/regs.scala 235:41 54:30]
  wire [63:0] _GEN_509 = io_rd_id == 12'h301 ? {{32'd0}, mcounteren} : _GEN_483; // @[playground/src/noop/regs.scala 233:38 53:30]
  wire [63:0] _GEN_510 = io_rd_id == 12'h301 ? {{32'd0}, scounteren} : _GEN_484; // @[playground/src/noop/regs.scala 233:38 54:30]
  wire [63:0] _GEN_535 = ~io_rd_en ? {{32'd0}, mcounteren} : _GEN_509; // @[playground/src/noop/regs.scala 232:20 53:30]
  wire [63:0] _GEN_536 = ~io_rd_en ? {{32'd0}, scounteren} : _GEN_510; // @[playground/src/noop/regs.scala 232:20 54:30]
  wire [73:0] _updateCsrs_io_mstatus_T = {10'h300,mstatus}; // @[playground/src/noop/regs.scala 300:35]
  wire [73:0] _updateCsrs_io_mepc_T = {10'h341,mepc}; // @[playground/src/noop/regs.scala 301:35]
  wire [73:0] _updateCsrs_io_mtval_T = {10'h343,mtval}; // @[playground/src/noop/regs.scala 302:35]
  wire [73:0] _updateCsrs_io_mscratch_T = {10'h340,mscratch}; // @[playground/src/noop/regs.scala 303:35]
  wire [73:0] _updateCsrs_io_mcause_T = {10'h342,mcause}; // @[playground/src/noop/regs.scala 304:35]
  wire [73:0] _updateCsrs_io_mtvec_T = {10'h305,mtvec}; // @[playground/src/noop/regs.scala 305:35]
  wire [73:0] _updateCsrs_io_mie_T = {10'h304,mie}; // @[playground/src/noop/regs.scala 306:35]
  wire [73:0] _updateCsrs_io_mip_T = {10'h344,mip}; // @[playground/src/noop/regs.scala 307:35]
  wire [73:0] _updateCsrs_io_medeleg_T = {10'h302,medeleg}; // @[playground/src/noop/regs.scala 308:35]
  wire [73:0] _updateCsrs_io_mideleg_T = {10'h303,mideleg}; // @[playground/src/noop/regs.scala 309:35]
  wire [72:0] _updateCsrs_io_sepc_T = {9'h141,sepc}; // @[playground/src/noop/regs.scala 310:35]
  wire [72:0] _updateCsrs_io_stval_T = {9'h143,stval}; // @[playground/src/noop/regs.scala 311:35]
  wire [72:0] _updateCsrs_io_sscratch_T = {9'h140,sscratch}; // @[playground/src/noop/regs.scala 312:35]
  wire [72:0] _updateCsrs_io_stvec_T = {9'h105,stvec}; // @[playground/src/noop/regs.scala 313:35]
  wire [72:0] _updateCsrs_io_satp_T = {9'h180,satp}; // @[playground/src/noop/regs.scala 314:35]
  wire [72:0] _updateCsrs_io_scause_T = {9'h142,scause}; // @[playground/src/noop/regs.scala 315:35]
  wire [63:0] _GEN_181 = reset ? 64'h0 : _GEN_535; // @[playground/src/noop/regs.scala 53:{30,30}]
  wire [63:0] _GEN_194 = reset ? 64'h0 : _GEN_536; // @[playground/src/noop/regs.scala 54:{30,30}]
  wire [66:0] _GEN_208 = reset ? 67'h0 : _GEN_30; // @[playground/src/noop/regs.scala 74:{34,34}]
  UpdateCsrs updateCsrs ( // @[playground/src/noop/regs.scala 298:28]
    .priv(updateCsrs_priv),
    .mstatus(updateCsrs_mstatus),
    .mepc(updateCsrs_mepc),
    .mtval(updateCsrs_mtval),
    .mscratch(updateCsrs_mscratch),
    .mcause(updateCsrs_mcause),
    .mtvec(updateCsrs_mtvec),
    .mie(updateCsrs_mie),
    .mip(updateCsrs_mip),
    .medeleg(updateCsrs_medeleg),
    .mideleg(updateCsrs_mideleg),
    .sepc(updateCsrs_sepc),
    .stval(updateCsrs_stval),
    .sscratch(updateCsrs_sscratch),
    .stvec(updateCsrs_stvec),
    .satp(updateCsrs_satp),
    .scause(updateCsrs_scause),
    .clock(updateCsrs_clock)
  );
  assign io_rs_data = io_rs_id == 12'h301 ? misa : _GEN_102; // @[playground/src/noop/regs.scala 170:32 171:20]
  assign io_rs_is_err = io_rs_id == 12'h301 ? 1'h0 : _GEN_103; // @[playground/src/noop/regs.scala 169:21 170:32]
  assign io_mmuState_priv = priv; // @[playground/src/noop/regs.scala 70:25]
  assign io_mmuState_mstatus = mstatus; // @[playground/src/noop/regs.scala 71:25]
  assign io_mmuState_satp = satp; // @[playground/src/noop/regs.scala 72:25]
  assign io_idState_priv = priv; // @[playground/src/noop/regs.scala 73:24]
  assign io_reg2if_seq_pc = forceJmp_seq_pc; // @[playground/src/noop/regs.scala 75:25]
  assign io_reg2if_valid = forceJmp_valid; // @[playground/src/noop/regs.scala 75:25]
  assign io_intr_out_en = intr_out_r_en; // @[playground/src/noop/regs.scala 124:17]
  assign io_intr_out_cause = intr_out_r_cause; // @[playground/src/noop/regs.scala 124:17]
  assign io_updateNextPc_seq_pc = forceJmp_seq_pc; // @[playground/src/noop/regs.scala 78:25]
  assign io_updateNextPc_valid = forceJmp_valid; // @[playground/src/noop/regs.scala 78:25]
  assign updateCsrs_priv = priv; // @[playground/src/noop/regs.scala 299:29]
  assign updateCsrs_mstatus = {{2'd0}, _updateCsrs_io_mstatus_T}; // @[playground/src/noop/regs.scala 300:29]
  assign updateCsrs_mepc = {{2'd0}, _updateCsrs_io_mepc_T}; // @[playground/src/noop/regs.scala 301:29]
  assign updateCsrs_mtval = {{2'd0}, _updateCsrs_io_mtval_T}; // @[playground/src/noop/regs.scala 302:29]
  assign updateCsrs_mscratch = {{2'd0}, _updateCsrs_io_mscratch_T}; // @[playground/src/noop/regs.scala 303:29]
  assign updateCsrs_mcause = {{2'd0}, _updateCsrs_io_mcause_T}; // @[playground/src/noop/regs.scala 304:29]
  assign updateCsrs_mtvec = {{2'd0}, _updateCsrs_io_mtvec_T}; // @[playground/src/noop/regs.scala 305:29]
  assign updateCsrs_mie = {{2'd0}, _updateCsrs_io_mie_T}; // @[playground/src/noop/regs.scala 306:29]
  assign updateCsrs_mip = {{2'd0}, _updateCsrs_io_mip_T}; // @[playground/src/noop/regs.scala 307:29]
  assign updateCsrs_medeleg = {{2'd0}, _updateCsrs_io_medeleg_T}; // @[playground/src/noop/regs.scala 308:29]
  assign updateCsrs_mideleg = {{2'd0}, _updateCsrs_io_mideleg_T}; // @[playground/src/noop/regs.scala 309:29]
  assign updateCsrs_sepc = {{3'd0}, _updateCsrs_io_sepc_T}; // @[playground/src/noop/regs.scala 310:29]
  assign updateCsrs_stval = {{3'd0}, _updateCsrs_io_stval_T}; // @[playground/src/noop/regs.scala 311:29]
  assign updateCsrs_sscratch = {{3'd0}, _updateCsrs_io_sscratch_T}; // @[playground/src/noop/regs.scala 312:29]
  assign updateCsrs_stvec = {{3'd0}, _updateCsrs_io_stvec_T}; // @[playground/src/noop/regs.scala 313:29]
  assign updateCsrs_satp = {{3'd0}, _updateCsrs_io_satp_T}; // @[playground/src/noop/regs.scala 314:29]
  assign updateCsrs_scause = {{3'd0}, _updateCsrs_io_scause_T}; // @[playground/src/noop/regs.scala 315:29]
  assign updateCsrs_clock = clock; // @[playground/src/noop/regs.scala 316:29]
  always @(posedge clock) begin
    if (reset) begin // @[playground/src/noop/regs.scala 41:30]
      priv <= 2'h3; // @[playground/src/noop/regs.scala 41:30]
    end else if (io_excep_en) begin // @[playground/src/noop/regs.scala 79:22]
      if (io_excep_etype == 2'h2) begin // @[playground/src/noop/regs.scala 80:44]
        priv <= _priv_T_1; // @[playground/src/noop/regs.scala 84:29]
      end else if (io_excep_etype == 2'h3) begin // @[playground/src/noop/regs.scala 87:50]
        priv <= mstatus[12:11]; // @[playground/src/noop/regs.scala 91:29]
      end else begin
        priv <= _GEN_6;
      end
    end
    if (reset) begin // @[playground/src/noop/regs.scala 42:30]
      misa <= 64'h800000000014112d; // @[playground/src/noop/regs.scala 42:30]
    end else if (!(~io_rd_en)) begin // @[playground/src/noop/regs.scala 232:20]
      if (io_rd_id == 12'h301) begin // @[playground/src/noop/regs.scala 233:38]
        misa <= io_rd_data; // @[playground/src/noop/regs.scala 234:14]
      end
    end
    if (reset) begin // @[playground/src/noop/regs.scala 43:30]
      mstatus <= 64'ha00000000; // @[playground/src/noop/regs.scala 43:30]
    end else if (~io_rd_en) begin // @[playground/src/noop/regs.scala 232:20]
      mstatus <= _GEN_33;
    end else if (io_rd_id == 12'h301) begin // @[playground/src/noop/regs.scala 233:38]
      mstatus <= _GEN_33;
    end else if (io_rd_id == 12'h300) begin // @[playground/src/noop/regs.scala 235:41]
      mstatus <= _mstatus_T_13; // @[playground/src/noop/regs.scala 238:17]
    end else begin
      mstatus <= _GEN_465;
    end
    if (reset) begin // @[playground/src/noop/regs.scala 44:30]
      mepc <= 64'h0; // @[playground/src/noop/regs.scala 44:30]
    end else if (~io_rd_en) begin // @[playground/src/noop/regs.scala 232:20]
      mepc <= _GEN_38;
    end else if (io_rd_id == 12'h301) begin // @[playground/src/noop/regs.scala 233:38]
      mepc <= _GEN_38;
    end else if (io_rd_id == 12'h300) begin // @[playground/src/noop/regs.scala 235:41]
      mepc <= _GEN_38;
    end else begin
      mepc <= _GEN_448;
    end
    if (reset) begin // @[playground/src/noop/regs.scala 45:30]
      mtval <= 64'h0; // @[playground/src/noop/regs.scala 45:30]
    end else if (~io_rd_en) begin // @[playground/src/noop/regs.scala 232:20]
      mtval <= _GEN_39;
    end else if (io_rd_id == 12'h301) begin // @[playground/src/noop/regs.scala 233:38]
      mtval <= _GEN_39;
    end else if (io_rd_id == 12'h300) begin // @[playground/src/noop/regs.scala 235:41]
      mtval <= _GEN_39;
    end else begin
      mtval <= _GEN_449;
    end
    if (reset) begin // @[playground/src/noop/regs.scala 46:30]
      mscratch <= 64'h0; // @[playground/src/noop/regs.scala 46:30]
    end else if (!(~io_rd_en)) begin // @[playground/src/noop/regs.scala 232:20]
      if (!(io_rd_id == 12'h301)) begin // @[playground/src/noop/regs.scala 233:38]
        if (!(io_rd_id == 12'h300)) begin // @[playground/src/noop/regs.scala 235:41]
          mscratch <= _GEN_450;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/regs.scala 47:30]
      mcause <= 64'h0; // @[playground/src/noop/regs.scala 47:30]
    end else if (~io_rd_en) begin // @[playground/src/noop/regs.scala 232:20]
      mcause <= _GEN_37;
    end else if (io_rd_id == 12'h301) begin // @[playground/src/noop/regs.scala 233:38]
      mcause <= _GEN_37;
    end else if (io_rd_id == 12'h300) begin // @[playground/src/noop/regs.scala 235:41]
      mcause <= _GEN_37;
    end else begin
      mcause <= _GEN_454;
    end
    if (reset) begin // @[playground/src/noop/regs.scala 48:30]
      mtvec <= 64'h0; // @[playground/src/noop/regs.scala 48:30]
    end else if (!(~io_rd_en)) begin // @[playground/src/noop/regs.scala 232:20]
      if (!(io_rd_id == 12'h301)) begin // @[playground/src/noop/regs.scala 233:38]
        if (!(io_rd_id == 12'h300)) begin // @[playground/src/noop/regs.scala 235:41]
          mtvec <= _GEN_451;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/regs.scala 49:30]
      mie <= 64'h0; // @[playground/src/noop/regs.scala 49:30]
    end else if (!(~io_rd_en)) begin // @[playground/src/noop/regs.scala 232:20]
      if (!(io_rd_id == 12'h301)) begin // @[playground/src/noop/regs.scala 233:38]
        if (!(io_rd_id == 12'h300)) begin // @[playground/src/noop/regs.scala 235:41]
          mie <= _GEN_452;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/regs.scala 50:30]
      mip <= 64'h0; // @[playground/src/noop/regs.scala 50:30]
    end else if (~io_rd_en) begin // @[playground/src/noop/regs.scala 232:20]
      mip <= _GEN_47;
    end else if (io_rd_id == 12'h301) begin // @[playground/src/noop/regs.scala 233:38]
      mip <= _GEN_47;
    end else if (io_rd_id == 12'h300) begin // @[playground/src/noop/regs.scala 235:41]
      mip <= _GEN_47;
    end else begin
      mip <= _GEN_453;
    end
    if (reset) begin // @[playground/src/noop/regs.scala 51:30]
      medeleg <= 64'h0; // @[playground/src/noop/regs.scala 51:30]
    end else if (!(~io_rd_en)) begin // @[playground/src/noop/regs.scala 232:20]
      if (!(io_rd_id == 12'h301)) begin // @[playground/src/noop/regs.scala 233:38]
        if (!(io_rd_id == 12'h300)) begin // @[playground/src/noop/regs.scala 235:41]
          medeleg <= _GEN_455;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/regs.scala 52:30]
      mideleg <= 64'h0; // @[playground/src/noop/regs.scala 52:30]
    end else if (!(~io_rd_en)) begin // @[playground/src/noop/regs.scala 232:20]
      if (!(io_rd_id == 12'h301)) begin // @[playground/src/noop/regs.scala 233:38]
        if (!(io_rd_id == 12'h300)) begin // @[playground/src/noop/regs.scala 235:41]
          mideleg <= _GEN_456;
        end
      end
    end
    mcounteren <= _GEN_181[31:0]; // @[playground/src/noop/regs.scala 53:{30,30}]
    scounteren <= _GEN_194[31:0]; // @[playground/src/noop/regs.scala 54:{30,30}]
    if (reset) begin // @[playground/src/noop/regs.scala 55:30]
      sepc <= 64'h0; // @[playground/src/noop/regs.scala 55:30]
    end else if (~io_rd_en) begin // @[playground/src/noop/regs.scala 232:20]
      sepc <= _GEN_35;
    end else if (io_rd_id == 12'h301) begin // @[playground/src/noop/regs.scala 233:38]
      sepc <= _GEN_35;
    end else if (io_rd_id == 12'h300) begin // @[playground/src/noop/regs.scala 235:41]
      sepc <= _GEN_35;
    end else begin
      sepc <= _GEN_459;
    end
    if (reset) begin // @[playground/src/noop/regs.scala 56:30]
      stval <= 64'h0; // @[playground/src/noop/regs.scala 56:30]
    end else if (~io_rd_en) begin // @[playground/src/noop/regs.scala 232:20]
      stval <= _GEN_36;
    end else if (io_rd_id == 12'h301) begin // @[playground/src/noop/regs.scala 233:38]
      stval <= _GEN_36;
    end else if (io_rd_id == 12'h300) begin // @[playground/src/noop/regs.scala 235:41]
      stval <= _GEN_36;
    end else begin
      stval <= _GEN_460;
    end
    if (reset) begin // @[playground/src/noop/regs.scala 57:30]
      sscratch <= 64'h0; // @[playground/src/noop/regs.scala 57:30]
    end else if (!(~io_rd_en)) begin // @[playground/src/noop/regs.scala 232:20]
      if (!(io_rd_id == 12'h301)) begin // @[playground/src/noop/regs.scala 233:38]
        if (!(io_rd_id == 12'h300)) begin // @[playground/src/noop/regs.scala 235:41]
          sscratch <= _GEN_461;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/regs.scala 58:30]
      stvec <= 64'h0; // @[playground/src/noop/regs.scala 58:30]
    end else if (!(~io_rd_en)) begin // @[playground/src/noop/regs.scala 232:20]
      if (!(io_rd_id == 12'h301)) begin // @[playground/src/noop/regs.scala 233:38]
        if (!(io_rd_id == 12'h300)) begin // @[playground/src/noop/regs.scala 235:41]
          stvec <= _GEN_462;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/regs.scala 59:30]
      satp <= 64'h0; // @[playground/src/noop/regs.scala 59:30]
    end else if (!(~io_rd_en)) begin // @[playground/src/noop/regs.scala 232:20]
      if (!(io_rd_id == 12'h301)) begin // @[playground/src/noop/regs.scala 233:38]
        if (!(io_rd_id == 12'h300)) begin // @[playground/src/noop/regs.scala 235:41]
          satp <= _GEN_463;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/regs.scala 60:30]
      scause <= 64'h0; // @[playground/src/noop/regs.scala 60:30]
    end else if (~io_rd_en) begin // @[playground/src/noop/regs.scala 232:20]
      scause <= _GEN_34;
    end else if (io_rd_id == 12'h301) begin // @[playground/src/noop/regs.scala 233:38]
      scause <= _GEN_34;
    end else if (io_rd_id == 12'h300) begin // @[playground/src/noop/regs.scala 235:41]
      scause <= _GEN_34;
    end else begin
      scause <= _GEN_464;
    end
    if (reset) begin // @[playground/src/noop/regs.scala 61:30]
      pmpaddr0 <= 64'h0; // @[playground/src/noop/regs.scala 61:30]
    end else if (!(~io_rd_en)) begin // @[playground/src/noop/regs.scala 232:20]
      if (!(io_rd_id == 12'h301)) begin // @[playground/src/noop/regs.scala 233:38]
        if (!(io_rd_id == 12'h300)) begin // @[playground/src/noop/regs.scala 235:41]
          pmpaddr0 <= _GEN_466;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/regs.scala 62:30]
      pmpaddr1 <= 64'h0; // @[playground/src/noop/regs.scala 62:30]
    end else if (!(~io_rd_en)) begin // @[playground/src/noop/regs.scala 232:20]
      if (!(io_rd_id == 12'h301)) begin // @[playground/src/noop/regs.scala 233:38]
        if (!(io_rd_id == 12'h300)) begin // @[playground/src/noop/regs.scala 235:41]
          pmpaddr1 <= _GEN_467;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/regs.scala 63:30]
      pmpaddr2 <= 64'h0; // @[playground/src/noop/regs.scala 63:30]
    end else if (!(~io_rd_en)) begin // @[playground/src/noop/regs.scala 232:20]
      if (!(io_rd_id == 12'h301)) begin // @[playground/src/noop/regs.scala 233:38]
        if (!(io_rd_id == 12'h300)) begin // @[playground/src/noop/regs.scala 235:41]
          pmpaddr2 <= _GEN_468;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/regs.scala 64:30]
      pmpaddr3 <= 64'h0; // @[playground/src/noop/regs.scala 64:30]
    end else if (!(~io_rd_en)) begin // @[playground/src/noop/regs.scala 232:20]
      if (!(io_rd_id == 12'h301)) begin // @[playground/src/noop/regs.scala 233:38]
        if (!(io_rd_id == 12'h300)) begin // @[playground/src/noop/regs.scala 235:41]
          pmpaddr3 <= _GEN_469;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/regs.scala 65:30]
      uscratch <= 64'h0; // @[playground/src/noop/regs.scala 65:30]
    end else if (!(~io_rd_en)) begin // @[playground/src/noop/regs.scala 232:20]
      if (!(io_rd_id == 12'h301)) begin // @[playground/src/noop/regs.scala 233:38]
        if (!(io_rd_id == 12'h300)) begin // @[playground/src/noop/regs.scala 235:41]
          uscratch <= _GEN_471;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/regs.scala 67:30]
      mhartid <= 64'h0; // @[playground/src/noop/regs.scala 67:30]
    end else if (!(~io_rd_en)) begin // @[playground/src/noop/regs.scala 232:20]
      if (!(io_rd_id == 12'h301)) begin // @[playground/src/noop/regs.scala 233:38]
        if (!(io_rd_id == 12'h300)) begin // @[playground/src/noop/regs.scala 235:41]
          mhartid <= _GEN_472;
        end
      end
    end
    forceJmp_seq_pc <= _GEN_208[63:0]; // @[playground/src/noop/regs.scala 74:{34,34}]
    if (reset) begin // @[playground/src/noop/regs.scala 74:34]
      forceJmp_valid <= 1'h0; // @[playground/src/noop/regs.scala 74:34]
    end else begin
      forceJmp_valid <= io_excep_en;
    end
    if (reset) begin // @[playground/src/noop/regs.scala 123:29]
      intr_out_r_en <= 1'h0; // @[playground/src/noop/regs.scala 123:29]
    end else begin
      intr_out_r_en <= enable_int != 64'h0; // @[playground/src/noop/regs.scala 157:19]
    end
    if (reset) begin // @[playground/src/noop/regs.scala 123:29]
      intr_out_r_cause <= 64'h0; // @[playground/src/noop/regs.scala 123:29]
    end else begin
      intr_out_r_cause <= _intr_out_r_cause_T_13; // @[playground/src/noop/regs.scala 159:22]
    end
    if (reset) begin // @[playground/src/noop/regs.scala 125:28]
      intr_seip <= 1'h0; // @[playground/src/noop/regs.scala 125:28]
    end else if (io_plic_s_clear) begin // @[playground/src/noop/regs.scala 141:26]
      intr_seip <= 1'h0; // @[playground/src/noop/regs.scala 142:19]
    end else begin
      intr_seip <= _GEN_44;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  priv = _RAND_0[1:0];
  _RAND_1 = {2{`RANDOM}};
  misa = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  mstatus = _RAND_2[63:0];
  _RAND_3 = {2{`RANDOM}};
  mepc = _RAND_3[63:0];
  _RAND_4 = {2{`RANDOM}};
  mtval = _RAND_4[63:0];
  _RAND_5 = {2{`RANDOM}};
  mscratch = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  mcause = _RAND_6[63:0];
  _RAND_7 = {2{`RANDOM}};
  mtvec = _RAND_7[63:0];
  _RAND_8 = {2{`RANDOM}};
  mie = _RAND_8[63:0];
  _RAND_9 = {2{`RANDOM}};
  mip = _RAND_9[63:0];
  _RAND_10 = {2{`RANDOM}};
  medeleg = _RAND_10[63:0];
  _RAND_11 = {2{`RANDOM}};
  mideleg = _RAND_11[63:0];
  _RAND_12 = {1{`RANDOM}};
  mcounteren = _RAND_12[31:0];
  _RAND_13 = {1{`RANDOM}};
  scounteren = _RAND_13[31:0];
  _RAND_14 = {2{`RANDOM}};
  sepc = _RAND_14[63:0];
  _RAND_15 = {2{`RANDOM}};
  stval = _RAND_15[63:0];
  _RAND_16 = {2{`RANDOM}};
  sscratch = _RAND_16[63:0];
  _RAND_17 = {2{`RANDOM}};
  stvec = _RAND_17[63:0];
  _RAND_18 = {2{`RANDOM}};
  satp = _RAND_18[63:0];
  _RAND_19 = {2{`RANDOM}};
  scause = _RAND_19[63:0];
  _RAND_20 = {2{`RANDOM}};
  pmpaddr0 = _RAND_20[63:0];
  _RAND_21 = {2{`RANDOM}};
  pmpaddr1 = _RAND_21[63:0];
  _RAND_22 = {2{`RANDOM}};
  pmpaddr2 = _RAND_22[63:0];
  _RAND_23 = {2{`RANDOM}};
  pmpaddr3 = _RAND_23[63:0];
  _RAND_24 = {2{`RANDOM}};
  uscratch = _RAND_24[63:0];
  _RAND_25 = {2{`RANDOM}};
  mhartid = _RAND_25[63:0];
  _RAND_26 = {2{`RANDOM}};
  forceJmp_seq_pc = _RAND_26[63:0];
  _RAND_27 = {1{`RANDOM}};
  forceJmp_valid = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  intr_out_r_en = _RAND_28[0:0];
  _RAND_29 = {2{`RANDOM}};
  intr_out_r_cause = _RAND_29[63:0];
  _RAND_30 = {1{`RANDOM}};
  intr_seip = _RAND_30[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module S011HD1P_X32Y2D128_BW(
  input          clock,
  input          reset,
  output [127:0] io_Q, // @[playground/src/ram/ram.scala 87:16]
  input          io_CEN, // @[playground/src/ram/ram.scala 87:16]
  input          io_WEN, // @[playground/src/ram/ram.scala 87:16]
  input  [127:0] io_BWEN, // @[playground/src/ram/ram.scala 87:16]
  input  [5:0]   io_A, // @[playground/src/ram/ram.scala 87:16]
  input  [127:0] io_D // @[playground/src/ram/ram.scala 87:16]
);
`ifdef RANDOMIZE_MEM_INIT
  reg [127:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [127:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg [127:0] ram [0:63]; // @[playground/src/ram/ram.scala 96:18]
  wire  ram_MPORT_1_en; // @[playground/src/ram/ram.scala 96:18]
  wire [5:0] ram_MPORT_1_addr; // @[playground/src/ram/ram.scala 96:18]
  wire [127:0] ram_MPORT_1_data; // @[playground/src/ram/ram.scala 96:18]
  wire  ram_output_MPORT_en; // @[playground/src/ram/ram.scala 96:18]
  wire [5:0] ram_output_MPORT_addr; // @[playground/src/ram/ram.scala 96:18]
  wire [127:0] ram_output_MPORT_data; // @[playground/src/ram/ram.scala 96:18]
  wire [127:0] ram_MPORT_data; // @[playground/src/ram/ram.scala 96:18]
  wire [5:0] ram_MPORT_addr; // @[playground/src/ram/ram.scala 96:18]
  wire  ram_MPORT_mask; // @[playground/src/ram/ram.scala 96:18]
  wire  ram_MPORT_en; // @[playground/src/ram/ram.scala 96:18]
  reg [127:0] output_; // @[playground/src/ram/ram.scala 97:25]
  wire  _T = ~io_CEN; // @[playground/src/ram/ram.scala 98:10]
  wire  _T_1 = ~io_WEN; // @[playground/src/ram/ram.scala 98:21]
  wire  _T_2 = ~io_CEN & ~io_WEN; // @[playground/src/ram/ram.scala 98:18]
  wire [127:0] _T_3 = ~io_BWEN; // @[playground/src/ram/ram.scala 99:30]
  wire [127:0] _T_4 = io_D & _T_3; // @[playground/src/ram/ram.scala 99:28]
  wire [127:0] _T_5 = ram_MPORT_1_data & io_BWEN; // @[playground/src/ram/ram.scala 99:53]
  assign ram_MPORT_1_en = _T & _T_1;
  assign ram_MPORT_1_addr = io_A;
  assign ram_MPORT_1_data = ram[ram_MPORT_1_addr]; // @[playground/src/ram/ram.scala 96:18]
  assign ram_output_MPORT_en = _T_2 ? 1'h0 : 1'h1;
  assign ram_output_MPORT_addr = io_A;
  assign ram_output_MPORT_data = ram[ram_output_MPORT_addr]; // @[playground/src/ram/ram.scala 96:18]
  assign ram_MPORT_data = _T_4 | _T_5;
  assign ram_MPORT_addr = io_A;
  assign ram_MPORT_mask = 1'h1;
  assign ram_MPORT_en = _T & _T_1;
  assign io_Q = output_; // @[playground/src/ram/ram.scala 104:10]
  always @(posedge clock) begin
    if (ram_MPORT_en & ram_MPORT_mask) begin
      ram[ram_MPORT_addr] <= ram_MPORT_data; // @[playground/src/ram/ram.scala 96:18]
    end
    if (reset) begin // @[playground/src/ram/ram.scala 97:25]
      output_ <= 128'h0; // @[playground/src/ram/ram.scala 97:25]
    end else if (~io_CEN & ~io_WEN) begin // @[playground/src/ram/ram.scala 98:30]
      output_ <= 128'h0; // @[playground/src/ram/ram.scala 100:16]
    end else begin
      output_ <= ram_output_MPORT_data; // @[playground/src/ram/ram.scala 102:16]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {4{`RANDOM}};
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    ram[initvar] = _RAND_0[127:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {4{`RANDOM}};
  output_ = _RAND_1[127:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Ram_bw(
  input          clock,
  input          reset,
  input          io_cen, // @[playground/src/ram/ram.scala 50:16]
  input          io_wen, // @[playground/src/ram/ram.scala 50:16]
  input  [5:0]   io_addr, // @[playground/src/ram/ram.scala 50:16]
  output [127:0] io_rdata, // @[playground/src/ram/ram.scala 50:16]
  input  [127:0] io_wdata, // @[playground/src/ram/ram.scala 50:16]
  input  [127:0] io_mask // @[playground/src/ram/ram.scala 50:16]
);
  wire  ram_clock; // @[playground/src/ram/ram.scala 51:21]
  wire  ram_reset; // @[playground/src/ram/ram.scala 51:21]
  wire [127:0] ram_io_Q; // @[playground/src/ram/ram.scala 51:21]
  wire  ram_io_CEN; // @[playground/src/ram/ram.scala 51:21]
  wire  ram_io_WEN; // @[playground/src/ram/ram.scala 51:21]
  wire [127:0] ram_io_BWEN; // @[playground/src/ram/ram.scala 51:21]
  wire [5:0] ram_io_A; // @[playground/src/ram/ram.scala 51:21]
  wire [127:0] ram_io_D; // @[playground/src/ram/ram.scala 51:21]
  S011HD1P_X32Y2D128_BW ram ( // @[playground/src/ram/ram.scala 51:21]
    .clock(ram_clock),
    .reset(ram_reset),
    .io_Q(ram_io_Q),
    .io_CEN(ram_io_CEN),
    .io_WEN(ram_io_WEN),
    .io_BWEN(ram_io_BWEN),
    .io_A(ram_io_A),
    .io_D(ram_io_D)
  );
  assign io_rdata = ram_io_Q; // @[playground/src/ram/ram.scala 52:14]
  assign ram_clock = clock;
  assign ram_reset = reset;
  assign ram_io_CEN = ~io_cen; // @[playground/src/ram/ram.scala 54:19]
  assign ram_io_WEN = ~io_wen; // @[playground/src/ram/ram.scala 55:19]
  assign ram_io_BWEN = ~io_mask; // @[playground/src/ram/ram.scala 58:20]
  assign ram_io_A = io_addr; // @[playground/src/ram/ram.scala 56:14]
  assign ram_io_D = io_wdata; // @[playground/src/ram/ram.scala 57:14]
endmodule
module MaxPeriodFibonacciLFSR(
  input   clock,
  input   reset,
  output  io_out_0, // @[src/main/scala/chisel3/util/random/PRNG.scala 42:22]
  output  io_out_1 // @[src/main/scala/chisel3/util/random/PRNG.scala 42:22]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  state_0; // @[src/main/scala/chisel3/util/random/PRNG.scala 55:49]
  reg  state_1; // @[src/main/scala/chisel3/util/random/PRNG.scala 55:49]
  wire  _T = state_1 ^ state_0; // @[src/main/scala/chisel3/util/random/LFSR.scala 15:41]
  assign io_out_0 = state_0; // @[src/main/scala/chisel3/util/random/PRNG.scala 78:10]
  assign io_out_1 = state_1; // @[src/main/scala/chisel3/util/random/PRNG.scala 78:10]
  always @(posedge clock) begin
    state_0 <= reset | _T; // @[src/main/scala/chisel3/util/random/PRNG.scala 55:{49,49}]
    if (reset) begin // @[src/main/scala/chisel3/util/random/PRNG.scala 55:49]
      state_1 <= 1'h0; // @[src/main/scala/chisel3/util/random/PRNG.scala 55:49]
    end else begin
      state_1 <= state_0;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state_0 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  state_1 = _RAND_1[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module InstCache(
  input         clock,
  input         reset,
  input         io_instAxi_ra_ready, // @[playground/src/noop/icache.scala 59:16]
  output        io_instAxi_ra_valid, // @[playground/src/noop/icache.scala 59:16]
  output [31:0] io_instAxi_ra_bits_addr, // @[playground/src/noop/icache.scala 59:16]
  input         io_instAxi_rd_valid, // @[playground/src/noop/icache.scala 59:16]
  input  [63:0] io_instAxi_rd_bits_data, // @[playground/src/noop/icache.scala 59:16]
  input         io_instAxi_rd_bits_last, // @[playground/src/noop/icache.scala 59:16]
  input  [31:0] io_icRead_addr, // @[playground/src/noop/icache.scala 59:16]
  output [63:0] io_icRead_inst, // @[playground/src/noop/icache.scala 59:16]
  input         io_icRead_arvalid, // @[playground/src/noop/icache.scala 59:16]
  output        io_icRead_ready, // @[playground/src/noop/icache.scala 59:16]
  output        io_icRead_rvalid, // @[playground/src/noop/icache.scala 59:16]
  input         io_flush // @[playground/src/noop/icache.scala 59:16]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [63:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
`endif // RANDOMIZE_REG_INIT
  wire  Ram_bw_clock; // @[playground/src/noop/icache.scala 67:57]
  wire  Ram_bw_reset; // @[playground/src/noop/icache.scala 67:57]
  wire  Ram_bw_io_cen; // @[playground/src/noop/icache.scala 67:57]
  wire  Ram_bw_io_wen; // @[playground/src/noop/icache.scala 67:57]
  wire [5:0] Ram_bw_io_addr; // @[playground/src/noop/icache.scala 67:57]
  wire [127:0] Ram_bw_io_rdata; // @[playground/src/noop/icache.scala 67:57]
  wire [127:0] Ram_bw_io_wdata; // @[playground/src/noop/icache.scala 67:57]
  wire [127:0] Ram_bw_io_mask; // @[playground/src/noop/icache.scala 67:57]
  wire  Ram_bw_1_clock; // @[playground/src/noop/icache.scala 67:57]
  wire  Ram_bw_1_reset; // @[playground/src/noop/icache.scala 67:57]
  wire  Ram_bw_1_io_cen; // @[playground/src/noop/icache.scala 67:57]
  wire  Ram_bw_1_io_wen; // @[playground/src/noop/icache.scala 67:57]
  wire [5:0] Ram_bw_1_io_addr; // @[playground/src/noop/icache.scala 67:57]
  wire [127:0] Ram_bw_1_io_rdata; // @[playground/src/noop/icache.scala 67:57]
  wire [127:0] Ram_bw_1_io_wdata; // @[playground/src/noop/icache.scala 67:57]
  wire [127:0] Ram_bw_1_io_mask; // @[playground/src/noop/icache.scala 67:57]
  wire  Ram_bw_2_clock; // @[playground/src/noop/icache.scala 67:57]
  wire  Ram_bw_2_reset; // @[playground/src/noop/icache.scala 67:57]
  wire  Ram_bw_2_io_cen; // @[playground/src/noop/icache.scala 67:57]
  wire  Ram_bw_2_io_wen; // @[playground/src/noop/icache.scala 67:57]
  wire [5:0] Ram_bw_2_io_addr; // @[playground/src/noop/icache.scala 67:57]
  wire [127:0] Ram_bw_2_io_rdata; // @[playground/src/noop/icache.scala 67:57]
  wire [127:0] Ram_bw_2_io_wdata; // @[playground/src/noop/icache.scala 67:57]
  wire [127:0] Ram_bw_2_io_mask; // @[playground/src/noop/icache.scala 67:57]
  wire  Ram_bw_3_clock; // @[playground/src/noop/icache.scala 67:57]
  wire  Ram_bw_3_reset; // @[playground/src/noop/icache.scala 67:57]
  wire  Ram_bw_3_io_cen; // @[playground/src/noop/icache.scala 67:57]
  wire  Ram_bw_3_io_wen; // @[playground/src/noop/icache.scala 67:57]
  wire [5:0] Ram_bw_3_io_addr; // @[playground/src/noop/icache.scala 67:57]
  wire [127:0] Ram_bw_3_io_rdata; // @[playground/src/noop/icache.scala 67:57]
  wire [127:0] Ram_bw_3_io_wdata; // @[playground/src/noop/icache.scala 67:57]
  wire [127:0] Ram_bw_3_io_mask; // @[playground/src/noop/icache.scala 67:57]
  wire  matchWay_prng_clock; // @[src/main/scala/chisel3/util/random/PRNG.scala 91:22]
  wire  matchWay_prng_reset; // @[src/main/scala/chisel3/util/random/PRNG.scala 91:22]
  wire  matchWay_prng_io_out_0; // @[src/main/scala/chisel3/util/random/PRNG.scala 91:22]
  wire  matchWay_prng_io_out_1; // @[src/main/scala/chisel3/util/random/PRNG.scala 91:22]
  reg [21:0] tag_0_0; // @[playground/src/noop/icache.scala 65:26]
  reg [21:0] tag_0_1; // @[playground/src/noop/icache.scala 65:26]
  reg [21:0] tag_0_2; // @[playground/src/noop/icache.scala 65:26]
  reg [21:0] tag_0_3; // @[playground/src/noop/icache.scala 65:26]
  reg [21:0] tag_0_4; // @[playground/src/noop/icache.scala 65:26]
  reg [21:0] tag_0_5; // @[playground/src/noop/icache.scala 65:26]
  reg [21:0] tag_0_6; // @[playground/src/noop/icache.scala 65:26]
  reg [21:0] tag_0_7; // @[playground/src/noop/icache.scala 65:26]
  reg [21:0] tag_0_8; // @[playground/src/noop/icache.scala 65:26]
  reg [21:0] tag_0_9; // @[playground/src/noop/icache.scala 65:26]
  reg [21:0] tag_0_10; // @[playground/src/noop/icache.scala 65:26]
  reg [21:0] tag_0_11; // @[playground/src/noop/icache.scala 65:26]
  reg [21:0] tag_0_12; // @[playground/src/noop/icache.scala 65:26]
  reg [21:0] tag_0_13; // @[playground/src/noop/icache.scala 65:26]
  reg [21:0] tag_0_14; // @[playground/src/noop/icache.scala 65:26]
  reg [21:0] tag_0_15; // @[playground/src/noop/icache.scala 65:26]
  reg [21:0] tag_1_0; // @[playground/src/noop/icache.scala 65:26]
  reg [21:0] tag_1_1; // @[playground/src/noop/icache.scala 65:26]
  reg [21:0] tag_1_2; // @[playground/src/noop/icache.scala 65:26]
  reg [21:0] tag_1_3; // @[playground/src/noop/icache.scala 65:26]
  reg [21:0] tag_1_4; // @[playground/src/noop/icache.scala 65:26]
  reg [21:0] tag_1_5; // @[playground/src/noop/icache.scala 65:26]
  reg [21:0] tag_1_6; // @[playground/src/noop/icache.scala 65:26]
  reg [21:0] tag_1_7; // @[playground/src/noop/icache.scala 65:26]
  reg [21:0] tag_1_8; // @[playground/src/noop/icache.scala 65:26]
  reg [21:0] tag_1_9; // @[playground/src/noop/icache.scala 65:26]
  reg [21:0] tag_1_10; // @[playground/src/noop/icache.scala 65:26]
  reg [21:0] tag_1_11; // @[playground/src/noop/icache.scala 65:26]
  reg [21:0] tag_1_12; // @[playground/src/noop/icache.scala 65:26]
  reg [21:0] tag_1_13; // @[playground/src/noop/icache.scala 65:26]
  reg [21:0] tag_1_14; // @[playground/src/noop/icache.scala 65:26]
  reg [21:0] tag_1_15; // @[playground/src/noop/icache.scala 65:26]
  reg [21:0] tag_2_0; // @[playground/src/noop/icache.scala 65:26]
  reg [21:0] tag_2_1; // @[playground/src/noop/icache.scala 65:26]
  reg [21:0] tag_2_2; // @[playground/src/noop/icache.scala 65:26]
  reg [21:0] tag_2_3; // @[playground/src/noop/icache.scala 65:26]
  reg [21:0] tag_2_4; // @[playground/src/noop/icache.scala 65:26]
  reg [21:0] tag_2_5; // @[playground/src/noop/icache.scala 65:26]
  reg [21:0] tag_2_6; // @[playground/src/noop/icache.scala 65:26]
  reg [21:0] tag_2_7; // @[playground/src/noop/icache.scala 65:26]
  reg [21:0] tag_2_8; // @[playground/src/noop/icache.scala 65:26]
  reg [21:0] tag_2_9; // @[playground/src/noop/icache.scala 65:26]
  reg [21:0] tag_2_10; // @[playground/src/noop/icache.scala 65:26]
  reg [21:0] tag_2_11; // @[playground/src/noop/icache.scala 65:26]
  reg [21:0] tag_2_12; // @[playground/src/noop/icache.scala 65:26]
  reg [21:0] tag_2_13; // @[playground/src/noop/icache.scala 65:26]
  reg [21:0] tag_2_14; // @[playground/src/noop/icache.scala 65:26]
  reg [21:0] tag_2_15; // @[playground/src/noop/icache.scala 65:26]
  reg [21:0] tag_3_0; // @[playground/src/noop/icache.scala 65:26]
  reg [21:0] tag_3_1; // @[playground/src/noop/icache.scala 65:26]
  reg [21:0] tag_3_2; // @[playground/src/noop/icache.scala 65:26]
  reg [21:0] tag_3_3; // @[playground/src/noop/icache.scala 65:26]
  reg [21:0] tag_3_4; // @[playground/src/noop/icache.scala 65:26]
  reg [21:0] tag_3_5; // @[playground/src/noop/icache.scala 65:26]
  reg [21:0] tag_3_6; // @[playground/src/noop/icache.scala 65:26]
  reg [21:0] tag_3_7; // @[playground/src/noop/icache.scala 65:26]
  reg [21:0] tag_3_8; // @[playground/src/noop/icache.scala 65:26]
  reg [21:0] tag_3_9; // @[playground/src/noop/icache.scala 65:26]
  reg [21:0] tag_3_10; // @[playground/src/noop/icache.scala 65:26]
  reg [21:0] tag_3_11; // @[playground/src/noop/icache.scala 65:26]
  reg [21:0] tag_3_12; // @[playground/src/noop/icache.scala 65:26]
  reg [21:0] tag_3_13; // @[playground/src/noop/icache.scala 65:26]
  reg [21:0] tag_3_14; // @[playground/src/noop/icache.scala 65:26]
  reg [21:0] tag_3_15; // @[playground/src/noop/icache.scala 65:26]
  reg  valid_0_0; // @[playground/src/noop/icache.scala 66:26]
  reg  valid_0_1; // @[playground/src/noop/icache.scala 66:26]
  reg  valid_0_2; // @[playground/src/noop/icache.scala 66:26]
  reg  valid_0_3; // @[playground/src/noop/icache.scala 66:26]
  reg  valid_0_4; // @[playground/src/noop/icache.scala 66:26]
  reg  valid_0_5; // @[playground/src/noop/icache.scala 66:26]
  reg  valid_0_6; // @[playground/src/noop/icache.scala 66:26]
  reg  valid_0_7; // @[playground/src/noop/icache.scala 66:26]
  reg  valid_0_8; // @[playground/src/noop/icache.scala 66:26]
  reg  valid_0_9; // @[playground/src/noop/icache.scala 66:26]
  reg  valid_0_10; // @[playground/src/noop/icache.scala 66:26]
  reg  valid_0_11; // @[playground/src/noop/icache.scala 66:26]
  reg  valid_0_12; // @[playground/src/noop/icache.scala 66:26]
  reg  valid_0_13; // @[playground/src/noop/icache.scala 66:26]
  reg  valid_0_14; // @[playground/src/noop/icache.scala 66:26]
  reg  valid_0_15; // @[playground/src/noop/icache.scala 66:26]
  reg  valid_1_0; // @[playground/src/noop/icache.scala 66:26]
  reg  valid_1_1; // @[playground/src/noop/icache.scala 66:26]
  reg  valid_1_2; // @[playground/src/noop/icache.scala 66:26]
  reg  valid_1_3; // @[playground/src/noop/icache.scala 66:26]
  reg  valid_1_4; // @[playground/src/noop/icache.scala 66:26]
  reg  valid_1_5; // @[playground/src/noop/icache.scala 66:26]
  reg  valid_1_6; // @[playground/src/noop/icache.scala 66:26]
  reg  valid_1_7; // @[playground/src/noop/icache.scala 66:26]
  reg  valid_1_8; // @[playground/src/noop/icache.scala 66:26]
  reg  valid_1_9; // @[playground/src/noop/icache.scala 66:26]
  reg  valid_1_10; // @[playground/src/noop/icache.scala 66:26]
  reg  valid_1_11; // @[playground/src/noop/icache.scala 66:26]
  reg  valid_1_12; // @[playground/src/noop/icache.scala 66:26]
  reg  valid_1_13; // @[playground/src/noop/icache.scala 66:26]
  reg  valid_1_14; // @[playground/src/noop/icache.scala 66:26]
  reg  valid_1_15; // @[playground/src/noop/icache.scala 66:26]
  reg  valid_2_0; // @[playground/src/noop/icache.scala 66:26]
  reg  valid_2_1; // @[playground/src/noop/icache.scala 66:26]
  reg  valid_2_2; // @[playground/src/noop/icache.scala 66:26]
  reg  valid_2_3; // @[playground/src/noop/icache.scala 66:26]
  reg  valid_2_4; // @[playground/src/noop/icache.scala 66:26]
  reg  valid_2_5; // @[playground/src/noop/icache.scala 66:26]
  reg  valid_2_6; // @[playground/src/noop/icache.scala 66:26]
  reg  valid_2_7; // @[playground/src/noop/icache.scala 66:26]
  reg  valid_2_8; // @[playground/src/noop/icache.scala 66:26]
  reg  valid_2_9; // @[playground/src/noop/icache.scala 66:26]
  reg  valid_2_10; // @[playground/src/noop/icache.scala 66:26]
  reg  valid_2_11; // @[playground/src/noop/icache.scala 66:26]
  reg  valid_2_12; // @[playground/src/noop/icache.scala 66:26]
  reg  valid_2_13; // @[playground/src/noop/icache.scala 66:26]
  reg  valid_2_14; // @[playground/src/noop/icache.scala 66:26]
  reg  valid_2_15; // @[playground/src/noop/icache.scala 66:26]
  reg  valid_3_0; // @[playground/src/noop/icache.scala 66:26]
  reg  valid_3_1; // @[playground/src/noop/icache.scala 66:26]
  reg  valid_3_2; // @[playground/src/noop/icache.scala 66:26]
  reg  valid_3_3; // @[playground/src/noop/icache.scala 66:26]
  reg  valid_3_4; // @[playground/src/noop/icache.scala 66:26]
  reg  valid_3_5; // @[playground/src/noop/icache.scala 66:26]
  reg  valid_3_6; // @[playground/src/noop/icache.scala 66:26]
  reg  valid_3_7; // @[playground/src/noop/icache.scala 66:26]
  reg  valid_3_8; // @[playground/src/noop/icache.scala 66:26]
  reg  valid_3_9; // @[playground/src/noop/icache.scala 66:26]
  reg  valid_3_10; // @[playground/src/noop/icache.scala 66:26]
  reg  valid_3_11; // @[playground/src/noop/icache.scala 66:26]
  reg  valid_3_12; // @[playground/src/noop/icache.scala 66:26]
  reg  valid_3_13; // @[playground/src/noop/icache.scala 66:26]
  reg  valid_3_14; // @[playground/src/noop/icache.scala 66:26]
  reg  valid_3_15; // @[playground/src/noop/icache.scala 66:26]
  reg  wait_r; // @[playground/src/noop/icache.scala 71:30]
  reg  valid_r; // @[playground/src/noop/icache.scala 72:30]
  wire  valid_in = io_icRead_arvalid & ~io_flush; // @[playground/src/noop/icache.scala 74:41]
  wire  hs_in = io_icRead_ready & io_icRead_arvalid; // @[playground/src/noop/icache.scala 75:39]
  wire  _io_icRead_ready_T = ~wait_r; // @[playground/src/noop/icache.scala 76:40]
  reg [31:0] addr_r; // @[playground/src/noop/icache.scala 78:34]
  reg [31:0] matchWay_r; // @[playground/src/noop/icache.scala 79:34]
  reg [2:0] axiOffset; // @[playground/src/noop/icache.scala 80:34]
  reg [63:0] databuf; // @[playground/src/noop/icache.scala 81:34]
  wire [31:0] cur_addr = hs_in ? io_icRead_addr : addr_r; // @[playground/src/noop/icache.scala 82:30]
  wire [21:0] instTag = cur_addr[31:10]; // @[playground/src/noop/icache.scala 83:35]
  wire [3:0] blockIdx = cur_addr[9:6]; // @[playground/src/noop/icache.scala 84:35]
  wire [5:0] cur_ram_addr = cur_addr[9:4]; // @[playground/src/noop/icache.scala 85:35]
  wire [5:0] cur_raddr = {blockIdx,axiOffset[2:1]}; // @[playground/src/noop/icache.scala 86:30]
  wire [21:0] _GEN_1 = 4'h1 == blockIdx ? tag_0_1 : tag_0_0; // @[playground/src/noop/icache.scala 87:{85,85}]
  wire [21:0] _GEN_2 = 4'h2 == blockIdx ? tag_0_2 : _GEN_1; // @[playground/src/noop/icache.scala 87:{85,85}]
  wire [21:0] _GEN_3 = 4'h3 == blockIdx ? tag_0_3 : _GEN_2; // @[playground/src/noop/icache.scala 87:{85,85}]
  wire [21:0] _GEN_4 = 4'h4 == blockIdx ? tag_0_4 : _GEN_3; // @[playground/src/noop/icache.scala 87:{85,85}]
  wire [21:0] _GEN_5 = 4'h5 == blockIdx ? tag_0_5 : _GEN_4; // @[playground/src/noop/icache.scala 87:{85,85}]
  wire [21:0] _GEN_6 = 4'h6 == blockIdx ? tag_0_6 : _GEN_5; // @[playground/src/noop/icache.scala 87:{85,85}]
  wire [21:0] _GEN_7 = 4'h7 == blockIdx ? tag_0_7 : _GEN_6; // @[playground/src/noop/icache.scala 87:{85,85}]
  wire [21:0] _GEN_8 = 4'h8 == blockIdx ? tag_0_8 : _GEN_7; // @[playground/src/noop/icache.scala 87:{85,85}]
  wire [21:0] _GEN_9 = 4'h9 == blockIdx ? tag_0_9 : _GEN_8; // @[playground/src/noop/icache.scala 87:{85,85}]
  wire [21:0] _GEN_10 = 4'ha == blockIdx ? tag_0_10 : _GEN_9; // @[playground/src/noop/icache.scala 87:{85,85}]
  wire [21:0] _GEN_11 = 4'hb == blockIdx ? tag_0_11 : _GEN_10; // @[playground/src/noop/icache.scala 87:{85,85}]
  wire [21:0] _GEN_12 = 4'hc == blockIdx ? tag_0_12 : _GEN_11; // @[playground/src/noop/icache.scala 87:{85,85}]
  wire [21:0] _GEN_13 = 4'hd == blockIdx ? tag_0_13 : _GEN_12; // @[playground/src/noop/icache.scala 87:{85,85}]
  wire [21:0] _GEN_14 = 4'he == blockIdx ? tag_0_14 : _GEN_13; // @[playground/src/noop/icache.scala 87:{85,85}]
  wire [21:0] _GEN_15 = 4'hf == blockIdx ? tag_0_15 : _GEN_14; // @[playground/src/noop/icache.scala 87:{85,85}]
  wire  _GEN_17 = 4'h1 == blockIdx ? valid_0_1 : valid_0_0; // @[playground/src/noop/icache.scala 87:{97,97}]
  wire  _GEN_18 = 4'h2 == blockIdx ? valid_0_2 : _GEN_17; // @[playground/src/noop/icache.scala 87:{97,97}]
  wire  _GEN_19 = 4'h3 == blockIdx ? valid_0_3 : _GEN_18; // @[playground/src/noop/icache.scala 87:{97,97}]
  wire  _GEN_20 = 4'h4 == blockIdx ? valid_0_4 : _GEN_19; // @[playground/src/noop/icache.scala 87:{97,97}]
  wire  _GEN_21 = 4'h5 == blockIdx ? valid_0_5 : _GEN_20; // @[playground/src/noop/icache.scala 87:{97,97}]
  wire  _GEN_22 = 4'h6 == blockIdx ? valid_0_6 : _GEN_21; // @[playground/src/noop/icache.scala 87:{97,97}]
  wire  _GEN_23 = 4'h7 == blockIdx ? valid_0_7 : _GEN_22; // @[playground/src/noop/icache.scala 87:{97,97}]
  wire  _GEN_24 = 4'h8 == blockIdx ? valid_0_8 : _GEN_23; // @[playground/src/noop/icache.scala 87:{97,97}]
  wire  _GEN_25 = 4'h9 == blockIdx ? valid_0_9 : _GEN_24; // @[playground/src/noop/icache.scala 87:{97,97}]
  wire  _GEN_26 = 4'ha == blockIdx ? valid_0_10 : _GEN_25; // @[playground/src/noop/icache.scala 87:{97,97}]
  wire  _GEN_27 = 4'hb == blockIdx ? valid_0_11 : _GEN_26; // @[playground/src/noop/icache.scala 87:{97,97}]
  wire  _GEN_28 = 4'hc == blockIdx ? valid_0_12 : _GEN_27; // @[playground/src/noop/icache.scala 87:{97,97}]
  wire  _GEN_29 = 4'hd == blockIdx ? valid_0_13 : _GEN_28; // @[playground/src/noop/icache.scala 87:{97,97}]
  wire  _GEN_30 = 4'he == blockIdx ? valid_0_14 : _GEN_29; // @[playground/src/noop/icache.scala 87:{97,97}]
  wire  _GEN_31 = 4'hf == blockIdx ? valid_0_15 : _GEN_30; // @[playground/src/noop/icache.scala 87:{97,97}]
  wire  cache_hit_vec_0 = _GEN_15 == instTag & _GEN_31; // @[playground/src/noop/icache.scala 87:97]
  wire [21:0] _GEN_33 = 4'h1 == blockIdx ? tag_1_1 : tag_1_0; // @[playground/src/noop/icache.scala 87:{85,85}]
  wire [21:0] _GEN_34 = 4'h2 == blockIdx ? tag_1_2 : _GEN_33; // @[playground/src/noop/icache.scala 87:{85,85}]
  wire [21:0] _GEN_35 = 4'h3 == blockIdx ? tag_1_3 : _GEN_34; // @[playground/src/noop/icache.scala 87:{85,85}]
  wire [21:0] _GEN_36 = 4'h4 == blockIdx ? tag_1_4 : _GEN_35; // @[playground/src/noop/icache.scala 87:{85,85}]
  wire [21:0] _GEN_37 = 4'h5 == blockIdx ? tag_1_5 : _GEN_36; // @[playground/src/noop/icache.scala 87:{85,85}]
  wire [21:0] _GEN_38 = 4'h6 == blockIdx ? tag_1_6 : _GEN_37; // @[playground/src/noop/icache.scala 87:{85,85}]
  wire [21:0] _GEN_39 = 4'h7 == blockIdx ? tag_1_7 : _GEN_38; // @[playground/src/noop/icache.scala 87:{85,85}]
  wire [21:0] _GEN_40 = 4'h8 == blockIdx ? tag_1_8 : _GEN_39; // @[playground/src/noop/icache.scala 87:{85,85}]
  wire [21:0] _GEN_41 = 4'h9 == blockIdx ? tag_1_9 : _GEN_40; // @[playground/src/noop/icache.scala 87:{85,85}]
  wire [21:0] _GEN_42 = 4'ha == blockIdx ? tag_1_10 : _GEN_41; // @[playground/src/noop/icache.scala 87:{85,85}]
  wire [21:0] _GEN_43 = 4'hb == blockIdx ? tag_1_11 : _GEN_42; // @[playground/src/noop/icache.scala 87:{85,85}]
  wire [21:0] _GEN_44 = 4'hc == blockIdx ? tag_1_12 : _GEN_43; // @[playground/src/noop/icache.scala 87:{85,85}]
  wire [21:0] _GEN_45 = 4'hd == blockIdx ? tag_1_13 : _GEN_44; // @[playground/src/noop/icache.scala 87:{85,85}]
  wire [21:0] _GEN_46 = 4'he == blockIdx ? tag_1_14 : _GEN_45; // @[playground/src/noop/icache.scala 87:{85,85}]
  wire [21:0] _GEN_47 = 4'hf == blockIdx ? tag_1_15 : _GEN_46; // @[playground/src/noop/icache.scala 87:{85,85}]
  wire  _GEN_49 = 4'h1 == blockIdx ? valid_1_1 : valid_1_0; // @[playground/src/noop/icache.scala 87:{97,97}]
  wire  _GEN_50 = 4'h2 == blockIdx ? valid_1_2 : _GEN_49; // @[playground/src/noop/icache.scala 87:{97,97}]
  wire  _GEN_51 = 4'h3 == blockIdx ? valid_1_3 : _GEN_50; // @[playground/src/noop/icache.scala 87:{97,97}]
  wire  _GEN_52 = 4'h4 == blockIdx ? valid_1_4 : _GEN_51; // @[playground/src/noop/icache.scala 87:{97,97}]
  wire  _GEN_53 = 4'h5 == blockIdx ? valid_1_5 : _GEN_52; // @[playground/src/noop/icache.scala 87:{97,97}]
  wire  _GEN_54 = 4'h6 == blockIdx ? valid_1_6 : _GEN_53; // @[playground/src/noop/icache.scala 87:{97,97}]
  wire  _GEN_55 = 4'h7 == blockIdx ? valid_1_7 : _GEN_54; // @[playground/src/noop/icache.scala 87:{97,97}]
  wire  _GEN_56 = 4'h8 == blockIdx ? valid_1_8 : _GEN_55; // @[playground/src/noop/icache.scala 87:{97,97}]
  wire  _GEN_57 = 4'h9 == blockIdx ? valid_1_9 : _GEN_56; // @[playground/src/noop/icache.scala 87:{97,97}]
  wire  _GEN_58 = 4'ha == blockIdx ? valid_1_10 : _GEN_57; // @[playground/src/noop/icache.scala 87:{97,97}]
  wire  _GEN_59 = 4'hb == blockIdx ? valid_1_11 : _GEN_58; // @[playground/src/noop/icache.scala 87:{97,97}]
  wire  _GEN_60 = 4'hc == blockIdx ? valid_1_12 : _GEN_59; // @[playground/src/noop/icache.scala 87:{97,97}]
  wire  _GEN_61 = 4'hd == blockIdx ? valid_1_13 : _GEN_60; // @[playground/src/noop/icache.scala 87:{97,97}]
  wire  _GEN_62 = 4'he == blockIdx ? valid_1_14 : _GEN_61; // @[playground/src/noop/icache.scala 87:{97,97}]
  wire  _GEN_63 = 4'hf == blockIdx ? valid_1_15 : _GEN_62; // @[playground/src/noop/icache.scala 87:{97,97}]
  wire  cache_hit_vec_1 = _GEN_47 == instTag & _GEN_63; // @[playground/src/noop/icache.scala 87:97]
  wire [21:0] _GEN_65 = 4'h1 == blockIdx ? tag_2_1 : tag_2_0; // @[playground/src/noop/icache.scala 87:{85,85}]
  wire [21:0] _GEN_66 = 4'h2 == blockIdx ? tag_2_2 : _GEN_65; // @[playground/src/noop/icache.scala 87:{85,85}]
  wire [21:0] _GEN_67 = 4'h3 == blockIdx ? tag_2_3 : _GEN_66; // @[playground/src/noop/icache.scala 87:{85,85}]
  wire [21:0] _GEN_68 = 4'h4 == blockIdx ? tag_2_4 : _GEN_67; // @[playground/src/noop/icache.scala 87:{85,85}]
  wire [21:0] _GEN_69 = 4'h5 == blockIdx ? tag_2_5 : _GEN_68; // @[playground/src/noop/icache.scala 87:{85,85}]
  wire [21:0] _GEN_70 = 4'h6 == blockIdx ? tag_2_6 : _GEN_69; // @[playground/src/noop/icache.scala 87:{85,85}]
  wire [21:0] _GEN_71 = 4'h7 == blockIdx ? tag_2_7 : _GEN_70; // @[playground/src/noop/icache.scala 87:{85,85}]
  wire [21:0] _GEN_72 = 4'h8 == blockIdx ? tag_2_8 : _GEN_71; // @[playground/src/noop/icache.scala 87:{85,85}]
  wire [21:0] _GEN_73 = 4'h9 == blockIdx ? tag_2_9 : _GEN_72; // @[playground/src/noop/icache.scala 87:{85,85}]
  wire [21:0] _GEN_74 = 4'ha == blockIdx ? tag_2_10 : _GEN_73; // @[playground/src/noop/icache.scala 87:{85,85}]
  wire [21:0] _GEN_75 = 4'hb == blockIdx ? tag_2_11 : _GEN_74; // @[playground/src/noop/icache.scala 87:{85,85}]
  wire [21:0] _GEN_76 = 4'hc == blockIdx ? tag_2_12 : _GEN_75; // @[playground/src/noop/icache.scala 87:{85,85}]
  wire [21:0] _GEN_77 = 4'hd == blockIdx ? tag_2_13 : _GEN_76; // @[playground/src/noop/icache.scala 87:{85,85}]
  wire [21:0] _GEN_78 = 4'he == blockIdx ? tag_2_14 : _GEN_77; // @[playground/src/noop/icache.scala 87:{85,85}]
  wire [21:0] _GEN_79 = 4'hf == blockIdx ? tag_2_15 : _GEN_78; // @[playground/src/noop/icache.scala 87:{85,85}]
  wire  _GEN_81 = 4'h1 == blockIdx ? valid_2_1 : valid_2_0; // @[playground/src/noop/icache.scala 87:{97,97}]
  wire  _GEN_82 = 4'h2 == blockIdx ? valid_2_2 : _GEN_81; // @[playground/src/noop/icache.scala 87:{97,97}]
  wire  _GEN_83 = 4'h3 == blockIdx ? valid_2_3 : _GEN_82; // @[playground/src/noop/icache.scala 87:{97,97}]
  wire  _GEN_84 = 4'h4 == blockIdx ? valid_2_4 : _GEN_83; // @[playground/src/noop/icache.scala 87:{97,97}]
  wire  _GEN_85 = 4'h5 == blockIdx ? valid_2_5 : _GEN_84; // @[playground/src/noop/icache.scala 87:{97,97}]
  wire  _GEN_86 = 4'h6 == blockIdx ? valid_2_6 : _GEN_85; // @[playground/src/noop/icache.scala 87:{97,97}]
  wire  _GEN_87 = 4'h7 == blockIdx ? valid_2_7 : _GEN_86; // @[playground/src/noop/icache.scala 87:{97,97}]
  wire  _GEN_88 = 4'h8 == blockIdx ? valid_2_8 : _GEN_87; // @[playground/src/noop/icache.scala 87:{97,97}]
  wire  _GEN_89 = 4'h9 == blockIdx ? valid_2_9 : _GEN_88; // @[playground/src/noop/icache.scala 87:{97,97}]
  wire  _GEN_90 = 4'ha == blockIdx ? valid_2_10 : _GEN_89; // @[playground/src/noop/icache.scala 87:{97,97}]
  wire  _GEN_91 = 4'hb == blockIdx ? valid_2_11 : _GEN_90; // @[playground/src/noop/icache.scala 87:{97,97}]
  wire  _GEN_92 = 4'hc == blockIdx ? valid_2_12 : _GEN_91; // @[playground/src/noop/icache.scala 87:{97,97}]
  wire  _GEN_93 = 4'hd == blockIdx ? valid_2_13 : _GEN_92; // @[playground/src/noop/icache.scala 87:{97,97}]
  wire  _GEN_94 = 4'he == blockIdx ? valid_2_14 : _GEN_93; // @[playground/src/noop/icache.scala 87:{97,97}]
  wire  _GEN_95 = 4'hf == blockIdx ? valid_2_15 : _GEN_94; // @[playground/src/noop/icache.scala 87:{97,97}]
  wire  cache_hit_vec_2 = _GEN_79 == instTag & _GEN_95; // @[playground/src/noop/icache.scala 87:97]
  wire [21:0] _GEN_97 = 4'h1 == blockIdx ? tag_3_1 : tag_3_0; // @[playground/src/noop/icache.scala 87:{85,85}]
  wire [21:0] _GEN_98 = 4'h2 == blockIdx ? tag_3_2 : _GEN_97; // @[playground/src/noop/icache.scala 87:{85,85}]
  wire [21:0] _GEN_99 = 4'h3 == blockIdx ? tag_3_3 : _GEN_98; // @[playground/src/noop/icache.scala 87:{85,85}]
  wire [21:0] _GEN_100 = 4'h4 == blockIdx ? tag_3_4 : _GEN_99; // @[playground/src/noop/icache.scala 87:{85,85}]
  wire [21:0] _GEN_101 = 4'h5 == blockIdx ? tag_3_5 : _GEN_100; // @[playground/src/noop/icache.scala 87:{85,85}]
  wire [21:0] _GEN_102 = 4'h6 == blockIdx ? tag_3_6 : _GEN_101; // @[playground/src/noop/icache.scala 87:{85,85}]
  wire [21:0] _GEN_103 = 4'h7 == blockIdx ? tag_3_7 : _GEN_102; // @[playground/src/noop/icache.scala 87:{85,85}]
  wire [21:0] _GEN_104 = 4'h8 == blockIdx ? tag_3_8 : _GEN_103; // @[playground/src/noop/icache.scala 87:{85,85}]
  wire [21:0] _GEN_105 = 4'h9 == blockIdx ? tag_3_9 : _GEN_104; // @[playground/src/noop/icache.scala 87:{85,85}]
  wire [21:0] _GEN_106 = 4'ha == blockIdx ? tag_3_10 : _GEN_105; // @[playground/src/noop/icache.scala 87:{85,85}]
  wire [21:0] _GEN_107 = 4'hb == blockIdx ? tag_3_11 : _GEN_106; // @[playground/src/noop/icache.scala 87:{85,85}]
  wire [21:0] _GEN_108 = 4'hc == blockIdx ? tag_3_12 : _GEN_107; // @[playground/src/noop/icache.scala 87:{85,85}]
  wire [21:0] _GEN_109 = 4'hd == blockIdx ? tag_3_13 : _GEN_108; // @[playground/src/noop/icache.scala 87:{85,85}]
  wire [21:0] _GEN_110 = 4'he == blockIdx ? tag_3_14 : _GEN_109; // @[playground/src/noop/icache.scala 87:{85,85}]
  wire [21:0] _GEN_111 = 4'hf == blockIdx ? tag_3_15 : _GEN_110; // @[playground/src/noop/icache.scala 87:{85,85}]
  wire  _GEN_113 = 4'h1 == blockIdx ? valid_3_1 : valid_3_0; // @[playground/src/noop/icache.scala 87:{97,97}]
  wire  _GEN_114 = 4'h2 == blockIdx ? valid_3_2 : _GEN_113; // @[playground/src/noop/icache.scala 87:{97,97}]
  wire  _GEN_115 = 4'h3 == blockIdx ? valid_3_3 : _GEN_114; // @[playground/src/noop/icache.scala 87:{97,97}]
  wire  _GEN_116 = 4'h4 == blockIdx ? valid_3_4 : _GEN_115; // @[playground/src/noop/icache.scala 87:{97,97}]
  wire  _GEN_117 = 4'h5 == blockIdx ? valid_3_5 : _GEN_116; // @[playground/src/noop/icache.scala 87:{97,97}]
  wire  _GEN_118 = 4'h6 == blockIdx ? valid_3_6 : _GEN_117; // @[playground/src/noop/icache.scala 87:{97,97}]
  wire  _GEN_119 = 4'h7 == blockIdx ? valid_3_7 : _GEN_118; // @[playground/src/noop/icache.scala 87:{97,97}]
  wire  _GEN_120 = 4'h8 == blockIdx ? valid_3_8 : _GEN_119; // @[playground/src/noop/icache.scala 87:{97,97}]
  wire  _GEN_121 = 4'h9 == blockIdx ? valid_3_9 : _GEN_120; // @[playground/src/noop/icache.scala 87:{97,97}]
  wire  _GEN_122 = 4'ha == blockIdx ? valid_3_10 : _GEN_121; // @[playground/src/noop/icache.scala 87:{97,97}]
  wire  _GEN_123 = 4'hb == blockIdx ? valid_3_11 : _GEN_122; // @[playground/src/noop/icache.scala 87:{97,97}]
  wire  _GEN_124 = 4'hc == blockIdx ? valid_3_12 : _GEN_123; // @[playground/src/noop/icache.scala 87:{97,97}]
  wire  _GEN_125 = 4'hd == blockIdx ? valid_3_13 : _GEN_124; // @[playground/src/noop/icache.scala 87:{97,97}]
  wire  _GEN_126 = 4'he == blockIdx ? valid_3_14 : _GEN_125; // @[playground/src/noop/icache.scala 87:{97,97}]
  wire  _GEN_127 = 4'hf == blockIdx ? valid_3_15 : _GEN_126; // @[playground/src/noop/icache.scala 87:{97,97}]
  wire  cache_hit_vec_3 = _GEN_111 == instTag & _GEN_127; // @[playground/src/noop/icache.scala 87:97]
  wire [3:0] _cacheHit_T = {cache_hit_vec_3,cache_hit_vec_2,cache_hit_vec_1,cache_hit_vec_0}; // @[playground/src/noop/icache.scala 88:41]
  wire  cacheHit = |_cacheHit_T; // @[playground/src/noop/icache.scala 88:48]
  wire [1:0] matchWay_hi_1 = _cacheHit_T[3:2]; // @[src/main/scala/chisel3/util/OneHot.scala 30:18]
  wire [1:0] matchWay_lo_1 = _cacheHit_T[1:0]; // @[src/main/scala/chisel3/util/OneHot.scala 31:18]
  wire [1:0] _matchWay_T_2 = matchWay_hi_1 | matchWay_lo_1; // @[src/main/scala/chisel3/util/OneHot.scala 32:28]
  wire [1:0] _matchWay_T_4 = {|matchWay_hi_1,_matchWay_T_2[1]}; // @[src/main/scala/chisel3/util/OneHot.scala 32:10]
  wire [1:0] _matchWay_T_5 = {matchWay_prng_io_out_1,matchWay_prng_io_out_0}; // @[src/main/scala/chisel3/util/random/PRNG.scala 95:17]
  wire [1:0] matchWay = cacheHit ? _matchWay_T_4 : _matchWay_T_5; // @[playground/src/noop/icache.scala 89:30]
  wire [31:0] cur_way = hs_in ? {{30'd0}, matchWay} : matchWay_r; // @[playground/src/noop/icache.scala 90:30]
  wire [3:0] pre_blockIdx = addr_r[9:6]; // @[playground/src/noop/icache.scala 91:33]
  wire [21:0] pre_instTag = addr_r[31:10]; // @[playground/src/noop/icache.scala 92:33]
  wire  _GEN_130 = io_flush ? 1'h0 : valid_0_0; // @[playground/src/noop/icache.scala 98:19 99:17 66:26]
  wire  _GEN_131 = io_flush ? 1'h0 : valid_0_1; // @[playground/src/noop/icache.scala 98:19 99:17 66:26]
  wire  _GEN_132 = io_flush ? 1'h0 : valid_0_2; // @[playground/src/noop/icache.scala 98:19 99:17 66:26]
  wire  _GEN_133 = io_flush ? 1'h0 : valid_0_3; // @[playground/src/noop/icache.scala 98:19 99:17 66:26]
  wire  _GEN_134 = io_flush ? 1'h0 : valid_0_4; // @[playground/src/noop/icache.scala 98:19 99:17 66:26]
  wire  _GEN_135 = io_flush ? 1'h0 : valid_0_5; // @[playground/src/noop/icache.scala 98:19 99:17 66:26]
  wire  _GEN_136 = io_flush ? 1'h0 : valid_0_6; // @[playground/src/noop/icache.scala 98:19 99:17 66:26]
  wire  _GEN_137 = io_flush ? 1'h0 : valid_0_7; // @[playground/src/noop/icache.scala 98:19 99:17 66:26]
  wire  _GEN_138 = io_flush ? 1'h0 : valid_0_8; // @[playground/src/noop/icache.scala 98:19 99:17 66:26]
  wire  _GEN_139 = io_flush ? 1'h0 : valid_0_9; // @[playground/src/noop/icache.scala 98:19 99:17 66:26]
  wire  _GEN_140 = io_flush ? 1'h0 : valid_0_10; // @[playground/src/noop/icache.scala 98:19 99:17 66:26]
  wire  _GEN_141 = io_flush ? 1'h0 : valid_0_11; // @[playground/src/noop/icache.scala 98:19 99:17 66:26]
  wire  _GEN_142 = io_flush ? 1'h0 : valid_0_12; // @[playground/src/noop/icache.scala 98:19 99:17 66:26]
  wire  _GEN_143 = io_flush ? 1'h0 : valid_0_13; // @[playground/src/noop/icache.scala 98:19 99:17 66:26]
  wire  _GEN_144 = io_flush ? 1'h0 : valid_0_14; // @[playground/src/noop/icache.scala 98:19 99:17 66:26]
  wire  _GEN_145 = io_flush ? 1'h0 : valid_0_15; // @[playground/src/noop/icache.scala 98:19 99:17 66:26]
  wire  _GEN_146 = io_flush ? 1'h0 : valid_1_0; // @[playground/src/noop/icache.scala 98:19 99:17 66:26]
  wire  _GEN_147 = io_flush ? 1'h0 : valid_1_1; // @[playground/src/noop/icache.scala 98:19 99:17 66:26]
  wire  _GEN_148 = io_flush ? 1'h0 : valid_1_2; // @[playground/src/noop/icache.scala 98:19 99:17 66:26]
  wire  _GEN_149 = io_flush ? 1'h0 : valid_1_3; // @[playground/src/noop/icache.scala 98:19 99:17 66:26]
  wire  _GEN_150 = io_flush ? 1'h0 : valid_1_4; // @[playground/src/noop/icache.scala 98:19 99:17 66:26]
  wire  _GEN_151 = io_flush ? 1'h0 : valid_1_5; // @[playground/src/noop/icache.scala 98:19 99:17 66:26]
  wire  _GEN_152 = io_flush ? 1'h0 : valid_1_6; // @[playground/src/noop/icache.scala 98:19 99:17 66:26]
  wire  _GEN_153 = io_flush ? 1'h0 : valid_1_7; // @[playground/src/noop/icache.scala 98:19 99:17 66:26]
  wire  _GEN_154 = io_flush ? 1'h0 : valid_1_8; // @[playground/src/noop/icache.scala 98:19 99:17 66:26]
  wire  _GEN_155 = io_flush ? 1'h0 : valid_1_9; // @[playground/src/noop/icache.scala 98:19 99:17 66:26]
  wire  _GEN_156 = io_flush ? 1'h0 : valid_1_10; // @[playground/src/noop/icache.scala 98:19 99:17 66:26]
  wire  _GEN_157 = io_flush ? 1'h0 : valid_1_11; // @[playground/src/noop/icache.scala 98:19 99:17 66:26]
  wire  _GEN_158 = io_flush ? 1'h0 : valid_1_12; // @[playground/src/noop/icache.scala 98:19 99:17 66:26]
  wire  _GEN_159 = io_flush ? 1'h0 : valid_1_13; // @[playground/src/noop/icache.scala 98:19 99:17 66:26]
  wire  _GEN_160 = io_flush ? 1'h0 : valid_1_14; // @[playground/src/noop/icache.scala 98:19 99:17 66:26]
  wire  _GEN_161 = io_flush ? 1'h0 : valid_1_15; // @[playground/src/noop/icache.scala 98:19 99:17 66:26]
  wire  _GEN_162 = io_flush ? 1'h0 : valid_2_0; // @[playground/src/noop/icache.scala 98:19 99:17 66:26]
  wire  _GEN_163 = io_flush ? 1'h0 : valid_2_1; // @[playground/src/noop/icache.scala 98:19 99:17 66:26]
  wire  _GEN_164 = io_flush ? 1'h0 : valid_2_2; // @[playground/src/noop/icache.scala 98:19 99:17 66:26]
  wire  _GEN_165 = io_flush ? 1'h0 : valid_2_3; // @[playground/src/noop/icache.scala 98:19 99:17 66:26]
  wire  _GEN_166 = io_flush ? 1'h0 : valid_2_4; // @[playground/src/noop/icache.scala 98:19 99:17 66:26]
  wire  _GEN_167 = io_flush ? 1'h0 : valid_2_5; // @[playground/src/noop/icache.scala 98:19 99:17 66:26]
  wire  _GEN_168 = io_flush ? 1'h0 : valid_2_6; // @[playground/src/noop/icache.scala 98:19 99:17 66:26]
  wire  _GEN_169 = io_flush ? 1'h0 : valid_2_7; // @[playground/src/noop/icache.scala 98:19 99:17 66:26]
  wire  _GEN_170 = io_flush ? 1'h0 : valid_2_8; // @[playground/src/noop/icache.scala 98:19 99:17 66:26]
  wire  _GEN_171 = io_flush ? 1'h0 : valid_2_9; // @[playground/src/noop/icache.scala 98:19 99:17 66:26]
  wire  _GEN_172 = io_flush ? 1'h0 : valid_2_10; // @[playground/src/noop/icache.scala 98:19 99:17 66:26]
  wire  _GEN_173 = io_flush ? 1'h0 : valid_2_11; // @[playground/src/noop/icache.scala 98:19 99:17 66:26]
  wire  _GEN_174 = io_flush ? 1'h0 : valid_2_12; // @[playground/src/noop/icache.scala 98:19 99:17 66:26]
  wire  _GEN_175 = io_flush ? 1'h0 : valid_2_13; // @[playground/src/noop/icache.scala 98:19 99:17 66:26]
  wire  _GEN_176 = io_flush ? 1'h0 : valid_2_14; // @[playground/src/noop/icache.scala 98:19 99:17 66:26]
  wire  _GEN_177 = io_flush ? 1'h0 : valid_2_15; // @[playground/src/noop/icache.scala 98:19 99:17 66:26]
  wire  _GEN_178 = io_flush ? 1'h0 : valid_3_0; // @[playground/src/noop/icache.scala 98:19 99:17 66:26]
  wire  _GEN_179 = io_flush ? 1'h0 : valid_3_1; // @[playground/src/noop/icache.scala 98:19 99:17 66:26]
  wire  _GEN_180 = io_flush ? 1'h0 : valid_3_2; // @[playground/src/noop/icache.scala 98:19 99:17 66:26]
  wire  _GEN_181 = io_flush ? 1'h0 : valid_3_3; // @[playground/src/noop/icache.scala 98:19 99:17 66:26]
  wire  _GEN_182 = io_flush ? 1'h0 : valid_3_4; // @[playground/src/noop/icache.scala 98:19 99:17 66:26]
  wire  _GEN_183 = io_flush ? 1'h0 : valid_3_5; // @[playground/src/noop/icache.scala 98:19 99:17 66:26]
  wire  _GEN_184 = io_flush ? 1'h0 : valid_3_6; // @[playground/src/noop/icache.scala 98:19 99:17 66:26]
  wire  _GEN_185 = io_flush ? 1'h0 : valid_3_7; // @[playground/src/noop/icache.scala 98:19 99:17 66:26]
  wire  _GEN_186 = io_flush ? 1'h0 : valid_3_8; // @[playground/src/noop/icache.scala 98:19 99:17 66:26]
  wire  _GEN_187 = io_flush ? 1'h0 : valid_3_9; // @[playground/src/noop/icache.scala 98:19 99:17 66:26]
  wire  _GEN_188 = io_flush ? 1'h0 : valid_3_10; // @[playground/src/noop/icache.scala 98:19 99:17 66:26]
  wire  _GEN_189 = io_flush ? 1'h0 : valid_3_11; // @[playground/src/noop/icache.scala 98:19 99:17 66:26]
  wire  _GEN_190 = io_flush ? 1'h0 : valid_3_12; // @[playground/src/noop/icache.scala 98:19 99:17 66:26]
  wire  _GEN_191 = io_flush ? 1'h0 : valid_3_13; // @[playground/src/noop/icache.scala 98:19 99:17 66:26]
  wire  _GEN_192 = io_flush ? 1'h0 : valid_3_14; // @[playground/src/noop/icache.scala 98:19 99:17 66:26]
  wire  _GEN_193 = io_flush ? 1'h0 : valid_3_15; // @[playground/src/noop/icache.scala 98:19 99:17 66:26]
  reg [1:0] state; // @[playground/src/noop/icache.scala 102:24]
  wire [127:0] data_0_rdata = Ram_bw_io_rdata; // @[playground/src/noop/icache.scala 67:{26,26}]
  wire [127:0] data_1_rdata = Ram_bw_1_io_rdata; // @[playground/src/noop/icache.scala 67:{26,26}]
  wire [127:0] _GEN_195 = 2'h1 == matchWay_r[1:0] ? data_1_rdata : data_0_rdata; // @[playground/src/noop/icache.scala 106:{28,28}]
  wire [127:0] data_2_rdata = Ram_bw_2_io_rdata; // @[playground/src/noop/icache.scala 67:{26,26}]
  wire [127:0] _GEN_196 = 2'h2 == matchWay_r[1:0] ? data_2_rdata : _GEN_195; // @[playground/src/noop/icache.scala 106:{28,28}]
  wire [127:0] data_3_rdata = Ram_bw_3_io_rdata; // @[playground/src/noop/icache.scala 67:{26,26}]
  wire [127:0] _GEN_197 = 2'h3 == matchWay_r[1:0] ? data_3_rdata : _GEN_196; // @[playground/src/noop/icache.scala 106:{28,28}]
  wire [5:0] _data_addr_T_1 = state == 2'h2 ? cur_raddr : cur_ram_addr; // @[playground/src/noop/icache.scala 110:31]
  wire  _GEN_1030 = 2'h0 == cur_way[1:0]; // @[playground/src/noop/icache.scala 111:{25,25} playground/src/ram/ram.scala 41:17]
  wire  _GEN_1031 = 2'h1 == cur_way[1:0]; // @[playground/src/noop/icache.scala 111:{25,25} playground/src/ram/ram.scala 41:17]
  wire  _GEN_1032 = 2'h2 == cur_way[1:0]; // @[playground/src/noop/icache.scala 111:{25,25} playground/src/ram/ram.scala 41:17]
  wire  _GEN_1033 = 2'h3 == cur_way[1:0]; // @[playground/src/noop/icache.scala 111:{25,25} playground/src/ram/ram.scala 41:17]
  reg  rdataEn; // @[playground/src/noop/icache.scala 119:30]
  wire  _GEN_494 = rdataEn & io_instAxi_rd_valid & axiOffset[0]; // @[playground/src/noop/icache.scala 115:13 145:49]
  wire  _GEN_763 = 2'h1 == state ? 1'h0 : 2'h2 == state & _GEN_494; // @[playground/src/noop/icache.scala 115:13 121:18]
  wire  wen = 2'h0 == state ? 1'h0 : _GEN_763; // @[playground/src/noop/icache.scala 115:13 121:18]
  wire [127:0] _data_wdata_T = {io_instAxi_rd_bits_data,databuf}; // @[playground/src/noop/icache.scala 113:31]
  reg  raddrEn; // @[playground/src/noop/icache.scala 117:30]
  reg [31:0] raddr; // @[playground/src/noop/icache.scala 118:30]
  wire [31:0] _raddr_T = cur_addr & 32'hffffffc0; // @[playground/src/noop/icache.scala 129:37]
  wire  _GEN_223 = ~hs_in & _io_icRead_ready_T ? 1'h0 : cacheHit; // @[playground/src/noop/icache.scala 123:36 73:13]
  wire  _GEN_230 = raddrEn & io_instAxi_ra_ready | rdataEn; // @[playground/src/noop/icache.scala 137:49 140:25 119:30]
  wire [2:0] _axiOffset_T_1 = axiOffset + 3'h1; // @[playground/src/noop/icache.scala 146:40]
  wire [63:0] _GEN_233 = axiOffset[0] ? databuf : io_instAxi_rd_bits_data; // @[playground/src/noop/icache.scala 147:35 150:29 81:34]
  wire  _GEN_1038 = 2'h0 == matchWay_r[1:0]; // @[playground/src/noop/icache.scala 154:{51,51} 65:26]
  wire  _GEN_1039 = 4'h0 == pre_blockIdx; // @[playground/src/noop/icache.scala 154:{51,51} 65:26]
  wire [21:0] _GEN_234 = 2'h0 == matchWay_r[1:0] & 4'h0 == pre_blockIdx ? pre_instTag : tag_0_0; // @[playground/src/noop/icache.scala 154:{51,51} 65:26]
  wire  _GEN_1041 = 4'h1 == pre_blockIdx; // @[playground/src/noop/icache.scala 154:{51,51} 65:26]
  wire [21:0] _GEN_235 = 2'h0 == matchWay_r[1:0] & 4'h1 == pre_blockIdx ? pre_instTag : tag_0_1; // @[playground/src/noop/icache.scala 154:{51,51} 65:26]
  wire  _GEN_1043 = 4'h2 == pre_blockIdx; // @[playground/src/noop/icache.scala 154:{51,51} 65:26]
  wire [21:0] _GEN_236 = 2'h0 == matchWay_r[1:0] & 4'h2 == pre_blockIdx ? pre_instTag : tag_0_2; // @[playground/src/noop/icache.scala 154:{51,51} 65:26]
  wire  _GEN_1045 = 4'h3 == pre_blockIdx; // @[playground/src/noop/icache.scala 154:{51,51} 65:26]
  wire [21:0] _GEN_237 = 2'h0 == matchWay_r[1:0] & 4'h3 == pre_blockIdx ? pre_instTag : tag_0_3; // @[playground/src/noop/icache.scala 154:{51,51} 65:26]
  wire  _GEN_1047 = 4'h4 == pre_blockIdx; // @[playground/src/noop/icache.scala 154:{51,51} 65:26]
  wire [21:0] _GEN_238 = 2'h0 == matchWay_r[1:0] & 4'h4 == pre_blockIdx ? pre_instTag : tag_0_4; // @[playground/src/noop/icache.scala 154:{51,51} 65:26]
  wire  _GEN_1049 = 4'h5 == pre_blockIdx; // @[playground/src/noop/icache.scala 154:{51,51} 65:26]
  wire [21:0] _GEN_239 = 2'h0 == matchWay_r[1:0] & 4'h5 == pre_blockIdx ? pre_instTag : tag_0_5; // @[playground/src/noop/icache.scala 154:{51,51} 65:26]
  wire  _GEN_1051 = 4'h6 == pre_blockIdx; // @[playground/src/noop/icache.scala 154:{51,51} 65:26]
  wire [21:0] _GEN_240 = 2'h0 == matchWay_r[1:0] & 4'h6 == pre_blockIdx ? pre_instTag : tag_0_6; // @[playground/src/noop/icache.scala 154:{51,51} 65:26]
  wire  _GEN_1053 = 4'h7 == pre_blockIdx; // @[playground/src/noop/icache.scala 154:{51,51} 65:26]
  wire [21:0] _GEN_241 = 2'h0 == matchWay_r[1:0] & 4'h7 == pre_blockIdx ? pre_instTag : tag_0_7; // @[playground/src/noop/icache.scala 154:{51,51} 65:26]
  wire  _GEN_1055 = 4'h8 == pre_blockIdx; // @[playground/src/noop/icache.scala 154:{51,51} 65:26]
  wire [21:0] _GEN_242 = 2'h0 == matchWay_r[1:0] & 4'h8 == pre_blockIdx ? pre_instTag : tag_0_8; // @[playground/src/noop/icache.scala 154:{51,51} 65:26]
  wire  _GEN_1057 = 4'h9 == pre_blockIdx; // @[playground/src/noop/icache.scala 154:{51,51} 65:26]
  wire [21:0] _GEN_243 = 2'h0 == matchWay_r[1:0] & 4'h9 == pre_blockIdx ? pre_instTag : tag_0_9; // @[playground/src/noop/icache.scala 154:{51,51} 65:26]
  wire  _GEN_1059 = 4'ha == pre_blockIdx; // @[playground/src/noop/icache.scala 154:{51,51} 65:26]
  wire [21:0] _GEN_244 = 2'h0 == matchWay_r[1:0] & 4'ha == pre_blockIdx ? pre_instTag : tag_0_10; // @[playground/src/noop/icache.scala 154:{51,51} 65:26]
  wire  _GEN_1061 = 4'hb == pre_blockIdx; // @[playground/src/noop/icache.scala 154:{51,51} 65:26]
  wire [21:0] _GEN_245 = 2'h0 == matchWay_r[1:0] & 4'hb == pre_blockIdx ? pre_instTag : tag_0_11; // @[playground/src/noop/icache.scala 154:{51,51} 65:26]
  wire  _GEN_1063 = 4'hc == pre_blockIdx; // @[playground/src/noop/icache.scala 154:{51,51} 65:26]
  wire [21:0] _GEN_246 = 2'h0 == matchWay_r[1:0] & 4'hc == pre_blockIdx ? pre_instTag : tag_0_12; // @[playground/src/noop/icache.scala 154:{51,51} 65:26]
  wire  _GEN_1065 = 4'hd == pre_blockIdx; // @[playground/src/noop/icache.scala 154:{51,51} 65:26]
  wire [21:0] _GEN_247 = 2'h0 == matchWay_r[1:0] & 4'hd == pre_blockIdx ? pre_instTag : tag_0_13; // @[playground/src/noop/icache.scala 154:{51,51} 65:26]
  wire  _GEN_1067 = 4'he == pre_blockIdx; // @[playground/src/noop/icache.scala 154:{51,51} 65:26]
  wire [21:0] _GEN_248 = 2'h0 == matchWay_r[1:0] & 4'he == pre_blockIdx ? pre_instTag : tag_0_14; // @[playground/src/noop/icache.scala 154:{51,51} 65:26]
  wire  _GEN_1069 = 4'hf == pre_blockIdx; // @[playground/src/noop/icache.scala 154:{51,51} 65:26]
  wire [21:0] _GEN_249 = 2'h0 == matchWay_r[1:0] & 4'hf == pre_blockIdx ? pre_instTag : tag_0_15; // @[playground/src/noop/icache.scala 154:{51,51} 65:26]
  wire  _GEN_1070 = 2'h1 == matchWay_r[1:0]; // @[playground/src/noop/icache.scala 154:{51,51} 65:26]
  wire [21:0] _GEN_250 = 2'h1 == matchWay_r[1:0] & 4'h0 == pre_blockIdx ? pre_instTag : tag_1_0; // @[playground/src/noop/icache.scala 154:{51,51} 65:26]
  wire [21:0] _GEN_251 = 2'h1 == matchWay_r[1:0] & 4'h1 == pre_blockIdx ? pre_instTag : tag_1_1; // @[playground/src/noop/icache.scala 154:{51,51} 65:26]
  wire [21:0] _GEN_252 = 2'h1 == matchWay_r[1:0] & 4'h2 == pre_blockIdx ? pre_instTag : tag_1_2; // @[playground/src/noop/icache.scala 154:{51,51} 65:26]
  wire [21:0] _GEN_253 = 2'h1 == matchWay_r[1:0] & 4'h3 == pre_blockIdx ? pre_instTag : tag_1_3; // @[playground/src/noop/icache.scala 154:{51,51} 65:26]
  wire [21:0] _GEN_254 = 2'h1 == matchWay_r[1:0] & 4'h4 == pre_blockIdx ? pre_instTag : tag_1_4; // @[playground/src/noop/icache.scala 154:{51,51} 65:26]
  wire [21:0] _GEN_255 = 2'h1 == matchWay_r[1:0] & 4'h5 == pre_blockIdx ? pre_instTag : tag_1_5; // @[playground/src/noop/icache.scala 154:{51,51} 65:26]
  wire [21:0] _GEN_256 = 2'h1 == matchWay_r[1:0] & 4'h6 == pre_blockIdx ? pre_instTag : tag_1_6; // @[playground/src/noop/icache.scala 154:{51,51} 65:26]
  wire [21:0] _GEN_257 = 2'h1 == matchWay_r[1:0] & 4'h7 == pre_blockIdx ? pre_instTag : tag_1_7; // @[playground/src/noop/icache.scala 154:{51,51} 65:26]
  wire [21:0] _GEN_258 = 2'h1 == matchWay_r[1:0] & 4'h8 == pre_blockIdx ? pre_instTag : tag_1_8; // @[playground/src/noop/icache.scala 154:{51,51} 65:26]
  wire [21:0] _GEN_259 = 2'h1 == matchWay_r[1:0] & 4'h9 == pre_blockIdx ? pre_instTag : tag_1_9; // @[playground/src/noop/icache.scala 154:{51,51} 65:26]
  wire [21:0] _GEN_260 = 2'h1 == matchWay_r[1:0] & 4'ha == pre_blockIdx ? pre_instTag : tag_1_10; // @[playground/src/noop/icache.scala 154:{51,51} 65:26]
  wire [21:0] _GEN_261 = 2'h1 == matchWay_r[1:0] & 4'hb == pre_blockIdx ? pre_instTag : tag_1_11; // @[playground/src/noop/icache.scala 154:{51,51} 65:26]
  wire [21:0] _GEN_262 = 2'h1 == matchWay_r[1:0] & 4'hc == pre_blockIdx ? pre_instTag : tag_1_12; // @[playground/src/noop/icache.scala 154:{51,51} 65:26]
  wire [21:0] _GEN_263 = 2'h1 == matchWay_r[1:0] & 4'hd == pre_blockIdx ? pre_instTag : tag_1_13; // @[playground/src/noop/icache.scala 154:{51,51} 65:26]
  wire [21:0] _GEN_264 = 2'h1 == matchWay_r[1:0] & 4'he == pre_blockIdx ? pre_instTag : tag_1_14; // @[playground/src/noop/icache.scala 154:{51,51} 65:26]
  wire [21:0] _GEN_265 = 2'h1 == matchWay_r[1:0] & 4'hf == pre_blockIdx ? pre_instTag : tag_1_15; // @[playground/src/noop/icache.scala 154:{51,51} 65:26]
  wire  _GEN_1102 = 2'h2 == matchWay_r[1:0]; // @[playground/src/noop/icache.scala 154:{51,51} 65:26]
  wire [21:0] _GEN_266 = 2'h2 == matchWay_r[1:0] & 4'h0 == pre_blockIdx ? pre_instTag : tag_2_0; // @[playground/src/noop/icache.scala 154:{51,51} 65:26]
  wire [21:0] _GEN_267 = 2'h2 == matchWay_r[1:0] & 4'h1 == pre_blockIdx ? pre_instTag : tag_2_1; // @[playground/src/noop/icache.scala 154:{51,51} 65:26]
  wire [21:0] _GEN_268 = 2'h2 == matchWay_r[1:0] & 4'h2 == pre_blockIdx ? pre_instTag : tag_2_2; // @[playground/src/noop/icache.scala 154:{51,51} 65:26]
  wire [21:0] _GEN_269 = 2'h2 == matchWay_r[1:0] & 4'h3 == pre_blockIdx ? pre_instTag : tag_2_3; // @[playground/src/noop/icache.scala 154:{51,51} 65:26]
  wire [21:0] _GEN_270 = 2'h2 == matchWay_r[1:0] & 4'h4 == pre_blockIdx ? pre_instTag : tag_2_4; // @[playground/src/noop/icache.scala 154:{51,51} 65:26]
  wire [21:0] _GEN_271 = 2'h2 == matchWay_r[1:0] & 4'h5 == pre_blockIdx ? pre_instTag : tag_2_5; // @[playground/src/noop/icache.scala 154:{51,51} 65:26]
  wire [21:0] _GEN_272 = 2'h2 == matchWay_r[1:0] & 4'h6 == pre_blockIdx ? pre_instTag : tag_2_6; // @[playground/src/noop/icache.scala 154:{51,51} 65:26]
  wire [21:0] _GEN_273 = 2'h2 == matchWay_r[1:0] & 4'h7 == pre_blockIdx ? pre_instTag : tag_2_7; // @[playground/src/noop/icache.scala 154:{51,51} 65:26]
  wire [21:0] _GEN_274 = 2'h2 == matchWay_r[1:0] & 4'h8 == pre_blockIdx ? pre_instTag : tag_2_8; // @[playground/src/noop/icache.scala 154:{51,51} 65:26]
  wire [21:0] _GEN_275 = 2'h2 == matchWay_r[1:0] & 4'h9 == pre_blockIdx ? pre_instTag : tag_2_9; // @[playground/src/noop/icache.scala 154:{51,51} 65:26]
  wire [21:0] _GEN_276 = 2'h2 == matchWay_r[1:0] & 4'ha == pre_blockIdx ? pre_instTag : tag_2_10; // @[playground/src/noop/icache.scala 154:{51,51} 65:26]
  wire [21:0] _GEN_277 = 2'h2 == matchWay_r[1:0] & 4'hb == pre_blockIdx ? pre_instTag : tag_2_11; // @[playground/src/noop/icache.scala 154:{51,51} 65:26]
  wire [21:0] _GEN_278 = 2'h2 == matchWay_r[1:0] & 4'hc == pre_blockIdx ? pre_instTag : tag_2_12; // @[playground/src/noop/icache.scala 154:{51,51} 65:26]
  wire [21:0] _GEN_279 = 2'h2 == matchWay_r[1:0] & 4'hd == pre_blockIdx ? pre_instTag : tag_2_13; // @[playground/src/noop/icache.scala 154:{51,51} 65:26]
  wire [21:0] _GEN_280 = 2'h2 == matchWay_r[1:0] & 4'he == pre_blockIdx ? pre_instTag : tag_2_14; // @[playground/src/noop/icache.scala 154:{51,51} 65:26]
  wire [21:0] _GEN_281 = 2'h2 == matchWay_r[1:0] & 4'hf == pre_blockIdx ? pre_instTag : tag_2_15; // @[playground/src/noop/icache.scala 154:{51,51} 65:26]
  wire  _GEN_1134 = 2'h3 == matchWay_r[1:0]; // @[playground/src/noop/icache.scala 154:{51,51} 65:26]
  wire [21:0] _GEN_282 = 2'h3 == matchWay_r[1:0] & 4'h0 == pre_blockIdx ? pre_instTag : tag_3_0; // @[playground/src/noop/icache.scala 154:{51,51} 65:26]
  wire [21:0] _GEN_283 = 2'h3 == matchWay_r[1:0] & 4'h1 == pre_blockIdx ? pre_instTag : tag_3_1; // @[playground/src/noop/icache.scala 154:{51,51} 65:26]
  wire [21:0] _GEN_284 = 2'h3 == matchWay_r[1:0] & 4'h2 == pre_blockIdx ? pre_instTag : tag_3_2; // @[playground/src/noop/icache.scala 154:{51,51} 65:26]
  wire [21:0] _GEN_285 = 2'h3 == matchWay_r[1:0] & 4'h3 == pre_blockIdx ? pre_instTag : tag_3_3; // @[playground/src/noop/icache.scala 154:{51,51} 65:26]
  wire [21:0] _GEN_286 = 2'h3 == matchWay_r[1:0] & 4'h4 == pre_blockIdx ? pre_instTag : tag_3_4; // @[playground/src/noop/icache.scala 154:{51,51} 65:26]
  wire [21:0] _GEN_287 = 2'h3 == matchWay_r[1:0] & 4'h5 == pre_blockIdx ? pre_instTag : tag_3_5; // @[playground/src/noop/icache.scala 154:{51,51} 65:26]
  wire [21:0] _GEN_288 = 2'h3 == matchWay_r[1:0] & 4'h6 == pre_blockIdx ? pre_instTag : tag_3_6; // @[playground/src/noop/icache.scala 154:{51,51} 65:26]
  wire [21:0] _GEN_289 = 2'h3 == matchWay_r[1:0] & 4'h7 == pre_blockIdx ? pre_instTag : tag_3_7; // @[playground/src/noop/icache.scala 154:{51,51} 65:26]
  wire [21:0] _GEN_290 = 2'h3 == matchWay_r[1:0] & 4'h8 == pre_blockIdx ? pre_instTag : tag_3_8; // @[playground/src/noop/icache.scala 154:{51,51} 65:26]
  wire [21:0] _GEN_291 = 2'h3 == matchWay_r[1:0] & 4'h9 == pre_blockIdx ? pre_instTag : tag_3_9; // @[playground/src/noop/icache.scala 154:{51,51} 65:26]
  wire [21:0] _GEN_292 = 2'h3 == matchWay_r[1:0] & 4'ha == pre_blockIdx ? pre_instTag : tag_3_10; // @[playground/src/noop/icache.scala 154:{51,51} 65:26]
  wire [21:0] _GEN_293 = 2'h3 == matchWay_r[1:0] & 4'hb == pre_blockIdx ? pre_instTag : tag_3_11; // @[playground/src/noop/icache.scala 154:{51,51} 65:26]
  wire [21:0] _GEN_294 = 2'h3 == matchWay_r[1:0] & 4'hc == pre_blockIdx ? pre_instTag : tag_3_12; // @[playground/src/noop/icache.scala 154:{51,51} 65:26]
  wire [21:0] _GEN_295 = 2'h3 == matchWay_r[1:0] & 4'hd == pre_blockIdx ? pre_instTag : tag_3_13; // @[playground/src/noop/icache.scala 154:{51,51} 65:26]
  wire [21:0] _GEN_296 = 2'h3 == matchWay_r[1:0] & 4'he == pre_blockIdx ? pre_instTag : tag_3_14; // @[playground/src/noop/icache.scala 154:{51,51} 65:26]
  wire [21:0] _GEN_297 = 2'h3 == matchWay_r[1:0] & 4'hf == pre_blockIdx ? pre_instTag : tag_3_15; // @[playground/src/noop/icache.scala 154:{51,51} 65:26]
  wire  _GEN_298 = _GEN_1038 & _GEN_1039 | _GEN_130; // @[playground/src/noop/icache.scala 155:{53,53}]
  wire  _GEN_299 = _GEN_1038 & _GEN_1041 | _GEN_131; // @[playground/src/noop/icache.scala 155:{53,53}]
  wire  _GEN_300 = _GEN_1038 & _GEN_1043 | _GEN_132; // @[playground/src/noop/icache.scala 155:{53,53}]
  wire  _GEN_301 = _GEN_1038 & _GEN_1045 | _GEN_133; // @[playground/src/noop/icache.scala 155:{53,53}]
  wire  _GEN_302 = _GEN_1038 & _GEN_1047 | _GEN_134; // @[playground/src/noop/icache.scala 155:{53,53}]
  wire  _GEN_303 = _GEN_1038 & _GEN_1049 | _GEN_135; // @[playground/src/noop/icache.scala 155:{53,53}]
  wire  _GEN_304 = _GEN_1038 & _GEN_1051 | _GEN_136; // @[playground/src/noop/icache.scala 155:{53,53}]
  wire  _GEN_305 = _GEN_1038 & _GEN_1053 | _GEN_137; // @[playground/src/noop/icache.scala 155:{53,53}]
  wire  _GEN_306 = _GEN_1038 & _GEN_1055 | _GEN_138; // @[playground/src/noop/icache.scala 155:{53,53}]
  wire  _GEN_307 = _GEN_1038 & _GEN_1057 | _GEN_139; // @[playground/src/noop/icache.scala 155:{53,53}]
  wire  _GEN_308 = _GEN_1038 & _GEN_1059 | _GEN_140; // @[playground/src/noop/icache.scala 155:{53,53}]
  wire  _GEN_309 = _GEN_1038 & _GEN_1061 | _GEN_141; // @[playground/src/noop/icache.scala 155:{53,53}]
  wire  _GEN_310 = _GEN_1038 & _GEN_1063 | _GEN_142; // @[playground/src/noop/icache.scala 155:{53,53}]
  wire  _GEN_311 = _GEN_1038 & _GEN_1065 | _GEN_143; // @[playground/src/noop/icache.scala 155:{53,53}]
  wire  _GEN_312 = _GEN_1038 & _GEN_1067 | _GEN_144; // @[playground/src/noop/icache.scala 155:{53,53}]
  wire  _GEN_313 = _GEN_1038 & _GEN_1069 | _GEN_145; // @[playground/src/noop/icache.scala 155:{53,53}]
  wire  _GEN_314 = _GEN_1070 & _GEN_1039 | _GEN_146; // @[playground/src/noop/icache.scala 155:{53,53}]
  wire  _GEN_315 = _GEN_1070 & _GEN_1041 | _GEN_147; // @[playground/src/noop/icache.scala 155:{53,53}]
  wire  _GEN_316 = _GEN_1070 & _GEN_1043 | _GEN_148; // @[playground/src/noop/icache.scala 155:{53,53}]
  wire  _GEN_317 = _GEN_1070 & _GEN_1045 | _GEN_149; // @[playground/src/noop/icache.scala 155:{53,53}]
  wire  _GEN_318 = _GEN_1070 & _GEN_1047 | _GEN_150; // @[playground/src/noop/icache.scala 155:{53,53}]
  wire  _GEN_319 = _GEN_1070 & _GEN_1049 | _GEN_151; // @[playground/src/noop/icache.scala 155:{53,53}]
  wire  _GEN_320 = _GEN_1070 & _GEN_1051 | _GEN_152; // @[playground/src/noop/icache.scala 155:{53,53}]
  wire  _GEN_321 = _GEN_1070 & _GEN_1053 | _GEN_153; // @[playground/src/noop/icache.scala 155:{53,53}]
  wire  _GEN_322 = _GEN_1070 & _GEN_1055 | _GEN_154; // @[playground/src/noop/icache.scala 155:{53,53}]
  wire  _GEN_323 = _GEN_1070 & _GEN_1057 | _GEN_155; // @[playground/src/noop/icache.scala 155:{53,53}]
  wire  _GEN_324 = _GEN_1070 & _GEN_1059 | _GEN_156; // @[playground/src/noop/icache.scala 155:{53,53}]
  wire  _GEN_325 = _GEN_1070 & _GEN_1061 | _GEN_157; // @[playground/src/noop/icache.scala 155:{53,53}]
  wire  _GEN_326 = _GEN_1070 & _GEN_1063 | _GEN_158; // @[playground/src/noop/icache.scala 155:{53,53}]
  wire  _GEN_327 = _GEN_1070 & _GEN_1065 | _GEN_159; // @[playground/src/noop/icache.scala 155:{53,53}]
  wire  _GEN_328 = _GEN_1070 & _GEN_1067 | _GEN_160; // @[playground/src/noop/icache.scala 155:{53,53}]
  wire  _GEN_329 = _GEN_1070 & _GEN_1069 | _GEN_161; // @[playground/src/noop/icache.scala 155:{53,53}]
  wire  _GEN_330 = _GEN_1102 & _GEN_1039 | _GEN_162; // @[playground/src/noop/icache.scala 155:{53,53}]
  wire  _GEN_331 = _GEN_1102 & _GEN_1041 | _GEN_163; // @[playground/src/noop/icache.scala 155:{53,53}]
  wire  _GEN_332 = _GEN_1102 & _GEN_1043 | _GEN_164; // @[playground/src/noop/icache.scala 155:{53,53}]
  wire  _GEN_333 = _GEN_1102 & _GEN_1045 | _GEN_165; // @[playground/src/noop/icache.scala 155:{53,53}]
  wire  _GEN_334 = _GEN_1102 & _GEN_1047 | _GEN_166; // @[playground/src/noop/icache.scala 155:{53,53}]
  wire  _GEN_335 = _GEN_1102 & _GEN_1049 | _GEN_167; // @[playground/src/noop/icache.scala 155:{53,53}]
  wire  _GEN_336 = _GEN_1102 & _GEN_1051 | _GEN_168; // @[playground/src/noop/icache.scala 155:{53,53}]
  wire  _GEN_337 = _GEN_1102 & _GEN_1053 | _GEN_169; // @[playground/src/noop/icache.scala 155:{53,53}]
  wire  _GEN_338 = _GEN_1102 & _GEN_1055 | _GEN_170; // @[playground/src/noop/icache.scala 155:{53,53}]
  wire  _GEN_339 = _GEN_1102 & _GEN_1057 | _GEN_171; // @[playground/src/noop/icache.scala 155:{53,53}]
  wire  _GEN_340 = _GEN_1102 & _GEN_1059 | _GEN_172; // @[playground/src/noop/icache.scala 155:{53,53}]
  wire  _GEN_341 = _GEN_1102 & _GEN_1061 | _GEN_173; // @[playground/src/noop/icache.scala 155:{53,53}]
  wire  _GEN_342 = _GEN_1102 & _GEN_1063 | _GEN_174; // @[playground/src/noop/icache.scala 155:{53,53}]
  wire  _GEN_343 = _GEN_1102 & _GEN_1065 | _GEN_175; // @[playground/src/noop/icache.scala 155:{53,53}]
  wire  _GEN_344 = _GEN_1102 & _GEN_1067 | _GEN_176; // @[playground/src/noop/icache.scala 155:{53,53}]
  wire  _GEN_345 = _GEN_1102 & _GEN_1069 | _GEN_177; // @[playground/src/noop/icache.scala 155:{53,53}]
  wire  _GEN_346 = _GEN_1134 & _GEN_1039 | _GEN_178; // @[playground/src/noop/icache.scala 155:{53,53}]
  wire  _GEN_347 = _GEN_1134 & _GEN_1041 | _GEN_179; // @[playground/src/noop/icache.scala 155:{53,53}]
  wire  _GEN_348 = _GEN_1134 & _GEN_1043 | _GEN_180; // @[playground/src/noop/icache.scala 155:{53,53}]
  wire  _GEN_349 = _GEN_1134 & _GEN_1045 | _GEN_181; // @[playground/src/noop/icache.scala 155:{53,53}]
  wire  _GEN_350 = _GEN_1134 & _GEN_1047 | _GEN_182; // @[playground/src/noop/icache.scala 155:{53,53}]
  wire  _GEN_351 = _GEN_1134 & _GEN_1049 | _GEN_183; // @[playground/src/noop/icache.scala 155:{53,53}]
  wire  _GEN_352 = _GEN_1134 & _GEN_1051 | _GEN_184; // @[playground/src/noop/icache.scala 155:{53,53}]
  wire  _GEN_353 = _GEN_1134 & _GEN_1053 | _GEN_185; // @[playground/src/noop/icache.scala 155:{53,53}]
  wire  _GEN_354 = _GEN_1134 & _GEN_1055 | _GEN_186; // @[playground/src/noop/icache.scala 155:{53,53}]
  wire  _GEN_355 = _GEN_1134 & _GEN_1057 | _GEN_187; // @[playground/src/noop/icache.scala 155:{53,53}]
  wire  _GEN_356 = _GEN_1134 & _GEN_1059 | _GEN_188; // @[playground/src/noop/icache.scala 155:{53,53}]
  wire  _GEN_357 = _GEN_1134 & _GEN_1061 | _GEN_189; // @[playground/src/noop/icache.scala 155:{53,53}]
  wire  _GEN_358 = _GEN_1134 & _GEN_1063 | _GEN_190; // @[playground/src/noop/icache.scala 155:{53,53}]
  wire  _GEN_359 = _GEN_1134 & _GEN_1065 | _GEN_191; // @[playground/src/noop/icache.scala 155:{53,53}]
  wire  _GEN_360 = _GEN_1134 & _GEN_1067 | _GEN_192; // @[playground/src/noop/icache.scala 155:{53,53}]
  wire  _GEN_361 = _GEN_1134 & _GEN_1069 | _GEN_193; // @[playground/src/noop/icache.scala 155:{53,53}]
  wire  _GEN_362 = io_instAxi_rd_bits_last ? 1'h0 : rdataEn; // @[playground/src/noop/icache.scala 152:46 153:29 119:30]
  wire [21:0] _GEN_363 = io_instAxi_rd_bits_last ? _GEN_234 : tag_0_0; // @[playground/src/noop/icache.scala 152:46 65:26]
  wire [21:0] _GEN_364 = io_instAxi_rd_bits_last ? _GEN_235 : tag_0_1; // @[playground/src/noop/icache.scala 152:46 65:26]
  wire [21:0] _GEN_365 = io_instAxi_rd_bits_last ? _GEN_236 : tag_0_2; // @[playground/src/noop/icache.scala 152:46 65:26]
  wire [21:0] _GEN_366 = io_instAxi_rd_bits_last ? _GEN_237 : tag_0_3; // @[playground/src/noop/icache.scala 152:46 65:26]
  wire [21:0] _GEN_367 = io_instAxi_rd_bits_last ? _GEN_238 : tag_0_4; // @[playground/src/noop/icache.scala 152:46 65:26]
  wire [21:0] _GEN_368 = io_instAxi_rd_bits_last ? _GEN_239 : tag_0_5; // @[playground/src/noop/icache.scala 152:46 65:26]
  wire [21:0] _GEN_369 = io_instAxi_rd_bits_last ? _GEN_240 : tag_0_6; // @[playground/src/noop/icache.scala 152:46 65:26]
  wire [21:0] _GEN_370 = io_instAxi_rd_bits_last ? _GEN_241 : tag_0_7; // @[playground/src/noop/icache.scala 152:46 65:26]
  wire [21:0] _GEN_371 = io_instAxi_rd_bits_last ? _GEN_242 : tag_0_8; // @[playground/src/noop/icache.scala 152:46 65:26]
  wire [21:0] _GEN_372 = io_instAxi_rd_bits_last ? _GEN_243 : tag_0_9; // @[playground/src/noop/icache.scala 152:46 65:26]
  wire [21:0] _GEN_373 = io_instAxi_rd_bits_last ? _GEN_244 : tag_0_10; // @[playground/src/noop/icache.scala 152:46 65:26]
  wire [21:0] _GEN_374 = io_instAxi_rd_bits_last ? _GEN_245 : tag_0_11; // @[playground/src/noop/icache.scala 152:46 65:26]
  wire [21:0] _GEN_375 = io_instAxi_rd_bits_last ? _GEN_246 : tag_0_12; // @[playground/src/noop/icache.scala 152:46 65:26]
  wire [21:0] _GEN_376 = io_instAxi_rd_bits_last ? _GEN_247 : tag_0_13; // @[playground/src/noop/icache.scala 152:46 65:26]
  wire [21:0] _GEN_377 = io_instAxi_rd_bits_last ? _GEN_248 : tag_0_14; // @[playground/src/noop/icache.scala 152:46 65:26]
  wire [21:0] _GEN_378 = io_instAxi_rd_bits_last ? _GEN_249 : tag_0_15; // @[playground/src/noop/icache.scala 152:46 65:26]
  wire [21:0] _GEN_379 = io_instAxi_rd_bits_last ? _GEN_250 : tag_1_0; // @[playground/src/noop/icache.scala 152:46 65:26]
  wire [21:0] _GEN_380 = io_instAxi_rd_bits_last ? _GEN_251 : tag_1_1; // @[playground/src/noop/icache.scala 152:46 65:26]
  wire [21:0] _GEN_381 = io_instAxi_rd_bits_last ? _GEN_252 : tag_1_2; // @[playground/src/noop/icache.scala 152:46 65:26]
  wire [21:0] _GEN_382 = io_instAxi_rd_bits_last ? _GEN_253 : tag_1_3; // @[playground/src/noop/icache.scala 152:46 65:26]
  wire [21:0] _GEN_383 = io_instAxi_rd_bits_last ? _GEN_254 : tag_1_4; // @[playground/src/noop/icache.scala 152:46 65:26]
  wire [21:0] _GEN_384 = io_instAxi_rd_bits_last ? _GEN_255 : tag_1_5; // @[playground/src/noop/icache.scala 152:46 65:26]
  wire [21:0] _GEN_385 = io_instAxi_rd_bits_last ? _GEN_256 : tag_1_6; // @[playground/src/noop/icache.scala 152:46 65:26]
  wire [21:0] _GEN_386 = io_instAxi_rd_bits_last ? _GEN_257 : tag_1_7; // @[playground/src/noop/icache.scala 152:46 65:26]
  wire [21:0] _GEN_387 = io_instAxi_rd_bits_last ? _GEN_258 : tag_1_8; // @[playground/src/noop/icache.scala 152:46 65:26]
  wire [21:0] _GEN_388 = io_instAxi_rd_bits_last ? _GEN_259 : tag_1_9; // @[playground/src/noop/icache.scala 152:46 65:26]
  wire [21:0] _GEN_389 = io_instAxi_rd_bits_last ? _GEN_260 : tag_1_10; // @[playground/src/noop/icache.scala 152:46 65:26]
  wire [21:0] _GEN_390 = io_instAxi_rd_bits_last ? _GEN_261 : tag_1_11; // @[playground/src/noop/icache.scala 152:46 65:26]
  wire [21:0] _GEN_391 = io_instAxi_rd_bits_last ? _GEN_262 : tag_1_12; // @[playground/src/noop/icache.scala 152:46 65:26]
  wire [21:0] _GEN_392 = io_instAxi_rd_bits_last ? _GEN_263 : tag_1_13; // @[playground/src/noop/icache.scala 152:46 65:26]
  wire [21:0] _GEN_393 = io_instAxi_rd_bits_last ? _GEN_264 : tag_1_14; // @[playground/src/noop/icache.scala 152:46 65:26]
  wire [21:0] _GEN_394 = io_instAxi_rd_bits_last ? _GEN_265 : tag_1_15; // @[playground/src/noop/icache.scala 152:46 65:26]
  wire [21:0] _GEN_395 = io_instAxi_rd_bits_last ? _GEN_266 : tag_2_0; // @[playground/src/noop/icache.scala 152:46 65:26]
  wire [21:0] _GEN_396 = io_instAxi_rd_bits_last ? _GEN_267 : tag_2_1; // @[playground/src/noop/icache.scala 152:46 65:26]
  wire [21:0] _GEN_397 = io_instAxi_rd_bits_last ? _GEN_268 : tag_2_2; // @[playground/src/noop/icache.scala 152:46 65:26]
  wire [21:0] _GEN_398 = io_instAxi_rd_bits_last ? _GEN_269 : tag_2_3; // @[playground/src/noop/icache.scala 152:46 65:26]
  wire [21:0] _GEN_399 = io_instAxi_rd_bits_last ? _GEN_270 : tag_2_4; // @[playground/src/noop/icache.scala 152:46 65:26]
  wire [21:0] _GEN_400 = io_instAxi_rd_bits_last ? _GEN_271 : tag_2_5; // @[playground/src/noop/icache.scala 152:46 65:26]
  wire [21:0] _GEN_401 = io_instAxi_rd_bits_last ? _GEN_272 : tag_2_6; // @[playground/src/noop/icache.scala 152:46 65:26]
  wire [21:0] _GEN_402 = io_instAxi_rd_bits_last ? _GEN_273 : tag_2_7; // @[playground/src/noop/icache.scala 152:46 65:26]
  wire [21:0] _GEN_403 = io_instAxi_rd_bits_last ? _GEN_274 : tag_2_8; // @[playground/src/noop/icache.scala 152:46 65:26]
  wire [21:0] _GEN_404 = io_instAxi_rd_bits_last ? _GEN_275 : tag_2_9; // @[playground/src/noop/icache.scala 152:46 65:26]
  wire [21:0] _GEN_405 = io_instAxi_rd_bits_last ? _GEN_276 : tag_2_10; // @[playground/src/noop/icache.scala 152:46 65:26]
  wire [21:0] _GEN_406 = io_instAxi_rd_bits_last ? _GEN_277 : tag_2_11; // @[playground/src/noop/icache.scala 152:46 65:26]
  wire [21:0] _GEN_407 = io_instAxi_rd_bits_last ? _GEN_278 : tag_2_12; // @[playground/src/noop/icache.scala 152:46 65:26]
  wire [21:0] _GEN_408 = io_instAxi_rd_bits_last ? _GEN_279 : tag_2_13; // @[playground/src/noop/icache.scala 152:46 65:26]
  wire [21:0] _GEN_409 = io_instAxi_rd_bits_last ? _GEN_280 : tag_2_14; // @[playground/src/noop/icache.scala 152:46 65:26]
  wire [21:0] _GEN_410 = io_instAxi_rd_bits_last ? _GEN_281 : tag_2_15; // @[playground/src/noop/icache.scala 152:46 65:26]
  wire [21:0] _GEN_411 = io_instAxi_rd_bits_last ? _GEN_282 : tag_3_0; // @[playground/src/noop/icache.scala 152:46 65:26]
  wire [21:0] _GEN_412 = io_instAxi_rd_bits_last ? _GEN_283 : tag_3_1; // @[playground/src/noop/icache.scala 152:46 65:26]
  wire [21:0] _GEN_413 = io_instAxi_rd_bits_last ? _GEN_284 : tag_3_2; // @[playground/src/noop/icache.scala 152:46 65:26]
  wire [21:0] _GEN_414 = io_instAxi_rd_bits_last ? _GEN_285 : tag_3_3; // @[playground/src/noop/icache.scala 152:46 65:26]
  wire [21:0] _GEN_415 = io_instAxi_rd_bits_last ? _GEN_286 : tag_3_4; // @[playground/src/noop/icache.scala 152:46 65:26]
  wire [21:0] _GEN_416 = io_instAxi_rd_bits_last ? _GEN_287 : tag_3_5; // @[playground/src/noop/icache.scala 152:46 65:26]
  wire [21:0] _GEN_417 = io_instAxi_rd_bits_last ? _GEN_288 : tag_3_6; // @[playground/src/noop/icache.scala 152:46 65:26]
  wire [21:0] _GEN_418 = io_instAxi_rd_bits_last ? _GEN_289 : tag_3_7; // @[playground/src/noop/icache.scala 152:46 65:26]
  wire [21:0] _GEN_419 = io_instAxi_rd_bits_last ? _GEN_290 : tag_3_8; // @[playground/src/noop/icache.scala 152:46 65:26]
  wire [21:0] _GEN_420 = io_instAxi_rd_bits_last ? _GEN_291 : tag_3_9; // @[playground/src/noop/icache.scala 152:46 65:26]
  wire [21:0] _GEN_421 = io_instAxi_rd_bits_last ? _GEN_292 : tag_3_10; // @[playground/src/noop/icache.scala 152:46 65:26]
  wire [21:0] _GEN_422 = io_instAxi_rd_bits_last ? _GEN_293 : tag_3_11; // @[playground/src/noop/icache.scala 152:46 65:26]
  wire [21:0] _GEN_423 = io_instAxi_rd_bits_last ? _GEN_294 : tag_3_12; // @[playground/src/noop/icache.scala 152:46 65:26]
  wire [21:0] _GEN_424 = io_instAxi_rd_bits_last ? _GEN_295 : tag_3_13; // @[playground/src/noop/icache.scala 152:46 65:26]
  wire [21:0] _GEN_425 = io_instAxi_rd_bits_last ? _GEN_296 : tag_3_14; // @[playground/src/noop/icache.scala 152:46 65:26]
  wire [21:0] _GEN_426 = io_instAxi_rd_bits_last ? _GEN_297 : tag_3_15; // @[playground/src/noop/icache.scala 152:46 65:26]
  wire  _GEN_427 = io_instAxi_rd_bits_last ? _GEN_298 : _GEN_130; // @[playground/src/noop/icache.scala 152:46]
  wire  _GEN_428 = io_instAxi_rd_bits_last ? _GEN_299 : _GEN_131; // @[playground/src/noop/icache.scala 152:46]
  wire  _GEN_429 = io_instAxi_rd_bits_last ? _GEN_300 : _GEN_132; // @[playground/src/noop/icache.scala 152:46]
  wire  _GEN_430 = io_instAxi_rd_bits_last ? _GEN_301 : _GEN_133; // @[playground/src/noop/icache.scala 152:46]
  wire  _GEN_431 = io_instAxi_rd_bits_last ? _GEN_302 : _GEN_134; // @[playground/src/noop/icache.scala 152:46]
  wire  _GEN_432 = io_instAxi_rd_bits_last ? _GEN_303 : _GEN_135; // @[playground/src/noop/icache.scala 152:46]
  wire  _GEN_433 = io_instAxi_rd_bits_last ? _GEN_304 : _GEN_136; // @[playground/src/noop/icache.scala 152:46]
  wire  _GEN_434 = io_instAxi_rd_bits_last ? _GEN_305 : _GEN_137; // @[playground/src/noop/icache.scala 152:46]
  wire  _GEN_435 = io_instAxi_rd_bits_last ? _GEN_306 : _GEN_138; // @[playground/src/noop/icache.scala 152:46]
  wire  _GEN_436 = io_instAxi_rd_bits_last ? _GEN_307 : _GEN_139; // @[playground/src/noop/icache.scala 152:46]
  wire  _GEN_437 = io_instAxi_rd_bits_last ? _GEN_308 : _GEN_140; // @[playground/src/noop/icache.scala 152:46]
  wire  _GEN_438 = io_instAxi_rd_bits_last ? _GEN_309 : _GEN_141; // @[playground/src/noop/icache.scala 152:46]
  wire  _GEN_439 = io_instAxi_rd_bits_last ? _GEN_310 : _GEN_142; // @[playground/src/noop/icache.scala 152:46]
  wire  _GEN_440 = io_instAxi_rd_bits_last ? _GEN_311 : _GEN_143; // @[playground/src/noop/icache.scala 152:46]
  wire  _GEN_441 = io_instAxi_rd_bits_last ? _GEN_312 : _GEN_144; // @[playground/src/noop/icache.scala 152:46]
  wire  _GEN_442 = io_instAxi_rd_bits_last ? _GEN_313 : _GEN_145; // @[playground/src/noop/icache.scala 152:46]
  wire  _GEN_443 = io_instAxi_rd_bits_last ? _GEN_314 : _GEN_146; // @[playground/src/noop/icache.scala 152:46]
  wire  _GEN_444 = io_instAxi_rd_bits_last ? _GEN_315 : _GEN_147; // @[playground/src/noop/icache.scala 152:46]
  wire  _GEN_445 = io_instAxi_rd_bits_last ? _GEN_316 : _GEN_148; // @[playground/src/noop/icache.scala 152:46]
  wire  _GEN_446 = io_instAxi_rd_bits_last ? _GEN_317 : _GEN_149; // @[playground/src/noop/icache.scala 152:46]
  wire  _GEN_447 = io_instAxi_rd_bits_last ? _GEN_318 : _GEN_150; // @[playground/src/noop/icache.scala 152:46]
  wire  _GEN_448 = io_instAxi_rd_bits_last ? _GEN_319 : _GEN_151; // @[playground/src/noop/icache.scala 152:46]
  wire  _GEN_449 = io_instAxi_rd_bits_last ? _GEN_320 : _GEN_152; // @[playground/src/noop/icache.scala 152:46]
  wire  _GEN_450 = io_instAxi_rd_bits_last ? _GEN_321 : _GEN_153; // @[playground/src/noop/icache.scala 152:46]
  wire  _GEN_451 = io_instAxi_rd_bits_last ? _GEN_322 : _GEN_154; // @[playground/src/noop/icache.scala 152:46]
  wire  _GEN_452 = io_instAxi_rd_bits_last ? _GEN_323 : _GEN_155; // @[playground/src/noop/icache.scala 152:46]
  wire  _GEN_453 = io_instAxi_rd_bits_last ? _GEN_324 : _GEN_156; // @[playground/src/noop/icache.scala 152:46]
  wire  _GEN_454 = io_instAxi_rd_bits_last ? _GEN_325 : _GEN_157; // @[playground/src/noop/icache.scala 152:46]
  wire  _GEN_455 = io_instAxi_rd_bits_last ? _GEN_326 : _GEN_158; // @[playground/src/noop/icache.scala 152:46]
  wire  _GEN_456 = io_instAxi_rd_bits_last ? _GEN_327 : _GEN_159; // @[playground/src/noop/icache.scala 152:46]
  wire  _GEN_457 = io_instAxi_rd_bits_last ? _GEN_328 : _GEN_160; // @[playground/src/noop/icache.scala 152:46]
  wire  _GEN_458 = io_instAxi_rd_bits_last ? _GEN_329 : _GEN_161; // @[playground/src/noop/icache.scala 152:46]
  wire  _GEN_459 = io_instAxi_rd_bits_last ? _GEN_330 : _GEN_162; // @[playground/src/noop/icache.scala 152:46]
  wire  _GEN_460 = io_instAxi_rd_bits_last ? _GEN_331 : _GEN_163; // @[playground/src/noop/icache.scala 152:46]
  wire  _GEN_461 = io_instAxi_rd_bits_last ? _GEN_332 : _GEN_164; // @[playground/src/noop/icache.scala 152:46]
  wire  _GEN_462 = io_instAxi_rd_bits_last ? _GEN_333 : _GEN_165; // @[playground/src/noop/icache.scala 152:46]
  wire  _GEN_463 = io_instAxi_rd_bits_last ? _GEN_334 : _GEN_166; // @[playground/src/noop/icache.scala 152:46]
  wire  _GEN_464 = io_instAxi_rd_bits_last ? _GEN_335 : _GEN_167; // @[playground/src/noop/icache.scala 152:46]
  wire  _GEN_465 = io_instAxi_rd_bits_last ? _GEN_336 : _GEN_168; // @[playground/src/noop/icache.scala 152:46]
  wire  _GEN_466 = io_instAxi_rd_bits_last ? _GEN_337 : _GEN_169; // @[playground/src/noop/icache.scala 152:46]
  wire  _GEN_467 = io_instAxi_rd_bits_last ? _GEN_338 : _GEN_170; // @[playground/src/noop/icache.scala 152:46]
  wire  _GEN_468 = io_instAxi_rd_bits_last ? _GEN_339 : _GEN_171; // @[playground/src/noop/icache.scala 152:46]
  wire  _GEN_469 = io_instAxi_rd_bits_last ? _GEN_340 : _GEN_172; // @[playground/src/noop/icache.scala 152:46]
  wire  _GEN_470 = io_instAxi_rd_bits_last ? _GEN_341 : _GEN_173; // @[playground/src/noop/icache.scala 152:46]
  wire  _GEN_471 = io_instAxi_rd_bits_last ? _GEN_342 : _GEN_174; // @[playground/src/noop/icache.scala 152:46]
  wire  _GEN_472 = io_instAxi_rd_bits_last ? _GEN_343 : _GEN_175; // @[playground/src/noop/icache.scala 152:46]
  wire  _GEN_473 = io_instAxi_rd_bits_last ? _GEN_344 : _GEN_176; // @[playground/src/noop/icache.scala 152:46]
  wire  _GEN_474 = io_instAxi_rd_bits_last ? _GEN_345 : _GEN_177; // @[playground/src/noop/icache.scala 152:46]
  wire  _GEN_475 = io_instAxi_rd_bits_last ? _GEN_346 : _GEN_178; // @[playground/src/noop/icache.scala 152:46]
  wire  _GEN_476 = io_instAxi_rd_bits_last ? _GEN_347 : _GEN_179; // @[playground/src/noop/icache.scala 152:46]
  wire  _GEN_477 = io_instAxi_rd_bits_last ? _GEN_348 : _GEN_180; // @[playground/src/noop/icache.scala 152:46]
  wire  _GEN_478 = io_instAxi_rd_bits_last ? _GEN_349 : _GEN_181; // @[playground/src/noop/icache.scala 152:46]
  wire  _GEN_479 = io_instAxi_rd_bits_last ? _GEN_350 : _GEN_182; // @[playground/src/noop/icache.scala 152:46]
  wire  _GEN_480 = io_instAxi_rd_bits_last ? _GEN_351 : _GEN_183; // @[playground/src/noop/icache.scala 152:46]
  wire  _GEN_481 = io_instAxi_rd_bits_last ? _GEN_352 : _GEN_184; // @[playground/src/noop/icache.scala 152:46]
  wire  _GEN_482 = io_instAxi_rd_bits_last ? _GEN_353 : _GEN_185; // @[playground/src/noop/icache.scala 152:46]
  wire  _GEN_483 = io_instAxi_rd_bits_last ? _GEN_354 : _GEN_186; // @[playground/src/noop/icache.scala 152:46]
  wire  _GEN_484 = io_instAxi_rd_bits_last ? _GEN_355 : _GEN_187; // @[playground/src/noop/icache.scala 152:46]
  wire  _GEN_485 = io_instAxi_rd_bits_last ? _GEN_356 : _GEN_188; // @[playground/src/noop/icache.scala 152:46]
  wire  _GEN_486 = io_instAxi_rd_bits_last ? _GEN_357 : _GEN_189; // @[playground/src/noop/icache.scala 152:46]
  wire  _GEN_487 = io_instAxi_rd_bits_last ? _GEN_358 : _GEN_190; // @[playground/src/noop/icache.scala 152:46]
  wire  _GEN_488 = io_instAxi_rd_bits_last ? _GEN_359 : _GEN_191; // @[playground/src/noop/icache.scala 152:46]
  wire  _GEN_489 = io_instAxi_rd_bits_last ? _GEN_360 : _GEN_192; // @[playground/src/noop/icache.scala 152:46]
  wire  _GEN_490 = io_instAxi_rd_bits_last ? _GEN_361 : _GEN_193; // @[playground/src/noop/icache.scala 152:46]
  wire [1:0] _GEN_491 = io_instAxi_rd_bits_last ? 2'h0 : state; // @[playground/src/noop/icache.scala 102:24 152:46 156:27]
  wire [2:0] _GEN_492 = io_instAxi_rd_bits_last ? 3'h0 : _axiOffset_T_1; // @[playground/src/noop/icache.scala 146:27 152:46 157:31]
  wire [2:0] _GEN_493 = rdataEn & io_instAxi_rd_valid ? _GEN_492 : axiOffset; // @[playground/src/noop/icache.scala 145:49 80:34]
  wire [63:0] _GEN_495 = rdataEn & io_instAxi_rd_valid ? _GEN_233 : databuf; // @[playground/src/noop/icache.scala 145:49 81:34]
  wire  _GEN_496 = rdataEn & io_instAxi_rd_valid ? _GEN_362 : rdataEn; // @[playground/src/noop/icache.scala 119:30 145:49]
  wire [21:0] _GEN_497 = rdataEn & io_instAxi_rd_valid ? _GEN_363 : tag_0_0; // @[playground/src/noop/icache.scala 145:49 65:26]
  wire [21:0] _GEN_498 = rdataEn & io_instAxi_rd_valid ? _GEN_364 : tag_0_1; // @[playground/src/noop/icache.scala 145:49 65:26]
  wire [21:0] _GEN_499 = rdataEn & io_instAxi_rd_valid ? _GEN_365 : tag_0_2; // @[playground/src/noop/icache.scala 145:49 65:26]
  wire [21:0] _GEN_500 = rdataEn & io_instAxi_rd_valid ? _GEN_366 : tag_0_3; // @[playground/src/noop/icache.scala 145:49 65:26]
  wire [21:0] _GEN_501 = rdataEn & io_instAxi_rd_valid ? _GEN_367 : tag_0_4; // @[playground/src/noop/icache.scala 145:49 65:26]
  wire [21:0] _GEN_502 = rdataEn & io_instAxi_rd_valid ? _GEN_368 : tag_0_5; // @[playground/src/noop/icache.scala 145:49 65:26]
  wire [21:0] _GEN_503 = rdataEn & io_instAxi_rd_valid ? _GEN_369 : tag_0_6; // @[playground/src/noop/icache.scala 145:49 65:26]
  wire [21:0] _GEN_504 = rdataEn & io_instAxi_rd_valid ? _GEN_370 : tag_0_7; // @[playground/src/noop/icache.scala 145:49 65:26]
  wire [21:0] _GEN_505 = rdataEn & io_instAxi_rd_valid ? _GEN_371 : tag_0_8; // @[playground/src/noop/icache.scala 145:49 65:26]
  wire [21:0] _GEN_506 = rdataEn & io_instAxi_rd_valid ? _GEN_372 : tag_0_9; // @[playground/src/noop/icache.scala 145:49 65:26]
  wire [21:0] _GEN_507 = rdataEn & io_instAxi_rd_valid ? _GEN_373 : tag_0_10; // @[playground/src/noop/icache.scala 145:49 65:26]
  wire [21:0] _GEN_508 = rdataEn & io_instAxi_rd_valid ? _GEN_374 : tag_0_11; // @[playground/src/noop/icache.scala 145:49 65:26]
  wire [21:0] _GEN_509 = rdataEn & io_instAxi_rd_valid ? _GEN_375 : tag_0_12; // @[playground/src/noop/icache.scala 145:49 65:26]
  wire [21:0] _GEN_510 = rdataEn & io_instAxi_rd_valid ? _GEN_376 : tag_0_13; // @[playground/src/noop/icache.scala 145:49 65:26]
  wire [21:0] _GEN_511 = rdataEn & io_instAxi_rd_valid ? _GEN_377 : tag_0_14; // @[playground/src/noop/icache.scala 145:49 65:26]
  wire [21:0] _GEN_512 = rdataEn & io_instAxi_rd_valid ? _GEN_378 : tag_0_15; // @[playground/src/noop/icache.scala 145:49 65:26]
  wire [21:0] _GEN_513 = rdataEn & io_instAxi_rd_valid ? _GEN_379 : tag_1_0; // @[playground/src/noop/icache.scala 145:49 65:26]
  wire [21:0] _GEN_514 = rdataEn & io_instAxi_rd_valid ? _GEN_380 : tag_1_1; // @[playground/src/noop/icache.scala 145:49 65:26]
  wire [21:0] _GEN_515 = rdataEn & io_instAxi_rd_valid ? _GEN_381 : tag_1_2; // @[playground/src/noop/icache.scala 145:49 65:26]
  wire [21:0] _GEN_516 = rdataEn & io_instAxi_rd_valid ? _GEN_382 : tag_1_3; // @[playground/src/noop/icache.scala 145:49 65:26]
  wire [21:0] _GEN_517 = rdataEn & io_instAxi_rd_valid ? _GEN_383 : tag_1_4; // @[playground/src/noop/icache.scala 145:49 65:26]
  wire [21:0] _GEN_518 = rdataEn & io_instAxi_rd_valid ? _GEN_384 : tag_1_5; // @[playground/src/noop/icache.scala 145:49 65:26]
  wire [21:0] _GEN_519 = rdataEn & io_instAxi_rd_valid ? _GEN_385 : tag_1_6; // @[playground/src/noop/icache.scala 145:49 65:26]
  wire [21:0] _GEN_520 = rdataEn & io_instAxi_rd_valid ? _GEN_386 : tag_1_7; // @[playground/src/noop/icache.scala 145:49 65:26]
  wire [21:0] _GEN_521 = rdataEn & io_instAxi_rd_valid ? _GEN_387 : tag_1_8; // @[playground/src/noop/icache.scala 145:49 65:26]
  wire [21:0] _GEN_522 = rdataEn & io_instAxi_rd_valid ? _GEN_388 : tag_1_9; // @[playground/src/noop/icache.scala 145:49 65:26]
  wire [21:0] _GEN_523 = rdataEn & io_instAxi_rd_valid ? _GEN_389 : tag_1_10; // @[playground/src/noop/icache.scala 145:49 65:26]
  wire [21:0] _GEN_524 = rdataEn & io_instAxi_rd_valid ? _GEN_390 : tag_1_11; // @[playground/src/noop/icache.scala 145:49 65:26]
  wire [21:0] _GEN_525 = rdataEn & io_instAxi_rd_valid ? _GEN_391 : tag_1_12; // @[playground/src/noop/icache.scala 145:49 65:26]
  wire [21:0] _GEN_526 = rdataEn & io_instAxi_rd_valid ? _GEN_392 : tag_1_13; // @[playground/src/noop/icache.scala 145:49 65:26]
  wire [21:0] _GEN_527 = rdataEn & io_instAxi_rd_valid ? _GEN_393 : tag_1_14; // @[playground/src/noop/icache.scala 145:49 65:26]
  wire [21:0] _GEN_528 = rdataEn & io_instAxi_rd_valid ? _GEN_394 : tag_1_15; // @[playground/src/noop/icache.scala 145:49 65:26]
  wire [21:0] _GEN_529 = rdataEn & io_instAxi_rd_valid ? _GEN_395 : tag_2_0; // @[playground/src/noop/icache.scala 145:49 65:26]
  wire [21:0] _GEN_530 = rdataEn & io_instAxi_rd_valid ? _GEN_396 : tag_2_1; // @[playground/src/noop/icache.scala 145:49 65:26]
  wire [21:0] _GEN_531 = rdataEn & io_instAxi_rd_valid ? _GEN_397 : tag_2_2; // @[playground/src/noop/icache.scala 145:49 65:26]
  wire [21:0] _GEN_532 = rdataEn & io_instAxi_rd_valid ? _GEN_398 : tag_2_3; // @[playground/src/noop/icache.scala 145:49 65:26]
  wire [21:0] _GEN_533 = rdataEn & io_instAxi_rd_valid ? _GEN_399 : tag_2_4; // @[playground/src/noop/icache.scala 145:49 65:26]
  wire [21:0] _GEN_534 = rdataEn & io_instAxi_rd_valid ? _GEN_400 : tag_2_5; // @[playground/src/noop/icache.scala 145:49 65:26]
  wire [21:0] _GEN_535 = rdataEn & io_instAxi_rd_valid ? _GEN_401 : tag_2_6; // @[playground/src/noop/icache.scala 145:49 65:26]
  wire [21:0] _GEN_536 = rdataEn & io_instAxi_rd_valid ? _GEN_402 : tag_2_7; // @[playground/src/noop/icache.scala 145:49 65:26]
  wire [21:0] _GEN_537 = rdataEn & io_instAxi_rd_valid ? _GEN_403 : tag_2_8; // @[playground/src/noop/icache.scala 145:49 65:26]
  wire [21:0] _GEN_538 = rdataEn & io_instAxi_rd_valid ? _GEN_404 : tag_2_9; // @[playground/src/noop/icache.scala 145:49 65:26]
  wire [21:0] _GEN_539 = rdataEn & io_instAxi_rd_valid ? _GEN_405 : tag_2_10; // @[playground/src/noop/icache.scala 145:49 65:26]
  wire [21:0] _GEN_540 = rdataEn & io_instAxi_rd_valid ? _GEN_406 : tag_2_11; // @[playground/src/noop/icache.scala 145:49 65:26]
  wire [21:0] _GEN_541 = rdataEn & io_instAxi_rd_valid ? _GEN_407 : tag_2_12; // @[playground/src/noop/icache.scala 145:49 65:26]
  wire [21:0] _GEN_542 = rdataEn & io_instAxi_rd_valid ? _GEN_408 : tag_2_13; // @[playground/src/noop/icache.scala 145:49 65:26]
  wire [21:0] _GEN_543 = rdataEn & io_instAxi_rd_valid ? _GEN_409 : tag_2_14; // @[playground/src/noop/icache.scala 145:49 65:26]
  wire [21:0] _GEN_544 = rdataEn & io_instAxi_rd_valid ? _GEN_410 : tag_2_15; // @[playground/src/noop/icache.scala 145:49 65:26]
  wire [21:0] _GEN_545 = rdataEn & io_instAxi_rd_valid ? _GEN_411 : tag_3_0; // @[playground/src/noop/icache.scala 145:49 65:26]
  wire [21:0] _GEN_546 = rdataEn & io_instAxi_rd_valid ? _GEN_412 : tag_3_1; // @[playground/src/noop/icache.scala 145:49 65:26]
  wire [21:0] _GEN_547 = rdataEn & io_instAxi_rd_valid ? _GEN_413 : tag_3_2; // @[playground/src/noop/icache.scala 145:49 65:26]
  wire [21:0] _GEN_548 = rdataEn & io_instAxi_rd_valid ? _GEN_414 : tag_3_3; // @[playground/src/noop/icache.scala 145:49 65:26]
  wire [21:0] _GEN_549 = rdataEn & io_instAxi_rd_valid ? _GEN_415 : tag_3_4; // @[playground/src/noop/icache.scala 145:49 65:26]
  wire [21:0] _GEN_550 = rdataEn & io_instAxi_rd_valid ? _GEN_416 : tag_3_5; // @[playground/src/noop/icache.scala 145:49 65:26]
  wire [21:0] _GEN_551 = rdataEn & io_instAxi_rd_valid ? _GEN_417 : tag_3_6; // @[playground/src/noop/icache.scala 145:49 65:26]
  wire [21:0] _GEN_552 = rdataEn & io_instAxi_rd_valid ? _GEN_418 : tag_3_7; // @[playground/src/noop/icache.scala 145:49 65:26]
  wire [21:0] _GEN_553 = rdataEn & io_instAxi_rd_valid ? _GEN_419 : tag_3_8; // @[playground/src/noop/icache.scala 145:49 65:26]
  wire [21:0] _GEN_554 = rdataEn & io_instAxi_rd_valid ? _GEN_420 : tag_3_9; // @[playground/src/noop/icache.scala 145:49 65:26]
  wire [21:0] _GEN_555 = rdataEn & io_instAxi_rd_valid ? _GEN_421 : tag_3_10; // @[playground/src/noop/icache.scala 145:49 65:26]
  wire [21:0] _GEN_556 = rdataEn & io_instAxi_rd_valid ? _GEN_422 : tag_3_11; // @[playground/src/noop/icache.scala 145:49 65:26]
  wire [21:0] _GEN_557 = rdataEn & io_instAxi_rd_valid ? _GEN_423 : tag_3_12; // @[playground/src/noop/icache.scala 145:49 65:26]
  wire [21:0] _GEN_558 = rdataEn & io_instAxi_rd_valid ? _GEN_424 : tag_3_13; // @[playground/src/noop/icache.scala 145:49 65:26]
  wire [21:0] _GEN_559 = rdataEn & io_instAxi_rd_valid ? _GEN_425 : tag_3_14; // @[playground/src/noop/icache.scala 145:49 65:26]
  wire [21:0] _GEN_560 = rdataEn & io_instAxi_rd_valid ? _GEN_426 : tag_3_15; // @[playground/src/noop/icache.scala 145:49 65:26]
  wire  _GEN_561 = rdataEn & io_instAxi_rd_valid ? _GEN_427 : _GEN_130; // @[playground/src/noop/icache.scala 145:49]
  wire  _GEN_562 = rdataEn & io_instAxi_rd_valid ? _GEN_428 : _GEN_131; // @[playground/src/noop/icache.scala 145:49]
  wire  _GEN_563 = rdataEn & io_instAxi_rd_valid ? _GEN_429 : _GEN_132; // @[playground/src/noop/icache.scala 145:49]
  wire  _GEN_564 = rdataEn & io_instAxi_rd_valid ? _GEN_430 : _GEN_133; // @[playground/src/noop/icache.scala 145:49]
  wire  _GEN_565 = rdataEn & io_instAxi_rd_valid ? _GEN_431 : _GEN_134; // @[playground/src/noop/icache.scala 145:49]
  wire  _GEN_566 = rdataEn & io_instAxi_rd_valid ? _GEN_432 : _GEN_135; // @[playground/src/noop/icache.scala 145:49]
  wire  _GEN_567 = rdataEn & io_instAxi_rd_valid ? _GEN_433 : _GEN_136; // @[playground/src/noop/icache.scala 145:49]
  wire  _GEN_568 = rdataEn & io_instAxi_rd_valid ? _GEN_434 : _GEN_137; // @[playground/src/noop/icache.scala 145:49]
  wire  _GEN_569 = rdataEn & io_instAxi_rd_valid ? _GEN_435 : _GEN_138; // @[playground/src/noop/icache.scala 145:49]
  wire  _GEN_570 = rdataEn & io_instAxi_rd_valid ? _GEN_436 : _GEN_139; // @[playground/src/noop/icache.scala 145:49]
  wire  _GEN_571 = rdataEn & io_instAxi_rd_valid ? _GEN_437 : _GEN_140; // @[playground/src/noop/icache.scala 145:49]
  wire  _GEN_572 = rdataEn & io_instAxi_rd_valid ? _GEN_438 : _GEN_141; // @[playground/src/noop/icache.scala 145:49]
  wire  _GEN_573 = rdataEn & io_instAxi_rd_valid ? _GEN_439 : _GEN_142; // @[playground/src/noop/icache.scala 145:49]
  wire  _GEN_574 = rdataEn & io_instAxi_rd_valid ? _GEN_440 : _GEN_143; // @[playground/src/noop/icache.scala 145:49]
  wire  _GEN_575 = rdataEn & io_instAxi_rd_valid ? _GEN_441 : _GEN_144; // @[playground/src/noop/icache.scala 145:49]
  wire  _GEN_576 = rdataEn & io_instAxi_rd_valid ? _GEN_442 : _GEN_145; // @[playground/src/noop/icache.scala 145:49]
  wire  _GEN_577 = rdataEn & io_instAxi_rd_valid ? _GEN_443 : _GEN_146; // @[playground/src/noop/icache.scala 145:49]
  wire  _GEN_578 = rdataEn & io_instAxi_rd_valid ? _GEN_444 : _GEN_147; // @[playground/src/noop/icache.scala 145:49]
  wire  _GEN_579 = rdataEn & io_instAxi_rd_valid ? _GEN_445 : _GEN_148; // @[playground/src/noop/icache.scala 145:49]
  wire  _GEN_580 = rdataEn & io_instAxi_rd_valid ? _GEN_446 : _GEN_149; // @[playground/src/noop/icache.scala 145:49]
  wire  _GEN_581 = rdataEn & io_instAxi_rd_valid ? _GEN_447 : _GEN_150; // @[playground/src/noop/icache.scala 145:49]
  wire  _GEN_582 = rdataEn & io_instAxi_rd_valid ? _GEN_448 : _GEN_151; // @[playground/src/noop/icache.scala 145:49]
  wire  _GEN_583 = rdataEn & io_instAxi_rd_valid ? _GEN_449 : _GEN_152; // @[playground/src/noop/icache.scala 145:49]
  wire  _GEN_584 = rdataEn & io_instAxi_rd_valid ? _GEN_450 : _GEN_153; // @[playground/src/noop/icache.scala 145:49]
  wire  _GEN_585 = rdataEn & io_instAxi_rd_valid ? _GEN_451 : _GEN_154; // @[playground/src/noop/icache.scala 145:49]
  wire  _GEN_586 = rdataEn & io_instAxi_rd_valid ? _GEN_452 : _GEN_155; // @[playground/src/noop/icache.scala 145:49]
  wire  _GEN_587 = rdataEn & io_instAxi_rd_valid ? _GEN_453 : _GEN_156; // @[playground/src/noop/icache.scala 145:49]
  wire  _GEN_588 = rdataEn & io_instAxi_rd_valid ? _GEN_454 : _GEN_157; // @[playground/src/noop/icache.scala 145:49]
  wire  _GEN_589 = rdataEn & io_instAxi_rd_valid ? _GEN_455 : _GEN_158; // @[playground/src/noop/icache.scala 145:49]
  wire  _GEN_590 = rdataEn & io_instAxi_rd_valid ? _GEN_456 : _GEN_159; // @[playground/src/noop/icache.scala 145:49]
  wire  _GEN_591 = rdataEn & io_instAxi_rd_valid ? _GEN_457 : _GEN_160; // @[playground/src/noop/icache.scala 145:49]
  wire  _GEN_592 = rdataEn & io_instAxi_rd_valid ? _GEN_458 : _GEN_161; // @[playground/src/noop/icache.scala 145:49]
  wire  _GEN_593 = rdataEn & io_instAxi_rd_valid ? _GEN_459 : _GEN_162; // @[playground/src/noop/icache.scala 145:49]
  wire  _GEN_594 = rdataEn & io_instAxi_rd_valid ? _GEN_460 : _GEN_163; // @[playground/src/noop/icache.scala 145:49]
  wire  _GEN_595 = rdataEn & io_instAxi_rd_valid ? _GEN_461 : _GEN_164; // @[playground/src/noop/icache.scala 145:49]
  wire  _GEN_596 = rdataEn & io_instAxi_rd_valid ? _GEN_462 : _GEN_165; // @[playground/src/noop/icache.scala 145:49]
  wire  _GEN_597 = rdataEn & io_instAxi_rd_valid ? _GEN_463 : _GEN_166; // @[playground/src/noop/icache.scala 145:49]
  wire  _GEN_598 = rdataEn & io_instAxi_rd_valid ? _GEN_464 : _GEN_167; // @[playground/src/noop/icache.scala 145:49]
  wire  _GEN_599 = rdataEn & io_instAxi_rd_valid ? _GEN_465 : _GEN_168; // @[playground/src/noop/icache.scala 145:49]
  wire  _GEN_600 = rdataEn & io_instAxi_rd_valid ? _GEN_466 : _GEN_169; // @[playground/src/noop/icache.scala 145:49]
  wire  _GEN_601 = rdataEn & io_instAxi_rd_valid ? _GEN_467 : _GEN_170; // @[playground/src/noop/icache.scala 145:49]
  wire  _GEN_602 = rdataEn & io_instAxi_rd_valid ? _GEN_468 : _GEN_171; // @[playground/src/noop/icache.scala 145:49]
  wire  _GEN_603 = rdataEn & io_instAxi_rd_valid ? _GEN_469 : _GEN_172; // @[playground/src/noop/icache.scala 145:49]
  wire  _GEN_604 = rdataEn & io_instAxi_rd_valid ? _GEN_470 : _GEN_173; // @[playground/src/noop/icache.scala 145:49]
  wire  _GEN_605 = rdataEn & io_instAxi_rd_valid ? _GEN_471 : _GEN_174; // @[playground/src/noop/icache.scala 145:49]
  wire  _GEN_606 = rdataEn & io_instAxi_rd_valid ? _GEN_472 : _GEN_175; // @[playground/src/noop/icache.scala 145:49]
  wire  _GEN_607 = rdataEn & io_instAxi_rd_valid ? _GEN_473 : _GEN_176; // @[playground/src/noop/icache.scala 145:49]
  wire  _GEN_608 = rdataEn & io_instAxi_rd_valid ? _GEN_474 : _GEN_177; // @[playground/src/noop/icache.scala 145:49]
  wire  _GEN_609 = rdataEn & io_instAxi_rd_valid ? _GEN_475 : _GEN_178; // @[playground/src/noop/icache.scala 145:49]
  wire  _GEN_610 = rdataEn & io_instAxi_rd_valid ? _GEN_476 : _GEN_179; // @[playground/src/noop/icache.scala 145:49]
  wire  _GEN_611 = rdataEn & io_instAxi_rd_valid ? _GEN_477 : _GEN_180; // @[playground/src/noop/icache.scala 145:49]
  wire  _GEN_612 = rdataEn & io_instAxi_rd_valid ? _GEN_478 : _GEN_181; // @[playground/src/noop/icache.scala 145:49]
  wire  _GEN_613 = rdataEn & io_instAxi_rd_valid ? _GEN_479 : _GEN_182; // @[playground/src/noop/icache.scala 145:49]
  wire  _GEN_614 = rdataEn & io_instAxi_rd_valid ? _GEN_480 : _GEN_183; // @[playground/src/noop/icache.scala 145:49]
  wire  _GEN_615 = rdataEn & io_instAxi_rd_valid ? _GEN_481 : _GEN_184; // @[playground/src/noop/icache.scala 145:49]
  wire  _GEN_616 = rdataEn & io_instAxi_rd_valid ? _GEN_482 : _GEN_185; // @[playground/src/noop/icache.scala 145:49]
  wire  _GEN_617 = rdataEn & io_instAxi_rd_valid ? _GEN_483 : _GEN_186; // @[playground/src/noop/icache.scala 145:49]
  wire  _GEN_618 = rdataEn & io_instAxi_rd_valid ? _GEN_484 : _GEN_187; // @[playground/src/noop/icache.scala 145:49]
  wire  _GEN_619 = rdataEn & io_instAxi_rd_valid ? _GEN_485 : _GEN_188; // @[playground/src/noop/icache.scala 145:49]
  wire  _GEN_620 = rdataEn & io_instAxi_rd_valid ? _GEN_486 : _GEN_189; // @[playground/src/noop/icache.scala 145:49]
  wire  _GEN_621 = rdataEn & io_instAxi_rd_valid ? _GEN_487 : _GEN_190; // @[playground/src/noop/icache.scala 145:49]
  wire  _GEN_622 = rdataEn & io_instAxi_rd_valid ? _GEN_488 : _GEN_191; // @[playground/src/noop/icache.scala 145:49]
  wire  _GEN_623 = rdataEn & io_instAxi_rd_valid ? _GEN_489 : _GEN_192; // @[playground/src/noop/icache.scala 145:49]
  wire  _GEN_624 = rdataEn & io_instAxi_rd_valid ? _GEN_490 : _GEN_193; // @[playground/src/noop/icache.scala 145:49]
  wire [1:0] _GEN_625 = rdataEn & io_instAxi_rd_valid ? _GEN_491 : state; // @[playground/src/noop/icache.scala 102:24 145:49]
  wire  _GEN_893 = 2'h0 == state & _GEN_223; // @[playground/src/noop/icache.scala 121:18 73:13]
  Ram_bw Ram_bw ( // @[playground/src/noop/icache.scala 67:57]
    .clock(Ram_bw_clock),
    .reset(Ram_bw_reset),
    .io_cen(Ram_bw_io_cen),
    .io_wen(Ram_bw_io_wen),
    .io_addr(Ram_bw_io_addr),
    .io_rdata(Ram_bw_io_rdata),
    .io_wdata(Ram_bw_io_wdata),
    .io_mask(Ram_bw_io_mask)
  );
  Ram_bw Ram_bw_1 ( // @[playground/src/noop/icache.scala 67:57]
    .clock(Ram_bw_1_clock),
    .reset(Ram_bw_1_reset),
    .io_cen(Ram_bw_1_io_cen),
    .io_wen(Ram_bw_1_io_wen),
    .io_addr(Ram_bw_1_io_addr),
    .io_rdata(Ram_bw_1_io_rdata),
    .io_wdata(Ram_bw_1_io_wdata),
    .io_mask(Ram_bw_1_io_mask)
  );
  Ram_bw Ram_bw_2 ( // @[playground/src/noop/icache.scala 67:57]
    .clock(Ram_bw_2_clock),
    .reset(Ram_bw_2_reset),
    .io_cen(Ram_bw_2_io_cen),
    .io_wen(Ram_bw_2_io_wen),
    .io_addr(Ram_bw_2_io_addr),
    .io_rdata(Ram_bw_2_io_rdata),
    .io_wdata(Ram_bw_2_io_wdata),
    .io_mask(Ram_bw_2_io_mask)
  );
  Ram_bw Ram_bw_3 ( // @[playground/src/noop/icache.scala 67:57]
    .clock(Ram_bw_3_clock),
    .reset(Ram_bw_3_reset),
    .io_cen(Ram_bw_3_io_cen),
    .io_wen(Ram_bw_3_io_wen),
    .io_addr(Ram_bw_3_io_addr),
    .io_rdata(Ram_bw_3_io_rdata),
    .io_wdata(Ram_bw_3_io_wdata),
    .io_mask(Ram_bw_3_io_mask)
  );
  MaxPeriodFibonacciLFSR matchWay_prng ( // @[src/main/scala/chisel3/util/random/PRNG.scala 91:22]
    .clock(matchWay_prng_clock),
    .reset(matchWay_prng_reset),
    .io_out_0(matchWay_prng_io_out_0),
    .io_out_1(matchWay_prng_io_out_1)
  );
  assign io_instAxi_ra_valid = raddrEn; // @[playground/src/noop/icache.scala 165:30]
  assign io_instAxi_ra_bits_addr = raddr; // @[playground/src/noop/icache.scala 166:30]
  assign io_icRead_inst = addr_r[3] ? _GEN_197[127:64] : _GEN_197[63:0]; // @[src/main/scala/chisel3/util/Mux.scala 81:58]
  assign io_icRead_ready = valid_in & ~wait_r; // @[playground/src/noop/icache.scala 76:37]
  assign io_icRead_rvalid = valid_r; // @[playground/src/noop/icache.scala 77:25]
  assign Ram_bw_clock = clock;
  assign Ram_bw_reset = reset;
  assign Ram_bw_io_cen = 2'h0 == cur_way[1:0] & (wait_r | hs_in); // @[playground/src/noop/icache.scala 111:{25,25} playground/src/ram/ram.scala 41:17]
  assign Ram_bw_io_wen = _GEN_1030 & wen; // @[playground/src/noop/icache.scala 112:{25,25} playground/src/ram/ram.scala 42:17]
  assign Ram_bw_io_addr = 2'h0 == cur_way[1:0] ? _data_addr_T_1 : 6'h0; // @[playground/src/noop/icache.scala 110:{25,25} playground/src/ram/ram.scala 43:17]
  assign Ram_bw_io_wdata = 2'h0 == cur_way[1:0] ? _data_wdata_T : 128'h0; // @[playground/src/noop/icache.scala 113:{25,25} playground/src/ram/ram.scala 44:17]
  assign Ram_bw_io_mask = 2'h0 == cur_way[1:0] ? 128'hffffffffffffffffffffffffffffffff : 128'h0; // @[playground/src/noop/icache.scala 114:{25,25} playground/src/ram/ram.scala 45:17]
  assign Ram_bw_1_clock = clock;
  assign Ram_bw_1_reset = reset;
  assign Ram_bw_1_io_cen = 2'h1 == cur_way[1:0] & (wait_r | hs_in); // @[playground/src/noop/icache.scala 111:{25,25} playground/src/ram/ram.scala 41:17]
  assign Ram_bw_1_io_wen = _GEN_1031 & wen; // @[playground/src/noop/icache.scala 112:{25,25} playground/src/ram/ram.scala 42:17]
  assign Ram_bw_1_io_addr = 2'h1 == cur_way[1:0] ? _data_addr_T_1 : 6'h0; // @[playground/src/noop/icache.scala 110:{25,25} playground/src/ram/ram.scala 43:17]
  assign Ram_bw_1_io_wdata = 2'h1 == cur_way[1:0] ? _data_wdata_T : 128'h0; // @[playground/src/noop/icache.scala 113:{25,25} playground/src/ram/ram.scala 44:17]
  assign Ram_bw_1_io_mask = 2'h1 == cur_way[1:0] ? 128'hffffffffffffffffffffffffffffffff : 128'h0; // @[playground/src/noop/icache.scala 114:{25,25} playground/src/ram/ram.scala 45:17]
  assign Ram_bw_2_clock = clock;
  assign Ram_bw_2_reset = reset;
  assign Ram_bw_2_io_cen = 2'h2 == cur_way[1:0] & (wait_r | hs_in); // @[playground/src/noop/icache.scala 111:{25,25} playground/src/ram/ram.scala 41:17]
  assign Ram_bw_2_io_wen = _GEN_1032 & wen; // @[playground/src/noop/icache.scala 112:{25,25} playground/src/ram/ram.scala 42:17]
  assign Ram_bw_2_io_addr = 2'h2 == cur_way[1:0] ? _data_addr_T_1 : 6'h0; // @[playground/src/noop/icache.scala 110:{25,25} playground/src/ram/ram.scala 43:17]
  assign Ram_bw_2_io_wdata = 2'h2 == cur_way[1:0] ? _data_wdata_T : 128'h0; // @[playground/src/noop/icache.scala 113:{25,25} playground/src/ram/ram.scala 44:17]
  assign Ram_bw_2_io_mask = 2'h2 == cur_way[1:0] ? 128'hffffffffffffffffffffffffffffffff : 128'h0; // @[playground/src/noop/icache.scala 114:{25,25} playground/src/ram/ram.scala 45:17]
  assign Ram_bw_3_clock = clock;
  assign Ram_bw_3_reset = reset;
  assign Ram_bw_3_io_cen = 2'h3 == cur_way[1:0] & (wait_r | hs_in); // @[playground/src/noop/icache.scala 111:{25,25} playground/src/ram/ram.scala 41:17]
  assign Ram_bw_3_io_wen = _GEN_1033 & wen; // @[playground/src/noop/icache.scala 112:{25,25} playground/src/ram/ram.scala 42:17]
  assign Ram_bw_3_io_addr = 2'h3 == cur_way[1:0] ? _data_addr_T_1 : 6'h0; // @[playground/src/noop/icache.scala 110:{25,25} playground/src/ram/ram.scala 43:17]
  assign Ram_bw_3_io_wdata = 2'h3 == cur_way[1:0] ? _data_wdata_T : 128'h0; // @[playground/src/noop/icache.scala 113:{25,25} playground/src/ram/ram.scala 44:17]
  assign Ram_bw_3_io_mask = 2'h3 == cur_way[1:0] ? 128'hffffffffffffffffffffffffffffffff : 128'h0; // @[playground/src/noop/icache.scala 114:{25,25} playground/src/ram/ram.scala 45:17]
  assign matchWay_prng_clock = clock;
  assign matchWay_prng_reset = reset;
  always @(posedge clock) begin
    if (reset) begin // @[playground/src/noop/icache.scala 65:26]
      tag_0_0 <= 22'h0; // @[playground/src/noop/icache.scala 65:26]
    end else if (!(2'h0 == state)) begin // @[playground/src/noop/icache.scala 121:18]
      if (!(2'h1 == state)) begin // @[playground/src/noop/icache.scala 121:18]
        if (2'h2 == state) begin // @[playground/src/noop/icache.scala 121:18]
          tag_0_0 <= _GEN_497;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/icache.scala 65:26]
      tag_0_1 <= 22'h0; // @[playground/src/noop/icache.scala 65:26]
    end else if (!(2'h0 == state)) begin // @[playground/src/noop/icache.scala 121:18]
      if (!(2'h1 == state)) begin // @[playground/src/noop/icache.scala 121:18]
        if (2'h2 == state) begin // @[playground/src/noop/icache.scala 121:18]
          tag_0_1 <= _GEN_498;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/icache.scala 65:26]
      tag_0_2 <= 22'h0; // @[playground/src/noop/icache.scala 65:26]
    end else if (!(2'h0 == state)) begin // @[playground/src/noop/icache.scala 121:18]
      if (!(2'h1 == state)) begin // @[playground/src/noop/icache.scala 121:18]
        if (2'h2 == state) begin // @[playground/src/noop/icache.scala 121:18]
          tag_0_2 <= _GEN_499;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/icache.scala 65:26]
      tag_0_3 <= 22'h0; // @[playground/src/noop/icache.scala 65:26]
    end else if (!(2'h0 == state)) begin // @[playground/src/noop/icache.scala 121:18]
      if (!(2'h1 == state)) begin // @[playground/src/noop/icache.scala 121:18]
        if (2'h2 == state) begin // @[playground/src/noop/icache.scala 121:18]
          tag_0_3 <= _GEN_500;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/icache.scala 65:26]
      tag_0_4 <= 22'h0; // @[playground/src/noop/icache.scala 65:26]
    end else if (!(2'h0 == state)) begin // @[playground/src/noop/icache.scala 121:18]
      if (!(2'h1 == state)) begin // @[playground/src/noop/icache.scala 121:18]
        if (2'h2 == state) begin // @[playground/src/noop/icache.scala 121:18]
          tag_0_4 <= _GEN_501;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/icache.scala 65:26]
      tag_0_5 <= 22'h0; // @[playground/src/noop/icache.scala 65:26]
    end else if (!(2'h0 == state)) begin // @[playground/src/noop/icache.scala 121:18]
      if (!(2'h1 == state)) begin // @[playground/src/noop/icache.scala 121:18]
        if (2'h2 == state) begin // @[playground/src/noop/icache.scala 121:18]
          tag_0_5 <= _GEN_502;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/icache.scala 65:26]
      tag_0_6 <= 22'h0; // @[playground/src/noop/icache.scala 65:26]
    end else if (!(2'h0 == state)) begin // @[playground/src/noop/icache.scala 121:18]
      if (!(2'h1 == state)) begin // @[playground/src/noop/icache.scala 121:18]
        if (2'h2 == state) begin // @[playground/src/noop/icache.scala 121:18]
          tag_0_6 <= _GEN_503;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/icache.scala 65:26]
      tag_0_7 <= 22'h0; // @[playground/src/noop/icache.scala 65:26]
    end else if (!(2'h0 == state)) begin // @[playground/src/noop/icache.scala 121:18]
      if (!(2'h1 == state)) begin // @[playground/src/noop/icache.scala 121:18]
        if (2'h2 == state) begin // @[playground/src/noop/icache.scala 121:18]
          tag_0_7 <= _GEN_504;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/icache.scala 65:26]
      tag_0_8 <= 22'h0; // @[playground/src/noop/icache.scala 65:26]
    end else if (!(2'h0 == state)) begin // @[playground/src/noop/icache.scala 121:18]
      if (!(2'h1 == state)) begin // @[playground/src/noop/icache.scala 121:18]
        if (2'h2 == state) begin // @[playground/src/noop/icache.scala 121:18]
          tag_0_8 <= _GEN_505;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/icache.scala 65:26]
      tag_0_9 <= 22'h0; // @[playground/src/noop/icache.scala 65:26]
    end else if (!(2'h0 == state)) begin // @[playground/src/noop/icache.scala 121:18]
      if (!(2'h1 == state)) begin // @[playground/src/noop/icache.scala 121:18]
        if (2'h2 == state) begin // @[playground/src/noop/icache.scala 121:18]
          tag_0_9 <= _GEN_506;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/icache.scala 65:26]
      tag_0_10 <= 22'h0; // @[playground/src/noop/icache.scala 65:26]
    end else if (!(2'h0 == state)) begin // @[playground/src/noop/icache.scala 121:18]
      if (!(2'h1 == state)) begin // @[playground/src/noop/icache.scala 121:18]
        if (2'h2 == state) begin // @[playground/src/noop/icache.scala 121:18]
          tag_0_10 <= _GEN_507;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/icache.scala 65:26]
      tag_0_11 <= 22'h0; // @[playground/src/noop/icache.scala 65:26]
    end else if (!(2'h0 == state)) begin // @[playground/src/noop/icache.scala 121:18]
      if (!(2'h1 == state)) begin // @[playground/src/noop/icache.scala 121:18]
        if (2'h2 == state) begin // @[playground/src/noop/icache.scala 121:18]
          tag_0_11 <= _GEN_508;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/icache.scala 65:26]
      tag_0_12 <= 22'h0; // @[playground/src/noop/icache.scala 65:26]
    end else if (!(2'h0 == state)) begin // @[playground/src/noop/icache.scala 121:18]
      if (!(2'h1 == state)) begin // @[playground/src/noop/icache.scala 121:18]
        if (2'h2 == state) begin // @[playground/src/noop/icache.scala 121:18]
          tag_0_12 <= _GEN_509;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/icache.scala 65:26]
      tag_0_13 <= 22'h0; // @[playground/src/noop/icache.scala 65:26]
    end else if (!(2'h0 == state)) begin // @[playground/src/noop/icache.scala 121:18]
      if (!(2'h1 == state)) begin // @[playground/src/noop/icache.scala 121:18]
        if (2'h2 == state) begin // @[playground/src/noop/icache.scala 121:18]
          tag_0_13 <= _GEN_510;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/icache.scala 65:26]
      tag_0_14 <= 22'h0; // @[playground/src/noop/icache.scala 65:26]
    end else if (!(2'h0 == state)) begin // @[playground/src/noop/icache.scala 121:18]
      if (!(2'h1 == state)) begin // @[playground/src/noop/icache.scala 121:18]
        if (2'h2 == state) begin // @[playground/src/noop/icache.scala 121:18]
          tag_0_14 <= _GEN_511;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/icache.scala 65:26]
      tag_0_15 <= 22'h0; // @[playground/src/noop/icache.scala 65:26]
    end else if (!(2'h0 == state)) begin // @[playground/src/noop/icache.scala 121:18]
      if (!(2'h1 == state)) begin // @[playground/src/noop/icache.scala 121:18]
        if (2'h2 == state) begin // @[playground/src/noop/icache.scala 121:18]
          tag_0_15 <= _GEN_512;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/icache.scala 65:26]
      tag_1_0 <= 22'h0; // @[playground/src/noop/icache.scala 65:26]
    end else if (!(2'h0 == state)) begin // @[playground/src/noop/icache.scala 121:18]
      if (!(2'h1 == state)) begin // @[playground/src/noop/icache.scala 121:18]
        if (2'h2 == state) begin // @[playground/src/noop/icache.scala 121:18]
          tag_1_0 <= _GEN_513;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/icache.scala 65:26]
      tag_1_1 <= 22'h0; // @[playground/src/noop/icache.scala 65:26]
    end else if (!(2'h0 == state)) begin // @[playground/src/noop/icache.scala 121:18]
      if (!(2'h1 == state)) begin // @[playground/src/noop/icache.scala 121:18]
        if (2'h2 == state) begin // @[playground/src/noop/icache.scala 121:18]
          tag_1_1 <= _GEN_514;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/icache.scala 65:26]
      tag_1_2 <= 22'h0; // @[playground/src/noop/icache.scala 65:26]
    end else if (!(2'h0 == state)) begin // @[playground/src/noop/icache.scala 121:18]
      if (!(2'h1 == state)) begin // @[playground/src/noop/icache.scala 121:18]
        if (2'h2 == state) begin // @[playground/src/noop/icache.scala 121:18]
          tag_1_2 <= _GEN_515;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/icache.scala 65:26]
      tag_1_3 <= 22'h0; // @[playground/src/noop/icache.scala 65:26]
    end else if (!(2'h0 == state)) begin // @[playground/src/noop/icache.scala 121:18]
      if (!(2'h1 == state)) begin // @[playground/src/noop/icache.scala 121:18]
        if (2'h2 == state) begin // @[playground/src/noop/icache.scala 121:18]
          tag_1_3 <= _GEN_516;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/icache.scala 65:26]
      tag_1_4 <= 22'h0; // @[playground/src/noop/icache.scala 65:26]
    end else if (!(2'h0 == state)) begin // @[playground/src/noop/icache.scala 121:18]
      if (!(2'h1 == state)) begin // @[playground/src/noop/icache.scala 121:18]
        if (2'h2 == state) begin // @[playground/src/noop/icache.scala 121:18]
          tag_1_4 <= _GEN_517;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/icache.scala 65:26]
      tag_1_5 <= 22'h0; // @[playground/src/noop/icache.scala 65:26]
    end else if (!(2'h0 == state)) begin // @[playground/src/noop/icache.scala 121:18]
      if (!(2'h1 == state)) begin // @[playground/src/noop/icache.scala 121:18]
        if (2'h2 == state) begin // @[playground/src/noop/icache.scala 121:18]
          tag_1_5 <= _GEN_518;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/icache.scala 65:26]
      tag_1_6 <= 22'h0; // @[playground/src/noop/icache.scala 65:26]
    end else if (!(2'h0 == state)) begin // @[playground/src/noop/icache.scala 121:18]
      if (!(2'h1 == state)) begin // @[playground/src/noop/icache.scala 121:18]
        if (2'h2 == state) begin // @[playground/src/noop/icache.scala 121:18]
          tag_1_6 <= _GEN_519;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/icache.scala 65:26]
      tag_1_7 <= 22'h0; // @[playground/src/noop/icache.scala 65:26]
    end else if (!(2'h0 == state)) begin // @[playground/src/noop/icache.scala 121:18]
      if (!(2'h1 == state)) begin // @[playground/src/noop/icache.scala 121:18]
        if (2'h2 == state) begin // @[playground/src/noop/icache.scala 121:18]
          tag_1_7 <= _GEN_520;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/icache.scala 65:26]
      tag_1_8 <= 22'h0; // @[playground/src/noop/icache.scala 65:26]
    end else if (!(2'h0 == state)) begin // @[playground/src/noop/icache.scala 121:18]
      if (!(2'h1 == state)) begin // @[playground/src/noop/icache.scala 121:18]
        if (2'h2 == state) begin // @[playground/src/noop/icache.scala 121:18]
          tag_1_8 <= _GEN_521;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/icache.scala 65:26]
      tag_1_9 <= 22'h0; // @[playground/src/noop/icache.scala 65:26]
    end else if (!(2'h0 == state)) begin // @[playground/src/noop/icache.scala 121:18]
      if (!(2'h1 == state)) begin // @[playground/src/noop/icache.scala 121:18]
        if (2'h2 == state) begin // @[playground/src/noop/icache.scala 121:18]
          tag_1_9 <= _GEN_522;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/icache.scala 65:26]
      tag_1_10 <= 22'h0; // @[playground/src/noop/icache.scala 65:26]
    end else if (!(2'h0 == state)) begin // @[playground/src/noop/icache.scala 121:18]
      if (!(2'h1 == state)) begin // @[playground/src/noop/icache.scala 121:18]
        if (2'h2 == state) begin // @[playground/src/noop/icache.scala 121:18]
          tag_1_10 <= _GEN_523;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/icache.scala 65:26]
      tag_1_11 <= 22'h0; // @[playground/src/noop/icache.scala 65:26]
    end else if (!(2'h0 == state)) begin // @[playground/src/noop/icache.scala 121:18]
      if (!(2'h1 == state)) begin // @[playground/src/noop/icache.scala 121:18]
        if (2'h2 == state) begin // @[playground/src/noop/icache.scala 121:18]
          tag_1_11 <= _GEN_524;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/icache.scala 65:26]
      tag_1_12 <= 22'h0; // @[playground/src/noop/icache.scala 65:26]
    end else if (!(2'h0 == state)) begin // @[playground/src/noop/icache.scala 121:18]
      if (!(2'h1 == state)) begin // @[playground/src/noop/icache.scala 121:18]
        if (2'h2 == state) begin // @[playground/src/noop/icache.scala 121:18]
          tag_1_12 <= _GEN_525;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/icache.scala 65:26]
      tag_1_13 <= 22'h0; // @[playground/src/noop/icache.scala 65:26]
    end else if (!(2'h0 == state)) begin // @[playground/src/noop/icache.scala 121:18]
      if (!(2'h1 == state)) begin // @[playground/src/noop/icache.scala 121:18]
        if (2'h2 == state) begin // @[playground/src/noop/icache.scala 121:18]
          tag_1_13 <= _GEN_526;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/icache.scala 65:26]
      tag_1_14 <= 22'h0; // @[playground/src/noop/icache.scala 65:26]
    end else if (!(2'h0 == state)) begin // @[playground/src/noop/icache.scala 121:18]
      if (!(2'h1 == state)) begin // @[playground/src/noop/icache.scala 121:18]
        if (2'h2 == state) begin // @[playground/src/noop/icache.scala 121:18]
          tag_1_14 <= _GEN_527;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/icache.scala 65:26]
      tag_1_15 <= 22'h0; // @[playground/src/noop/icache.scala 65:26]
    end else if (!(2'h0 == state)) begin // @[playground/src/noop/icache.scala 121:18]
      if (!(2'h1 == state)) begin // @[playground/src/noop/icache.scala 121:18]
        if (2'h2 == state) begin // @[playground/src/noop/icache.scala 121:18]
          tag_1_15 <= _GEN_528;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/icache.scala 65:26]
      tag_2_0 <= 22'h0; // @[playground/src/noop/icache.scala 65:26]
    end else if (!(2'h0 == state)) begin // @[playground/src/noop/icache.scala 121:18]
      if (!(2'h1 == state)) begin // @[playground/src/noop/icache.scala 121:18]
        if (2'h2 == state) begin // @[playground/src/noop/icache.scala 121:18]
          tag_2_0 <= _GEN_529;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/icache.scala 65:26]
      tag_2_1 <= 22'h0; // @[playground/src/noop/icache.scala 65:26]
    end else if (!(2'h0 == state)) begin // @[playground/src/noop/icache.scala 121:18]
      if (!(2'h1 == state)) begin // @[playground/src/noop/icache.scala 121:18]
        if (2'h2 == state) begin // @[playground/src/noop/icache.scala 121:18]
          tag_2_1 <= _GEN_530;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/icache.scala 65:26]
      tag_2_2 <= 22'h0; // @[playground/src/noop/icache.scala 65:26]
    end else if (!(2'h0 == state)) begin // @[playground/src/noop/icache.scala 121:18]
      if (!(2'h1 == state)) begin // @[playground/src/noop/icache.scala 121:18]
        if (2'h2 == state) begin // @[playground/src/noop/icache.scala 121:18]
          tag_2_2 <= _GEN_531;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/icache.scala 65:26]
      tag_2_3 <= 22'h0; // @[playground/src/noop/icache.scala 65:26]
    end else if (!(2'h0 == state)) begin // @[playground/src/noop/icache.scala 121:18]
      if (!(2'h1 == state)) begin // @[playground/src/noop/icache.scala 121:18]
        if (2'h2 == state) begin // @[playground/src/noop/icache.scala 121:18]
          tag_2_3 <= _GEN_532;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/icache.scala 65:26]
      tag_2_4 <= 22'h0; // @[playground/src/noop/icache.scala 65:26]
    end else if (!(2'h0 == state)) begin // @[playground/src/noop/icache.scala 121:18]
      if (!(2'h1 == state)) begin // @[playground/src/noop/icache.scala 121:18]
        if (2'h2 == state) begin // @[playground/src/noop/icache.scala 121:18]
          tag_2_4 <= _GEN_533;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/icache.scala 65:26]
      tag_2_5 <= 22'h0; // @[playground/src/noop/icache.scala 65:26]
    end else if (!(2'h0 == state)) begin // @[playground/src/noop/icache.scala 121:18]
      if (!(2'h1 == state)) begin // @[playground/src/noop/icache.scala 121:18]
        if (2'h2 == state) begin // @[playground/src/noop/icache.scala 121:18]
          tag_2_5 <= _GEN_534;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/icache.scala 65:26]
      tag_2_6 <= 22'h0; // @[playground/src/noop/icache.scala 65:26]
    end else if (!(2'h0 == state)) begin // @[playground/src/noop/icache.scala 121:18]
      if (!(2'h1 == state)) begin // @[playground/src/noop/icache.scala 121:18]
        if (2'h2 == state) begin // @[playground/src/noop/icache.scala 121:18]
          tag_2_6 <= _GEN_535;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/icache.scala 65:26]
      tag_2_7 <= 22'h0; // @[playground/src/noop/icache.scala 65:26]
    end else if (!(2'h0 == state)) begin // @[playground/src/noop/icache.scala 121:18]
      if (!(2'h1 == state)) begin // @[playground/src/noop/icache.scala 121:18]
        if (2'h2 == state) begin // @[playground/src/noop/icache.scala 121:18]
          tag_2_7 <= _GEN_536;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/icache.scala 65:26]
      tag_2_8 <= 22'h0; // @[playground/src/noop/icache.scala 65:26]
    end else if (!(2'h0 == state)) begin // @[playground/src/noop/icache.scala 121:18]
      if (!(2'h1 == state)) begin // @[playground/src/noop/icache.scala 121:18]
        if (2'h2 == state) begin // @[playground/src/noop/icache.scala 121:18]
          tag_2_8 <= _GEN_537;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/icache.scala 65:26]
      tag_2_9 <= 22'h0; // @[playground/src/noop/icache.scala 65:26]
    end else if (!(2'h0 == state)) begin // @[playground/src/noop/icache.scala 121:18]
      if (!(2'h1 == state)) begin // @[playground/src/noop/icache.scala 121:18]
        if (2'h2 == state) begin // @[playground/src/noop/icache.scala 121:18]
          tag_2_9 <= _GEN_538;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/icache.scala 65:26]
      tag_2_10 <= 22'h0; // @[playground/src/noop/icache.scala 65:26]
    end else if (!(2'h0 == state)) begin // @[playground/src/noop/icache.scala 121:18]
      if (!(2'h1 == state)) begin // @[playground/src/noop/icache.scala 121:18]
        if (2'h2 == state) begin // @[playground/src/noop/icache.scala 121:18]
          tag_2_10 <= _GEN_539;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/icache.scala 65:26]
      tag_2_11 <= 22'h0; // @[playground/src/noop/icache.scala 65:26]
    end else if (!(2'h0 == state)) begin // @[playground/src/noop/icache.scala 121:18]
      if (!(2'h1 == state)) begin // @[playground/src/noop/icache.scala 121:18]
        if (2'h2 == state) begin // @[playground/src/noop/icache.scala 121:18]
          tag_2_11 <= _GEN_540;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/icache.scala 65:26]
      tag_2_12 <= 22'h0; // @[playground/src/noop/icache.scala 65:26]
    end else if (!(2'h0 == state)) begin // @[playground/src/noop/icache.scala 121:18]
      if (!(2'h1 == state)) begin // @[playground/src/noop/icache.scala 121:18]
        if (2'h2 == state) begin // @[playground/src/noop/icache.scala 121:18]
          tag_2_12 <= _GEN_541;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/icache.scala 65:26]
      tag_2_13 <= 22'h0; // @[playground/src/noop/icache.scala 65:26]
    end else if (!(2'h0 == state)) begin // @[playground/src/noop/icache.scala 121:18]
      if (!(2'h1 == state)) begin // @[playground/src/noop/icache.scala 121:18]
        if (2'h2 == state) begin // @[playground/src/noop/icache.scala 121:18]
          tag_2_13 <= _GEN_542;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/icache.scala 65:26]
      tag_2_14 <= 22'h0; // @[playground/src/noop/icache.scala 65:26]
    end else if (!(2'h0 == state)) begin // @[playground/src/noop/icache.scala 121:18]
      if (!(2'h1 == state)) begin // @[playground/src/noop/icache.scala 121:18]
        if (2'h2 == state) begin // @[playground/src/noop/icache.scala 121:18]
          tag_2_14 <= _GEN_543;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/icache.scala 65:26]
      tag_2_15 <= 22'h0; // @[playground/src/noop/icache.scala 65:26]
    end else if (!(2'h0 == state)) begin // @[playground/src/noop/icache.scala 121:18]
      if (!(2'h1 == state)) begin // @[playground/src/noop/icache.scala 121:18]
        if (2'h2 == state) begin // @[playground/src/noop/icache.scala 121:18]
          tag_2_15 <= _GEN_544;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/icache.scala 65:26]
      tag_3_0 <= 22'h0; // @[playground/src/noop/icache.scala 65:26]
    end else if (!(2'h0 == state)) begin // @[playground/src/noop/icache.scala 121:18]
      if (!(2'h1 == state)) begin // @[playground/src/noop/icache.scala 121:18]
        if (2'h2 == state) begin // @[playground/src/noop/icache.scala 121:18]
          tag_3_0 <= _GEN_545;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/icache.scala 65:26]
      tag_3_1 <= 22'h0; // @[playground/src/noop/icache.scala 65:26]
    end else if (!(2'h0 == state)) begin // @[playground/src/noop/icache.scala 121:18]
      if (!(2'h1 == state)) begin // @[playground/src/noop/icache.scala 121:18]
        if (2'h2 == state) begin // @[playground/src/noop/icache.scala 121:18]
          tag_3_1 <= _GEN_546;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/icache.scala 65:26]
      tag_3_2 <= 22'h0; // @[playground/src/noop/icache.scala 65:26]
    end else if (!(2'h0 == state)) begin // @[playground/src/noop/icache.scala 121:18]
      if (!(2'h1 == state)) begin // @[playground/src/noop/icache.scala 121:18]
        if (2'h2 == state) begin // @[playground/src/noop/icache.scala 121:18]
          tag_3_2 <= _GEN_547;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/icache.scala 65:26]
      tag_3_3 <= 22'h0; // @[playground/src/noop/icache.scala 65:26]
    end else if (!(2'h0 == state)) begin // @[playground/src/noop/icache.scala 121:18]
      if (!(2'h1 == state)) begin // @[playground/src/noop/icache.scala 121:18]
        if (2'h2 == state) begin // @[playground/src/noop/icache.scala 121:18]
          tag_3_3 <= _GEN_548;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/icache.scala 65:26]
      tag_3_4 <= 22'h0; // @[playground/src/noop/icache.scala 65:26]
    end else if (!(2'h0 == state)) begin // @[playground/src/noop/icache.scala 121:18]
      if (!(2'h1 == state)) begin // @[playground/src/noop/icache.scala 121:18]
        if (2'h2 == state) begin // @[playground/src/noop/icache.scala 121:18]
          tag_3_4 <= _GEN_549;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/icache.scala 65:26]
      tag_3_5 <= 22'h0; // @[playground/src/noop/icache.scala 65:26]
    end else if (!(2'h0 == state)) begin // @[playground/src/noop/icache.scala 121:18]
      if (!(2'h1 == state)) begin // @[playground/src/noop/icache.scala 121:18]
        if (2'h2 == state) begin // @[playground/src/noop/icache.scala 121:18]
          tag_3_5 <= _GEN_550;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/icache.scala 65:26]
      tag_3_6 <= 22'h0; // @[playground/src/noop/icache.scala 65:26]
    end else if (!(2'h0 == state)) begin // @[playground/src/noop/icache.scala 121:18]
      if (!(2'h1 == state)) begin // @[playground/src/noop/icache.scala 121:18]
        if (2'h2 == state) begin // @[playground/src/noop/icache.scala 121:18]
          tag_3_6 <= _GEN_551;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/icache.scala 65:26]
      tag_3_7 <= 22'h0; // @[playground/src/noop/icache.scala 65:26]
    end else if (!(2'h0 == state)) begin // @[playground/src/noop/icache.scala 121:18]
      if (!(2'h1 == state)) begin // @[playground/src/noop/icache.scala 121:18]
        if (2'h2 == state) begin // @[playground/src/noop/icache.scala 121:18]
          tag_3_7 <= _GEN_552;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/icache.scala 65:26]
      tag_3_8 <= 22'h0; // @[playground/src/noop/icache.scala 65:26]
    end else if (!(2'h0 == state)) begin // @[playground/src/noop/icache.scala 121:18]
      if (!(2'h1 == state)) begin // @[playground/src/noop/icache.scala 121:18]
        if (2'h2 == state) begin // @[playground/src/noop/icache.scala 121:18]
          tag_3_8 <= _GEN_553;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/icache.scala 65:26]
      tag_3_9 <= 22'h0; // @[playground/src/noop/icache.scala 65:26]
    end else if (!(2'h0 == state)) begin // @[playground/src/noop/icache.scala 121:18]
      if (!(2'h1 == state)) begin // @[playground/src/noop/icache.scala 121:18]
        if (2'h2 == state) begin // @[playground/src/noop/icache.scala 121:18]
          tag_3_9 <= _GEN_554;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/icache.scala 65:26]
      tag_3_10 <= 22'h0; // @[playground/src/noop/icache.scala 65:26]
    end else if (!(2'h0 == state)) begin // @[playground/src/noop/icache.scala 121:18]
      if (!(2'h1 == state)) begin // @[playground/src/noop/icache.scala 121:18]
        if (2'h2 == state) begin // @[playground/src/noop/icache.scala 121:18]
          tag_3_10 <= _GEN_555;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/icache.scala 65:26]
      tag_3_11 <= 22'h0; // @[playground/src/noop/icache.scala 65:26]
    end else if (!(2'h0 == state)) begin // @[playground/src/noop/icache.scala 121:18]
      if (!(2'h1 == state)) begin // @[playground/src/noop/icache.scala 121:18]
        if (2'h2 == state) begin // @[playground/src/noop/icache.scala 121:18]
          tag_3_11 <= _GEN_556;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/icache.scala 65:26]
      tag_3_12 <= 22'h0; // @[playground/src/noop/icache.scala 65:26]
    end else if (!(2'h0 == state)) begin // @[playground/src/noop/icache.scala 121:18]
      if (!(2'h1 == state)) begin // @[playground/src/noop/icache.scala 121:18]
        if (2'h2 == state) begin // @[playground/src/noop/icache.scala 121:18]
          tag_3_12 <= _GEN_557;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/icache.scala 65:26]
      tag_3_13 <= 22'h0; // @[playground/src/noop/icache.scala 65:26]
    end else if (!(2'h0 == state)) begin // @[playground/src/noop/icache.scala 121:18]
      if (!(2'h1 == state)) begin // @[playground/src/noop/icache.scala 121:18]
        if (2'h2 == state) begin // @[playground/src/noop/icache.scala 121:18]
          tag_3_13 <= _GEN_558;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/icache.scala 65:26]
      tag_3_14 <= 22'h0; // @[playground/src/noop/icache.scala 65:26]
    end else if (!(2'h0 == state)) begin // @[playground/src/noop/icache.scala 121:18]
      if (!(2'h1 == state)) begin // @[playground/src/noop/icache.scala 121:18]
        if (2'h2 == state) begin // @[playground/src/noop/icache.scala 121:18]
          tag_3_14 <= _GEN_559;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/icache.scala 65:26]
      tag_3_15 <= 22'h0; // @[playground/src/noop/icache.scala 65:26]
    end else if (!(2'h0 == state)) begin // @[playground/src/noop/icache.scala 121:18]
      if (!(2'h1 == state)) begin // @[playground/src/noop/icache.scala 121:18]
        if (2'h2 == state) begin // @[playground/src/noop/icache.scala 121:18]
          tag_3_15 <= _GEN_560;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/icache.scala 66:26]
      valid_0_0 <= 1'h0; // @[playground/src/noop/icache.scala 66:26]
    end else if (2'h0 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_0_0 <= _GEN_130;
    end else if (2'h1 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_0_0 <= _GEN_130;
    end else if (2'h2 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_0_0 <= _GEN_561;
    end else begin
      valid_0_0 <= _GEN_130;
    end
    if (reset) begin // @[playground/src/noop/icache.scala 66:26]
      valid_0_1 <= 1'h0; // @[playground/src/noop/icache.scala 66:26]
    end else if (2'h0 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_0_1 <= _GEN_131;
    end else if (2'h1 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_0_1 <= _GEN_131;
    end else if (2'h2 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_0_1 <= _GEN_562;
    end else begin
      valid_0_1 <= _GEN_131;
    end
    if (reset) begin // @[playground/src/noop/icache.scala 66:26]
      valid_0_2 <= 1'h0; // @[playground/src/noop/icache.scala 66:26]
    end else if (2'h0 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_0_2 <= _GEN_132;
    end else if (2'h1 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_0_2 <= _GEN_132;
    end else if (2'h2 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_0_2 <= _GEN_563;
    end else begin
      valid_0_2 <= _GEN_132;
    end
    if (reset) begin // @[playground/src/noop/icache.scala 66:26]
      valid_0_3 <= 1'h0; // @[playground/src/noop/icache.scala 66:26]
    end else if (2'h0 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_0_3 <= _GEN_133;
    end else if (2'h1 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_0_3 <= _GEN_133;
    end else if (2'h2 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_0_3 <= _GEN_564;
    end else begin
      valid_0_3 <= _GEN_133;
    end
    if (reset) begin // @[playground/src/noop/icache.scala 66:26]
      valid_0_4 <= 1'h0; // @[playground/src/noop/icache.scala 66:26]
    end else if (2'h0 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_0_4 <= _GEN_134;
    end else if (2'h1 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_0_4 <= _GEN_134;
    end else if (2'h2 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_0_4 <= _GEN_565;
    end else begin
      valid_0_4 <= _GEN_134;
    end
    if (reset) begin // @[playground/src/noop/icache.scala 66:26]
      valid_0_5 <= 1'h0; // @[playground/src/noop/icache.scala 66:26]
    end else if (2'h0 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_0_5 <= _GEN_135;
    end else if (2'h1 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_0_5 <= _GEN_135;
    end else if (2'h2 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_0_5 <= _GEN_566;
    end else begin
      valid_0_5 <= _GEN_135;
    end
    if (reset) begin // @[playground/src/noop/icache.scala 66:26]
      valid_0_6 <= 1'h0; // @[playground/src/noop/icache.scala 66:26]
    end else if (2'h0 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_0_6 <= _GEN_136;
    end else if (2'h1 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_0_6 <= _GEN_136;
    end else if (2'h2 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_0_6 <= _GEN_567;
    end else begin
      valid_0_6 <= _GEN_136;
    end
    if (reset) begin // @[playground/src/noop/icache.scala 66:26]
      valid_0_7 <= 1'h0; // @[playground/src/noop/icache.scala 66:26]
    end else if (2'h0 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_0_7 <= _GEN_137;
    end else if (2'h1 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_0_7 <= _GEN_137;
    end else if (2'h2 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_0_7 <= _GEN_568;
    end else begin
      valid_0_7 <= _GEN_137;
    end
    if (reset) begin // @[playground/src/noop/icache.scala 66:26]
      valid_0_8 <= 1'h0; // @[playground/src/noop/icache.scala 66:26]
    end else if (2'h0 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_0_8 <= _GEN_138;
    end else if (2'h1 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_0_8 <= _GEN_138;
    end else if (2'h2 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_0_8 <= _GEN_569;
    end else begin
      valid_0_8 <= _GEN_138;
    end
    if (reset) begin // @[playground/src/noop/icache.scala 66:26]
      valid_0_9 <= 1'h0; // @[playground/src/noop/icache.scala 66:26]
    end else if (2'h0 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_0_9 <= _GEN_139;
    end else if (2'h1 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_0_9 <= _GEN_139;
    end else if (2'h2 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_0_9 <= _GEN_570;
    end else begin
      valid_0_9 <= _GEN_139;
    end
    if (reset) begin // @[playground/src/noop/icache.scala 66:26]
      valid_0_10 <= 1'h0; // @[playground/src/noop/icache.scala 66:26]
    end else if (2'h0 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_0_10 <= _GEN_140;
    end else if (2'h1 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_0_10 <= _GEN_140;
    end else if (2'h2 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_0_10 <= _GEN_571;
    end else begin
      valid_0_10 <= _GEN_140;
    end
    if (reset) begin // @[playground/src/noop/icache.scala 66:26]
      valid_0_11 <= 1'h0; // @[playground/src/noop/icache.scala 66:26]
    end else if (2'h0 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_0_11 <= _GEN_141;
    end else if (2'h1 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_0_11 <= _GEN_141;
    end else if (2'h2 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_0_11 <= _GEN_572;
    end else begin
      valid_0_11 <= _GEN_141;
    end
    if (reset) begin // @[playground/src/noop/icache.scala 66:26]
      valid_0_12 <= 1'h0; // @[playground/src/noop/icache.scala 66:26]
    end else if (2'h0 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_0_12 <= _GEN_142;
    end else if (2'h1 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_0_12 <= _GEN_142;
    end else if (2'h2 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_0_12 <= _GEN_573;
    end else begin
      valid_0_12 <= _GEN_142;
    end
    if (reset) begin // @[playground/src/noop/icache.scala 66:26]
      valid_0_13 <= 1'h0; // @[playground/src/noop/icache.scala 66:26]
    end else if (2'h0 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_0_13 <= _GEN_143;
    end else if (2'h1 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_0_13 <= _GEN_143;
    end else if (2'h2 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_0_13 <= _GEN_574;
    end else begin
      valid_0_13 <= _GEN_143;
    end
    if (reset) begin // @[playground/src/noop/icache.scala 66:26]
      valid_0_14 <= 1'h0; // @[playground/src/noop/icache.scala 66:26]
    end else if (2'h0 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_0_14 <= _GEN_144;
    end else if (2'h1 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_0_14 <= _GEN_144;
    end else if (2'h2 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_0_14 <= _GEN_575;
    end else begin
      valid_0_14 <= _GEN_144;
    end
    if (reset) begin // @[playground/src/noop/icache.scala 66:26]
      valid_0_15 <= 1'h0; // @[playground/src/noop/icache.scala 66:26]
    end else if (2'h0 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_0_15 <= _GEN_145;
    end else if (2'h1 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_0_15 <= _GEN_145;
    end else if (2'h2 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_0_15 <= _GEN_576;
    end else begin
      valid_0_15 <= _GEN_145;
    end
    if (reset) begin // @[playground/src/noop/icache.scala 66:26]
      valid_1_0 <= 1'h0; // @[playground/src/noop/icache.scala 66:26]
    end else if (2'h0 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_1_0 <= _GEN_146;
    end else if (2'h1 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_1_0 <= _GEN_146;
    end else if (2'h2 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_1_0 <= _GEN_577;
    end else begin
      valid_1_0 <= _GEN_146;
    end
    if (reset) begin // @[playground/src/noop/icache.scala 66:26]
      valid_1_1 <= 1'h0; // @[playground/src/noop/icache.scala 66:26]
    end else if (2'h0 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_1_1 <= _GEN_147;
    end else if (2'h1 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_1_1 <= _GEN_147;
    end else if (2'h2 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_1_1 <= _GEN_578;
    end else begin
      valid_1_1 <= _GEN_147;
    end
    if (reset) begin // @[playground/src/noop/icache.scala 66:26]
      valid_1_2 <= 1'h0; // @[playground/src/noop/icache.scala 66:26]
    end else if (2'h0 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_1_2 <= _GEN_148;
    end else if (2'h1 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_1_2 <= _GEN_148;
    end else if (2'h2 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_1_2 <= _GEN_579;
    end else begin
      valid_1_2 <= _GEN_148;
    end
    if (reset) begin // @[playground/src/noop/icache.scala 66:26]
      valid_1_3 <= 1'h0; // @[playground/src/noop/icache.scala 66:26]
    end else if (2'h0 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_1_3 <= _GEN_149;
    end else if (2'h1 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_1_3 <= _GEN_149;
    end else if (2'h2 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_1_3 <= _GEN_580;
    end else begin
      valid_1_3 <= _GEN_149;
    end
    if (reset) begin // @[playground/src/noop/icache.scala 66:26]
      valid_1_4 <= 1'h0; // @[playground/src/noop/icache.scala 66:26]
    end else if (2'h0 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_1_4 <= _GEN_150;
    end else if (2'h1 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_1_4 <= _GEN_150;
    end else if (2'h2 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_1_4 <= _GEN_581;
    end else begin
      valid_1_4 <= _GEN_150;
    end
    if (reset) begin // @[playground/src/noop/icache.scala 66:26]
      valid_1_5 <= 1'h0; // @[playground/src/noop/icache.scala 66:26]
    end else if (2'h0 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_1_5 <= _GEN_151;
    end else if (2'h1 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_1_5 <= _GEN_151;
    end else if (2'h2 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_1_5 <= _GEN_582;
    end else begin
      valid_1_5 <= _GEN_151;
    end
    if (reset) begin // @[playground/src/noop/icache.scala 66:26]
      valid_1_6 <= 1'h0; // @[playground/src/noop/icache.scala 66:26]
    end else if (2'h0 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_1_6 <= _GEN_152;
    end else if (2'h1 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_1_6 <= _GEN_152;
    end else if (2'h2 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_1_6 <= _GEN_583;
    end else begin
      valid_1_6 <= _GEN_152;
    end
    if (reset) begin // @[playground/src/noop/icache.scala 66:26]
      valid_1_7 <= 1'h0; // @[playground/src/noop/icache.scala 66:26]
    end else if (2'h0 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_1_7 <= _GEN_153;
    end else if (2'h1 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_1_7 <= _GEN_153;
    end else if (2'h2 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_1_7 <= _GEN_584;
    end else begin
      valid_1_7 <= _GEN_153;
    end
    if (reset) begin // @[playground/src/noop/icache.scala 66:26]
      valid_1_8 <= 1'h0; // @[playground/src/noop/icache.scala 66:26]
    end else if (2'h0 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_1_8 <= _GEN_154;
    end else if (2'h1 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_1_8 <= _GEN_154;
    end else if (2'h2 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_1_8 <= _GEN_585;
    end else begin
      valid_1_8 <= _GEN_154;
    end
    if (reset) begin // @[playground/src/noop/icache.scala 66:26]
      valid_1_9 <= 1'h0; // @[playground/src/noop/icache.scala 66:26]
    end else if (2'h0 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_1_9 <= _GEN_155;
    end else if (2'h1 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_1_9 <= _GEN_155;
    end else if (2'h2 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_1_9 <= _GEN_586;
    end else begin
      valid_1_9 <= _GEN_155;
    end
    if (reset) begin // @[playground/src/noop/icache.scala 66:26]
      valid_1_10 <= 1'h0; // @[playground/src/noop/icache.scala 66:26]
    end else if (2'h0 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_1_10 <= _GEN_156;
    end else if (2'h1 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_1_10 <= _GEN_156;
    end else if (2'h2 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_1_10 <= _GEN_587;
    end else begin
      valid_1_10 <= _GEN_156;
    end
    if (reset) begin // @[playground/src/noop/icache.scala 66:26]
      valid_1_11 <= 1'h0; // @[playground/src/noop/icache.scala 66:26]
    end else if (2'h0 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_1_11 <= _GEN_157;
    end else if (2'h1 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_1_11 <= _GEN_157;
    end else if (2'h2 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_1_11 <= _GEN_588;
    end else begin
      valid_1_11 <= _GEN_157;
    end
    if (reset) begin // @[playground/src/noop/icache.scala 66:26]
      valid_1_12 <= 1'h0; // @[playground/src/noop/icache.scala 66:26]
    end else if (2'h0 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_1_12 <= _GEN_158;
    end else if (2'h1 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_1_12 <= _GEN_158;
    end else if (2'h2 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_1_12 <= _GEN_589;
    end else begin
      valid_1_12 <= _GEN_158;
    end
    if (reset) begin // @[playground/src/noop/icache.scala 66:26]
      valid_1_13 <= 1'h0; // @[playground/src/noop/icache.scala 66:26]
    end else if (2'h0 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_1_13 <= _GEN_159;
    end else if (2'h1 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_1_13 <= _GEN_159;
    end else if (2'h2 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_1_13 <= _GEN_590;
    end else begin
      valid_1_13 <= _GEN_159;
    end
    if (reset) begin // @[playground/src/noop/icache.scala 66:26]
      valid_1_14 <= 1'h0; // @[playground/src/noop/icache.scala 66:26]
    end else if (2'h0 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_1_14 <= _GEN_160;
    end else if (2'h1 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_1_14 <= _GEN_160;
    end else if (2'h2 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_1_14 <= _GEN_591;
    end else begin
      valid_1_14 <= _GEN_160;
    end
    if (reset) begin // @[playground/src/noop/icache.scala 66:26]
      valid_1_15 <= 1'h0; // @[playground/src/noop/icache.scala 66:26]
    end else if (2'h0 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_1_15 <= _GEN_161;
    end else if (2'h1 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_1_15 <= _GEN_161;
    end else if (2'h2 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_1_15 <= _GEN_592;
    end else begin
      valid_1_15 <= _GEN_161;
    end
    if (reset) begin // @[playground/src/noop/icache.scala 66:26]
      valid_2_0 <= 1'h0; // @[playground/src/noop/icache.scala 66:26]
    end else if (2'h0 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_2_0 <= _GEN_162;
    end else if (2'h1 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_2_0 <= _GEN_162;
    end else if (2'h2 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_2_0 <= _GEN_593;
    end else begin
      valid_2_0 <= _GEN_162;
    end
    if (reset) begin // @[playground/src/noop/icache.scala 66:26]
      valid_2_1 <= 1'h0; // @[playground/src/noop/icache.scala 66:26]
    end else if (2'h0 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_2_1 <= _GEN_163;
    end else if (2'h1 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_2_1 <= _GEN_163;
    end else if (2'h2 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_2_1 <= _GEN_594;
    end else begin
      valid_2_1 <= _GEN_163;
    end
    if (reset) begin // @[playground/src/noop/icache.scala 66:26]
      valid_2_2 <= 1'h0; // @[playground/src/noop/icache.scala 66:26]
    end else if (2'h0 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_2_2 <= _GEN_164;
    end else if (2'h1 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_2_2 <= _GEN_164;
    end else if (2'h2 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_2_2 <= _GEN_595;
    end else begin
      valid_2_2 <= _GEN_164;
    end
    if (reset) begin // @[playground/src/noop/icache.scala 66:26]
      valid_2_3 <= 1'h0; // @[playground/src/noop/icache.scala 66:26]
    end else if (2'h0 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_2_3 <= _GEN_165;
    end else if (2'h1 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_2_3 <= _GEN_165;
    end else if (2'h2 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_2_3 <= _GEN_596;
    end else begin
      valid_2_3 <= _GEN_165;
    end
    if (reset) begin // @[playground/src/noop/icache.scala 66:26]
      valid_2_4 <= 1'h0; // @[playground/src/noop/icache.scala 66:26]
    end else if (2'h0 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_2_4 <= _GEN_166;
    end else if (2'h1 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_2_4 <= _GEN_166;
    end else if (2'h2 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_2_4 <= _GEN_597;
    end else begin
      valid_2_4 <= _GEN_166;
    end
    if (reset) begin // @[playground/src/noop/icache.scala 66:26]
      valid_2_5 <= 1'h0; // @[playground/src/noop/icache.scala 66:26]
    end else if (2'h0 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_2_5 <= _GEN_167;
    end else if (2'h1 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_2_5 <= _GEN_167;
    end else if (2'h2 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_2_5 <= _GEN_598;
    end else begin
      valid_2_5 <= _GEN_167;
    end
    if (reset) begin // @[playground/src/noop/icache.scala 66:26]
      valid_2_6 <= 1'h0; // @[playground/src/noop/icache.scala 66:26]
    end else if (2'h0 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_2_6 <= _GEN_168;
    end else if (2'h1 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_2_6 <= _GEN_168;
    end else if (2'h2 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_2_6 <= _GEN_599;
    end else begin
      valid_2_6 <= _GEN_168;
    end
    if (reset) begin // @[playground/src/noop/icache.scala 66:26]
      valid_2_7 <= 1'h0; // @[playground/src/noop/icache.scala 66:26]
    end else if (2'h0 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_2_7 <= _GEN_169;
    end else if (2'h1 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_2_7 <= _GEN_169;
    end else if (2'h2 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_2_7 <= _GEN_600;
    end else begin
      valid_2_7 <= _GEN_169;
    end
    if (reset) begin // @[playground/src/noop/icache.scala 66:26]
      valid_2_8 <= 1'h0; // @[playground/src/noop/icache.scala 66:26]
    end else if (2'h0 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_2_8 <= _GEN_170;
    end else if (2'h1 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_2_8 <= _GEN_170;
    end else if (2'h2 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_2_8 <= _GEN_601;
    end else begin
      valid_2_8 <= _GEN_170;
    end
    if (reset) begin // @[playground/src/noop/icache.scala 66:26]
      valid_2_9 <= 1'h0; // @[playground/src/noop/icache.scala 66:26]
    end else if (2'h0 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_2_9 <= _GEN_171;
    end else if (2'h1 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_2_9 <= _GEN_171;
    end else if (2'h2 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_2_9 <= _GEN_602;
    end else begin
      valid_2_9 <= _GEN_171;
    end
    if (reset) begin // @[playground/src/noop/icache.scala 66:26]
      valid_2_10 <= 1'h0; // @[playground/src/noop/icache.scala 66:26]
    end else if (2'h0 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_2_10 <= _GEN_172;
    end else if (2'h1 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_2_10 <= _GEN_172;
    end else if (2'h2 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_2_10 <= _GEN_603;
    end else begin
      valid_2_10 <= _GEN_172;
    end
    if (reset) begin // @[playground/src/noop/icache.scala 66:26]
      valid_2_11 <= 1'h0; // @[playground/src/noop/icache.scala 66:26]
    end else if (2'h0 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_2_11 <= _GEN_173;
    end else if (2'h1 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_2_11 <= _GEN_173;
    end else if (2'h2 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_2_11 <= _GEN_604;
    end else begin
      valid_2_11 <= _GEN_173;
    end
    if (reset) begin // @[playground/src/noop/icache.scala 66:26]
      valid_2_12 <= 1'h0; // @[playground/src/noop/icache.scala 66:26]
    end else if (2'h0 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_2_12 <= _GEN_174;
    end else if (2'h1 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_2_12 <= _GEN_174;
    end else if (2'h2 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_2_12 <= _GEN_605;
    end else begin
      valid_2_12 <= _GEN_174;
    end
    if (reset) begin // @[playground/src/noop/icache.scala 66:26]
      valid_2_13 <= 1'h0; // @[playground/src/noop/icache.scala 66:26]
    end else if (2'h0 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_2_13 <= _GEN_175;
    end else if (2'h1 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_2_13 <= _GEN_175;
    end else if (2'h2 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_2_13 <= _GEN_606;
    end else begin
      valid_2_13 <= _GEN_175;
    end
    if (reset) begin // @[playground/src/noop/icache.scala 66:26]
      valid_2_14 <= 1'h0; // @[playground/src/noop/icache.scala 66:26]
    end else if (2'h0 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_2_14 <= _GEN_176;
    end else if (2'h1 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_2_14 <= _GEN_176;
    end else if (2'h2 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_2_14 <= _GEN_607;
    end else begin
      valid_2_14 <= _GEN_176;
    end
    if (reset) begin // @[playground/src/noop/icache.scala 66:26]
      valid_2_15 <= 1'h0; // @[playground/src/noop/icache.scala 66:26]
    end else if (2'h0 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_2_15 <= _GEN_177;
    end else if (2'h1 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_2_15 <= _GEN_177;
    end else if (2'h2 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_2_15 <= _GEN_608;
    end else begin
      valid_2_15 <= _GEN_177;
    end
    if (reset) begin // @[playground/src/noop/icache.scala 66:26]
      valid_3_0 <= 1'h0; // @[playground/src/noop/icache.scala 66:26]
    end else if (2'h0 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_3_0 <= _GEN_178;
    end else if (2'h1 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_3_0 <= _GEN_178;
    end else if (2'h2 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_3_0 <= _GEN_609;
    end else begin
      valid_3_0 <= _GEN_178;
    end
    if (reset) begin // @[playground/src/noop/icache.scala 66:26]
      valid_3_1 <= 1'h0; // @[playground/src/noop/icache.scala 66:26]
    end else if (2'h0 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_3_1 <= _GEN_179;
    end else if (2'h1 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_3_1 <= _GEN_179;
    end else if (2'h2 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_3_1 <= _GEN_610;
    end else begin
      valid_3_1 <= _GEN_179;
    end
    if (reset) begin // @[playground/src/noop/icache.scala 66:26]
      valid_3_2 <= 1'h0; // @[playground/src/noop/icache.scala 66:26]
    end else if (2'h0 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_3_2 <= _GEN_180;
    end else if (2'h1 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_3_2 <= _GEN_180;
    end else if (2'h2 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_3_2 <= _GEN_611;
    end else begin
      valid_3_2 <= _GEN_180;
    end
    if (reset) begin // @[playground/src/noop/icache.scala 66:26]
      valid_3_3 <= 1'h0; // @[playground/src/noop/icache.scala 66:26]
    end else if (2'h0 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_3_3 <= _GEN_181;
    end else if (2'h1 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_3_3 <= _GEN_181;
    end else if (2'h2 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_3_3 <= _GEN_612;
    end else begin
      valid_3_3 <= _GEN_181;
    end
    if (reset) begin // @[playground/src/noop/icache.scala 66:26]
      valid_3_4 <= 1'h0; // @[playground/src/noop/icache.scala 66:26]
    end else if (2'h0 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_3_4 <= _GEN_182;
    end else if (2'h1 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_3_4 <= _GEN_182;
    end else if (2'h2 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_3_4 <= _GEN_613;
    end else begin
      valid_3_4 <= _GEN_182;
    end
    if (reset) begin // @[playground/src/noop/icache.scala 66:26]
      valid_3_5 <= 1'h0; // @[playground/src/noop/icache.scala 66:26]
    end else if (2'h0 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_3_5 <= _GEN_183;
    end else if (2'h1 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_3_5 <= _GEN_183;
    end else if (2'h2 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_3_5 <= _GEN_614;
    end else begin
      valid_3_5 <= _GEN_183;
    end
    if (reset) begin // @[playground/src/noop/icache.scala 66:26]
      valid_3_6 <= 1'h0; // @[playground/src/noop/icache.scala 66:26]
    end else if (2'h0 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_3_6 <= _GEN_184;
    end else if (2'h1 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_3_6 <= _GEN_184;
    end else if (2'h2 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_3_6 <= _GEN_615;
    end else begin
      valid_3_6 <= _GEN_184;
    end
    if (reset) begin // @[playground/src/noop/icache.scala 66:26]
      valid_3_7 <= 1'h0; // @[playground/src/noop/icache.scala 66:26]
    end else if (2'h0 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_3_7 <= _GEN_185;
    end else if (2'h1 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_3_7 <= _GEN_185;
    end else if (2'h2 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_3_7 <= _GEN_616;
    end else begin
      valid_3_7 <= _GEN_185;
    end
    if (reset) begin // @[playground/src/noop/icache.scala 66:26]
      valid_3_8 <= 1'h0; // @[playground/src/noop/icache.scala 66:26]
    end else if (2'h0 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_3_8 <= _GEN_186;
    end else if (2'h1 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_3_8 <= _GEN_186;
    end else if (2'h2 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_3_8 <= _GEN_617;
    end else begin
      valid_3_8 <= _GEN_186;
    end
    if (reset) begin // @[playground/src/noop/icache.scala 66:26]
      valid_3_9 <= 1'h0; // @[playground/src/noop/icache.scala 66:26]
    end else if (2'h0 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_3_9 <= _GEN_187;
    end else if (2'h1 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_3_9 <= _GEN_187;
    end else if (2'h2 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_3_9 <= _GEN_618;
    end else begin
      valid_3_9 <= _GEN_187;
    end
    if (reset) begin // @[playground/src/noop/icache.scala 66:26]
      valid_3_10 <= 1'h0; // @[playground/src/noop/icache.scala 66:26]
    end else if (2'h0 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_3_10 <= _GEN_188;
    end else if (2'h1 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_3_10 <= _GEN_188;
    end else if (2'h2 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_3_10 <= _GEN_619;
    end else begin
      valid_3_10 <= _GEN_188;
    end
    if (reset) begin // @[playground/src/noop/icache.scala 66:26]
      valid_3_11 <= 1'h0; // @[playground/src/noop/icache.scala 66:26]
    end else if (2'h0 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_3_11 <= _GEN_189;
    end else if (2'h1 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_3_11 <= _GEN_189;
    end else if (2'h2 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_3_11 <= _GEN_620;
    end else begin
      valid_3_11 <= _GEN_189;
    end
    if (reset) begin // @[playground/src/noop/icache.scala 66:26]
      valid_3_12 <= 1'h0; // @[playground/src/noop/icache.scala 66:26]
    end else if (2'h0 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_3_12 <= _GEN_190;
    end else if (2'h1 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_3_12 <= _GEN_190;
    end else if (2'h2 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_3_12 <= _GEN_621;
    end else begin
      valid_3_12 <= _GEN_190;
    end
    if (reset) begin // @[playground/src/noop/icache.scala 66:26]
      valid_3_13 <= 1'h0; // @[playground/src/noop/icache.scala 66:26]
    end else if (2'h0 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_3_13 <= _GEN_191;
    end else if (2'h1 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_3_13 <= _GEN_191;
    end else if (2'h2 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_3_13 <= _GEN_622;
    end else begin
      valid_3_13 <= _GEN_191;
    end
    if (reset) begin // @[playground/src/noop/icache.scala 66:26]
      valid_3_14 <= 1'h0; // @[playground/src/noop/icache.scala 66:26]
    end else if (2'h0 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_3_14 <= _GEN_192;
    end else if (2'h1 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_3_14 <= _GEN_192;
    end else if (2'h2 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_3_14 <= _GEN_623;
    end else begin
      valid_3_14 <= _GEN_192;
    end
    if (reset) begin // @[playground/src/noop/icache.scala 66:26]
      valid_3_15 <= 1'h0; // @[playground/src/noop/icache.scala 66:26]
    end else if (2'h0 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_3_15 <= _GEN_193;
    end else if (2'h1 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_3_15 <= _GEN_193;
    end else if (2'h2 == state) begin // @[playground/src/noop/icache.scala 121:18]
      valid_3_15 <= _GEN_624;
    end else begin
      valid_3_15 <= _GEN_193;
    end
    if (reset) begin // @[playground/src/noop/icache.scala 71:30]
      wait_r <= 1'h0; // @[playground/src/noop/icache.scala 71:30]
    end else if (2'h0 == state) begin // @[playground/src/noop/icache.scala 121:18]
      if (!(~hs_in & _io_icRead_ready_T)) begin // @[playground/src/noop/icache.scala 123:36]
        if (cacheHit) begin // @[playground/src/noop/icache.scala 125:33]
          wait_r <= 1'h0; // @[playground/src/noop/icache.scala 127:25]
        end else begin
          wait_r <= 1'h1; // @[playground/src/noop/icache.scala 133:25]
        end
      end
    end
    if (reset) begin // @[playground/src/noop/icache.scala 72:30]
      valid_r <= 1'h0; // @[playground/src/noop/icache.scala 72:30]
    end else begin
      valid_r <= _GEN_893;
    end
    if (reset) begin // @[playground/src/noop/icache.scala 78:34]
      addr_r <= 32'h0; // @[playground/src/noop/icache.scala 78:34]
    end else if (hs_in) begin // @[playground/src/noop/icache.scala 82:30]
      addr_r <= io_icRead_addr;
    end
    if (reset) begin // @[playground/src/noop/icache.scala 79:34]
      matchWay_r <= 32'h0; // @[playground/src/noop/icache.scala 79:34]
    end else if (hs_in) begin // @[playground/src/noop/icache.scala 90:30]
      matchWay_r <= {{30'd0}, matchWay};
    end
    if (reset) begin // @[playground/src/noop/icache.scala 80:34]
      axiOffset <= 3'h0; // @[playground/src/noop/icache.scala 80:34]
    end else if (!(2'h0 == state)) begin // @[playground/src/noop/icache.scala 121:18]
      if (2'h1 == state) begin // @[playground/src/noop/icache.scala 121:18]
        if (raddrEn & io_instAxi_ra_ready) begin // @[playground/src/noop/icache.scala 137:49]
          axiOffset <= 3'h0; // @[playground/src/noop/icache.scala 141:27]
        end
      end else if (2'h2 == state) begin // @[playground/src/noop/icache.scala 121:18]
        axiOffset <= _GEN_493;
      end
    end
    if (reset) begin // @[playground/src/noop/icache.scala 81:34]
      databuf <= 64'h0; // @[playground/src/noop/icache.scala 81:34]
    end else if (!(2'h0 == state)) begin // @[playground/src/noop/icache.scala 121:18]
      if (!(2'h1 == state)) begin // @[playground/src/noop/icache.scala 121:18]
        if (2'h2 == state) begin // @[playground/src/noop/icache.scala 121:18]
          databuf <= _GEN_495;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/icache.scala 102:24]
      state <= 2'h0; // @[playground/src/noop/icache.scala 102:24]
    end else if (2'h0 == state) begin // @[playground/src/noop/icache.scala 121:18]
      if (!(~hs_in & _io_icRead_ready_T)) begin // @[playground/src/noop/icache.scala 123:36]
        if (!(cacheHit)) begin // @[playground/src/noop/icache.scala 125:33]
          state <= 2'h1; // @[playground/src/noop/icache.scala 131:25]
        end
      end
    end else if (2'h1 == state) begin // @[playground/src/noop/icache.scala 121:18]
      if (raddrEn & io_instAxi_ra_ready) begin // @[playground/src/noop/icache.scala 137:49]
        state <= 2'h2; // @[playground/src/noop/icache.scala 138:25]
      end
    end else if (2'h2 == state) begin // @[playground/src/noop/icache.scala 121:18]
      state <= _GEN_625;
    end
    if (reset) begin // @[playground/src/noop/icache.scala 119:30]
      rdataEn <= 1'h0; // @[playground/src/noop/icache.scala 119:30]
    end else if (!(2'h0 == state)) begin // @[playground/src/noop/icache.scala 121:18]
      if (2'h1 == state) begin // @[playground/src/noop/icache.scala 121:18]
        rdataEn <= _GEN_230;
      end else if (2'h2 == state) begin // @[playground/src/noop/icache.scala 121:18]
        rdataEn <= _GEN_496;
      end
    end
    if (reset) begin // @[playground/src/noop/icache.scala 117:30]
      raddrEn <= 1'h0; // @[playground/src/noop/icache.scala 117:30]
    end else if (2'h0 == state) begin // @[playground/src/noop/icache.scala 121:18]
      if (!(~hs_in & _io_icRead_ready_T)) begin // @[playground/src/noop/icache.scala 123:36]
        if (!(cacheHit)) begin // @[playground/src/noop/icache.scala 125:33]
          raddrEn <= 1'h1; // @[playground/src/noop/icache.scala 130:25]
        end
      end
    end else if (2'h1 == state) begin // @[playground/src/noop/icache.scala 121:18]
      if (raddrEn & io_instAxi_ra_ready) begin // @[playground/src/noop/icache.scala 137:49]
        raddrEn <= 1'h0; // @[playground/src/noop/icache.scala 139:25]
      end
    end
    if (reset) begin // @[playground/src/noop/icache.scala 118:30]
      raddr <= 32'h0; // @[playground/src/noop/icache.scala 118:30]
    end else if (2'h0 == state) begin // @[playground/src/noop/icache.scala 121:18]
      if (!(~hs_in & _io_icRead_ready_T)) begin // @[playground/src/noop/icache.scala 123:36]
        if (!(cacheHit)) begin // @[playground/src/noop/icache.scala 125:33]
          raddr <= _raddr_T; // @[playground/src/noop/icache.scala 129:25]
        end
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  tag_0_0 = _RAND_0[21:0];
  _RAND_1 = {1{`RANDOM}};
  tag_0_1 = _RAND_1[21:0];
  _RAND_2 = {1{`RANDOM}};
  tag_0_2 = _RAND_2[21:0];
  _RAND_3 = {1{`RANDOM}};
  tag_0_3 = _RAND_3[21:0];
  _RAND_4 = {1{`RANDOM}};
  tag_0_4 = _RAND_4[21:0];
  _RAND_5 = {1{`RANDOM}};
  tag_0_5 = _RAND_5[21:0];
  _RAND_6 = {1{`RANDOM}};
  tag_0_6 = _RAND_6[21:0];
  _RAND_7 = {1{`RANDOM}};
  tag_0_7 = _RAND_7[21:0];
  _RAND_8 = {1{`RANDOM}};
  tag_0_8 = _RAND_8[21:0];
  _RAND_9 = {1{`RANDOM}};
  tag_0_9 = _RAND_9[21:0];
  _RAND_10 = {1{`RANDOM}};
  tag_0_10 = _RAND_10[21:0];
  _RAND_11 = {1{`RANDOM}};
  tag_0_11 = _RAND_11[21:0];
  _RAND_12 = {1{`RANDOM}};
  tag_0_12 = _RAND_12[21:0];
  _RAND_13 = {1{`RANDOM}};
  tag_0_13 = _RAND_13[21:0];
  _RAND_14 = {1{`RANDOM}};
  tag_0_14 = _RAND_14[21:0];
  _RAND_15 = {1{`RANDOM}};
  tag_0_15 = _RAND_15[21:0];
  _RAND_16 = {1{`RANDOM}};
  tag_1_0 = _RAND_16[21:0];
  _RAND_17 = {1{`RANDOM}};
  tag_1_1 = _RAND_17[21:0];
  _RAND_18 = {1{`RANDOM}};
  tag_1_2 = _RAND_18[21:0];
  _RAND_19 = {1{`RANDOM}};
  tag_1_3 = _RAND_19[21:0];
  _RAND_20 = {1{`RANDOM}};
  tag_1_4 = _RAND_20[21:0];
  _RAND_21 = {1{`RANDOM}};
  tag_1_5 = _RAND_21[21:0];
  _RAND_22 = {1{`RANDOM}};
  tag_1_6 = _RAND_22[21:0];
  _RAND_23 = {1{`RANDOM}};
  tag_1_7 = _RAND_23[21:0];
  _RAND_24 = {1{`RANDOM}};
  tag_1_8 = _RAND_24[21:0];
  _RAND_25 = {1{`RANDOM}};
  tag_1_9 = _RAND_25[21:0];
  _RAND_26 = {1{`RANDOM}};
  tag_1_10 = _RAND_26[21:0];
  _RAND_27 = {1{`RANDOM}};
  tag_1_11 = _RAND_27[21:0];
  _RAND_28 = {1{`RANDOM}};
  tag_1_12 = _RAND_28[21:0];
  _RAND_29 = {1{`RANDOM}};
  tag_1_13 = _RAND_29[21:0];
  _RAND_30 = {1{`RANDOM}};
  tag_1_14 = _RAND_30[21:0];
  _RAND_31 = {1{`RANDOM}};
  tag_1_15 = _RAND_31[21:0];
  _RAND_32 = {1{`RANDOM}};
  tag_2_0 = _RAND_32[21:0];
  _RAND_33 = {1{`RANDOM}};
  tag_2_1 = _RAND_33[21:0];
  _RAND_34 = {1{`RANDOM}};
  tag_2_2 = _RAND_34[21:0];
  _RAND_35 = {1{`RANDOM}};
  tag_2_3 = _RAND_35[21:0];
  _RAND_36 = {1{`RANDOM}};
  tag_2_4 = _RAND_36[21:0];
  _RAND_37 = {1{`RANDOM}};
  tag_2_5 = _RAND_37[21:0];
  _RAND_38 = {1{`RANDOM}};
  tag_2_6 = _RAND_38[21:0];
  _RAND_39 = {1{`RANDOM}};
  tag_2_7 = _RAND_39[21:0];
  _RAND_40 = {1{`RANDOM}};
  tag_2_8 = _RAND_40[21:0];
  _RAND_41 = {1{`RANDOM}};
  tag_2_9 = _RAND_41[21:0];
  _RAND_42 = {1{`RANDOM}};
  tag_2_10 = _RAND_42[21:0];
  _RAND_43 = {1{`RANDOM}};
  tag_2_11 = _RAND_43[21:0];
  _RAND_44 = {1{`RANDOM}};
  tag_2_12 = _RAND_44[21:0];
  _RAND_45 = {1{`RANDOM}};
  tag_2_13 = _RAND_45[21:0];
  _RAND_46 = {1{`RANDOM}};
  tag_2_14 = _RAND_46[21:0];
  _RAND_47 = {1{`RANDOM}};
  tag_2_15 = _RAND_47[21:0];
  _RAND_48 = {1{`RANDOM}};
  tag_3_0 = _RAND_48[21:0];
  _RAND_49 = {1{`RANDOM}};
  tag_3_1 = _RAND_49[21:0];
  _RAND_50 = {1{`RANDOM}};
  tag_3_2 = _RAND_50[21:0];
  _RAND_51 = {1{`RANDOM}};
  tag_3_3 = _RAND_51[21:0];
  _RAND_52 = {1{`RANDOM}};
  tag_3_4 = _RAND_52[21:0];
  _RAND_53 = {1{`RANDOM}};
  tag_3_5 = _RAND_53[21:0];
  _RAND_54 = {1{`RANDOM}};
  tag_3_6 = _RAND_54[21:0];
  _RAND_55 = {1{`RANDOM}};
  tag_3_7 = _RAND_55[21:0];
  _RAND_56 = {1{`RANDOM}};
  tag_3_8 = _RAND_56[21:0];
  _RAND_57 = {1{`RANDOM}};
  tag_3_9 = _RAND_57[21:0];
  _RAND_58 = {1{`RANDOM}};
  tag_3_10 = _RAND_58[21:0];
  _RAND_59 = {1{`RANDOM}};
  tag_3_11 = _RAND_59[21:0];
  _RAND_60 = {1{`RANDOM}};
  tag_3_12 = _RAND_60[21:0];
  _RAND_61 = {1{`RANDOM}};
  tag_3_13 = _RAND_61[21:0];
  _RAND_62 = {1{`RANDOM}};
  tag_3_14 = _RAND_62[21:0];
  _RAND_63 = {1{`RANDOM}};
  tag_3_15 = _RAND_63[21:0];
  _RAND_64 = {1{`RANDOM}};
  valid_0_0 = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  valid_0_1 = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  valid_0_2 = _RAND_66[0:0];
  _RAND_67 = {1{`RANDOM}};
  valid_0_3 = _RAND_67[0:0];
  _RAND_68 = {1{`RANDOM}};
  valid_0_4 = _RAND_68[0:0];
  _RAND_69 = {1{`RANDOM}};
  valid_0_5 = _RAND_69[0:0];
  _RAND_70 = {1{`RANDOM}};
  valid_0_6 = _RAND_70[0:0];
  _RAND_71 = {1{`RANDOM}};
  valid_0_7 = _RAND_71[0:0];
  _RAND_72 = {1{`RANDOM}};
  valid_0_8 = _RAND_72[0:0];
  _RAND_73 = {1{`RANDOM}};
  valid_0_9 = _RAND_73[0:0];
  _RAND_74 = {1{`RANDOM}};
  valid_0_10 = _RAND_74[0:0];
  _RAND_75 = {1{`RANDOM}};
  valid_0_11 = _RAND_75[0:0];
  _RAND_76 = {1{`RANDOM}};
  valid_0_12 = _RAND_76[0:0];
  _RAND_77 = {1{`RANDOM}};
  valid_0_13 = _RAND_77[0:0];
  _RAND_78 = {1{`RANDOM}};
  valid_0_14 = _RAND_78[0:0];
  _RAND_79 = {1{`RANDOM}};
  valid_0_15 = _RAND_79[0:0];
  _RAND_80 = {1{`RANDOM}};
  valid_1_0 = _RAND_80[0:0];
  _RAND_81 = {1{`RANDOM}};
  valid_1_1 = _RAND_81[0:0];
  _RAND_82 = {1{`RANDOM}};
  valid_1_2 = _RAND_82[0:0];
  _RAND_83 = {1{`RANDOM}};
  valid_1_3 = _RAND_83[0:0];
  _RAND_84 = {1{`RANDOM}};
  valid_1_4 = _RAND_84[0:0];
  _RAND_85 = {1{`RANDOM}};
  valid_1_5 = _RAND_85[0:0];
  _RAND_86 = {1{`RANDOM}};
  valid_1_6 = _RAND_86[0:0];
  _RAND_87 = {1{`RANDOM}};
  valid_1_7 = _RAND_87[0:0];
  _RAND_88 = {1{`RANDOM}};
  valid_1_8 = _RAND_88[0:0];
  _RAND_89 = {1{`RANDOM}};
  valid_1_9 = _RAND_89[0:0];
  _RAND_90 = {1{`RANDOM}};
  valid_1_10 = _RAND_90[0:0];
  _RAND_91 = {1{`RANDOM}};
  valid_1_11 = _RAND_91[0:0];
  _RAND_92 = {1{`RANDOM}};
  valid_1_12 = _RAND_92[0:0];
  _RAND_93 = {1{`RANDOM}};
  valid_1_13 = _RAND_93[0:0];
  _RAND_94 = {1{`RANDOM}};
  valid_1_14 = _RAND_94[0:0];
  _RAND_95 = {1{`RANDOM}};
  valid_1_15 = _RAND_95[0:0];
  _RAND_96 = {1{`RANDOM}};
  valid_2_0 = _RAND_96[0:0];
  _RAND_97 = {1{`RANDOM}};
  valid_2_1 = _RAND_97[0:0];
  _RAND_98 = {1{`RANDOM}};
  valid_2_2 = _RAND_98[0:0];
  _RAND_99 = {1{`RANDOM}};
  valid_2_3 = _RAND_99[0:0];
  _RAND_100 = {1{`RANDOM}};
  valid_2_4 = _RAND_100[0:0];
  _RAND_101 = {1{`RANDOM}};
  valid_2_5 = _RAND_101[0:0];
  _RAND_102 = {1{`RANDOM}};
  valid_2_6 = _RAND_102[0:0];
  _RAND_103 = {1{`RANDOM}};
  valid_2_7 = _RAND_103[0:0];
  _RAND_104 = {1{`RANDOM}};
  valid_2_8 = _RAND_104[0:0];
  _RAND_105 = {1{`RANDOM}};
  valid_2_9 = _RAND_105[0:0];
  _RAND_106 = {1{`RANDOM}};
  valid_2_10 = _RAND_106[0:0];
  _RAND_107 = {1{`RANDOM}};
  valid_2_11 = _RAND_107[0:0];
  _RAND_108 = {1{`RANDOM}};
  valid_2_12 = _RAND_108[0:0];
  _RAND_109 = {1{`RANDOM}};
  valid_2_13 = _RAND_109[0:0];
  _RAND_110 = {1{`RANDOM}};
  valid_2_14 = _RAND_110[0:0];
  _RAND_111 = {1{`RANDOM}};
  valid_2_15 = _RAND_111[0:0];
  _RAND_112 = {1{`RANDOM}};
  valid_3_0 = _RAND_112[0:0];
  _RAND_113 = {1{`RANDOM}};
  valid_3_1 = _RAND_113[0:0];
  _RAND_114 = {1{`RANDOM}};
  valid_3_2 = _RAND_114[0:0];
  _RAND_115 = {1{`RANDOM}};
  valid_3_3 = _RAND_115[0:0];
  _RAND_116 = {1{`RANDOM}};
  valid_3_4 = _RAND_116[0:0];
  _RAND_117 = {1{`RANDOM}};
  valid_3_5 = _RAND_117[0:0];
  _RAND_118 = {1{`RANDOM}};
  valid_3_6 = _RAND_118[0:0];
  _RAND_119 = {1{`RANDOM}};
  valid_3_7 = _RAND_119[0:0];
  _RAND_120 = {1{`RANDOM}};
  valid_3_8 = _RAND_120[0:0];
  _RAND_121 = {1{`RANDOM}};
  valid_3_9 = _RAND_121[0:0];
  _RAND_122 = {1{`RANDOM}};
  valid_3_10 = _RAND_122[0:0];
  _RAND_123 = {1{`RANDOM}};
  valid_3_11 = _RAND_123[0:0];
  _RAND_124 = {1{`RANDOM}};
  valid_3_12 = _RAND_124[0:0];
  _RAND_125 = {1{`RANDOM}};
  valid_3_13 = _RAND_125[0:0];
  _RAND_126 = {1{`RANDOM}};
  valid_3_14 = _RAND_126[0:0];
  _RAND_127 = {1{`RANDOM}};
  valid_3_15 = _RAND_127[0:0];
  _RAND_128 = {1{`RANDOM}};
  wait_r = _RAND_128[0:0];
  _RAND_129 = {1{`RANDOM}};
  valid_r = _RAND_129[0:0];
  _RAND_130 = {1{`RANDOM}};
  addr_r = _RAND_130[31:0];
  _RAND_131 = {1{`RANDOM}};
  matchWay_r = _RAND_131[31:0];
  _RAND_132 = {1{`RANDOM}};
  axiOffset = _RAND_132[2:0];
  _RAND_133 = {2{`RANDOM}};
  databuf = _RAND_133[63:0];
  _RAND_134 = {1{`RANDOM}};
  state = _RAND_134[1:0];
  _RAND_135 = {1{`RANDOM}};
  rdataEn = _RAND_135[0:0];
  _RAND_136 = {1{`RANDOM}};
  raddrEn = _RAND_136[0:0];
  _RAND_137 = {1{`RANDOM}};
  raddr = _RAND_137[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module DataCache(
  input         clock,
  input         reset,
  input         io_dataAxi_wa_ready, // @[playground/src/noop/dcache.scala 81:16]
  output        io_dataAxi_wa_valid, // @[playground/src/noop/dcache.scala 81:16]
  output [31:0] io_dataAxi_wa_bits_addr, // @[playground/src/noop/dcache.scala 81:16]
  input         io_dataAxi_wd_ready, // @[playground/src/noop/dcache.scala 81:16]
  output        io_dataAxi_wd_valid, // @[playground/src/noop/dcache.scala 81:16]
  output [63:0] io_dataAxi_wd_bits_data, // @[playground/src/noop/dcache.scala 81:16]
  output        io_dataAxi_wd_bits_last, // @[playground/src/noop/dcache.scala 81:16]
  input         io_dataAxi_ra_ready, // @[playground/src/noop/dcache.scala 81:16]
  output        io_dataAxi_ra_valid, // @[playground/src/noop/dcache.scala 81:16]
  output [31:0] io_dataAxi_ra_bits_addr, // @[playground/src/noop/dcache.scala 81:16]
  input         io_dataAxi_rd_valid, // @[playground/src/noop/dcache.scala 81:16]
  input  [63:0] io_dataAxi_rd_bits_data, // @[playground/src/noop/dcache.scala 81:16]
  input         io_dataAxi_rd_bits_last, // @[playground/src/noop/dcache.scala 81:16]
  input  [31:0] io_dcRW_addr, // @[playground/src/noop/dcache.scala 81:16]
  output [63:0] io_dcRW_rdata, // @[playground/src/noop/dcache.scala 81:16]
  output        io_dcRW_rvalid, // @[playground/src/noop/dcache.scala 81:16]
  input  [63:0] io_dcRW_wdata, // @[playground/src/noop/dcache.scala 81:16]
  input  [4:0]  io_dcRW_dc_mode, // @[playground/src/noop/dcache.scala 81:16]
  input  [4:0]  io_dcRW_amo, // @[playground/src/noop/dcache.scala 81:16]
  output        io_dcRW_ready, // @[playground/src/noop/dcache.scala 81:16]
  input         io_flush, // @[playground/src/noop/dcache.scala 81:16]
  output        io_flush_out // @[playground/src/noop/dcache.scala 81:16]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [63:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [63:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
`endif // RANDOMIZE_REG_INIT
  wire  Ram_bw_clock; // @[playground/src/noop/dcache.scala 91:57]
  wire  Ram_bw_reset; // @[playground/src/noop/dcache.scala 91:57]
  wire  Ram_bw_io_cen; // @[playground/src/noop/dcache.scala 91:57]
  wire  Ram_bw_io_wen; // @[playground/src/noop/dcache.scala 91:57]
  wire [5:0] Ram_bw_io_addr; // @[playground/src/noop/dcache.scala 91:57]
  wire [127:0] Ram_bw_io_rdata; // @[playground/src/noop/dcache.scala 91:57]
  wire [127:0] Ram_bw_io_wdata; // @[playground/src/noop/dcache.scala 91:57]
  wire [127:0] Ram_bw_io_mask; // @[playground/src/noop/dcache.scala 91:57]
  wire  Ram_bw_1_clock; // @[playground/src/noop/dcache.scala 91:57]
  wire  Ram_bw_1_reset; // @[playground/src/noop/dcache.scala 91:57]
  wire  Ram_bw_1_io_cen; // @[playground/src/noop/dcache.scala 91:57]
  wire  Ram_bw_1_io_wen; // @[playground/src/noop/dcache.scala 91:57]
  wire [5:0] Ram_bw_1_io_addr; // @[playground/src/noop/dcache.scala 91:57]
  wire [127:0] Ram_bw_1_io_rdata; // @[playground/src/noop/dcache.scala 91:57]
  wire [127:0] Ram_bw_1_io_wdata; // @[playground/src/noop/dcache.scala 91:57]
  wire [127:0] Ram_bw_1_io_mask; // @[playground/src/noop/dcache.scala 91:57]
  wire  Ram_bw_2_clock; // @[playground/src/noop/dcache.scala 91:57]
  wire  Ram_bw_2_reset; // @[playground/src/noop/dcache.scala 91:57]
  wire  Ram_bw_2_io_cen; // @[playground/src/noop/dcache.scala 91:57]
  wire  Ram_bw_2_io_wen; // @[playground/src/noop/dcache.scala 91:57]
  wire [5:0] Ram_bw_2_io_addr; // @[playground/src/noop/dcache.scala 91:57]
  wire [127:0] Ram_bw_2_io_rdata; // @[playground/src/noop/dcache.scala 91:57]
  wire [127:0] Ram_bw_2_io_wdata; // @[playground/src/noop/dcache.scala 91:57]
  wire [127:0] Ram_bw_2_io_mask; // @[playground/src/noop/dcache.scala 91:57]
  wire  Ram_bw_3_clock; // @[playground/src/noop/dcache.scala 91:57]
  wire  Ram_bw_3_reset; // @[playground/src/noop/dcache.scala 91:57]
  wire  Ram_bw_3_io_cen; // @[playground/src/noop/dcache.scala 91:57]
  wire  Ram_bw_3_io_wen; // @[playground/src/noop/dcache.scala 91:57]
  wire [5:0] Ram_bw_3_io_addr; // @[playground/src/noop/dcache.scala 91:57]
  wire [127:0] Ram_bw_3_io_rdata; // @[playground/src/noop/dcache.scala 91:57]
  wire [127:0] Ram_bw_3_io_wdata; // @[playground/src/noop/dcache.scala 91:57]
  wire [127:0] Ram_bw_3_io_mask; // @[playground/src/noop/dcache.scala 91:57]
  wire  matchWay_prng_clock; // @[src/main/scala/chisel3/util/random/PRNG.scala 91:22]
  wire  matchWay_prng_reset; // @[src/main/scala/chisel3/util/random/PRNG.scala 91:22]
  wire  matchWay_prng_io_out_0; // @[src/main/scala/chisel3/util/random/PRNG.scala 91:22]
  wire  matchWay_prng_io_out_1; // @[src/main/scala/chisel3/util/random/PRNG.scala 91:22]
  reg [21:0] tag_0_0; // @[playground/src/noop/dcache.scala 88:26]
  reg [21:0] tag_0_1; // @[playground/src/noop/dcache.scala 88:26]
  reg [21:0] tag_0_2; // @[playground/src/noop/dcache.scala 88:26]
  reg [21:0] tag_0_3; // @[playground/src/noop/dcache.scala 88:26]
  reg [21:0] tag_0_4; // @[playground/src/noop/dcache.scala 88:26]
  reg [21:0] tag_0_5; // @[playground/src/noop/dcache.scala 88:26]
  reg [21:0] tag_0_6; // @[playground/src/noop/dcache.scala 88:26]
  reg [21:0] tag_0_7; // @[playground/src/noop/dcache.scala 88:26]
  reg [21:0] tag_0_8; // @[playground/src/noop/dcache.scala 88:26]
  reg [21:0] tag_0_9; // @[playground/src/noop/dcache.scala 88:26]
  reg [21:0] tag_0_10; // @[playground/src/noop/dcache.scala 88:26]
  reg [21:0] tag_0_11; // @[playground/src/noop/dcache.scala 88:26]
  reg [21:0] tag_0_12; // @[playground/src/noop/dcache.scala 88:26]
  reg [21:0] tag_0_13; // @[playground/src/noop/dcache.scala 88:26]
  reg [21:0] tag_0_14; // @[playground/src/noop/dcache.scala 88:26]
  reg [21:0] tag_0_15; // @[playground/src/noop/dcache.scala 88:26]
  reg [21:0] tag_1_0; // @[playground/src/noop/dcache.scala 88:26]
  reg [21:0] tag_1_1; // @[playground/src/noop/dcache.scala 88:26]
  reg [21:0] tag_1_2; // @[playground/src/noop/dcache.scala 88:26]
  reg [21:0] tag_1_3; // @[playground/src/noop/dcache.scala 88:26]
  reg [21:0] tag_1_4; // @[playground/src/noop/dcache.scala 88:26]
  reg [21:0] tag_1_5; // @[playground/src/noop/dcache.scala 88:26]
  reg [21:0] tag_1_6; // @[playground/src/noop/dcache.scala 88:26]
  reg [21:0] tag_1_7; // @[playground/src/noop/dcache.scala 88:26]
  reg [21:0] tag_1_8; // @[playground/src/noop/dcache.scala 88:26]
  reg [21:0] tag_1_9; // @[playground/src/noop/dcache.scala 88:26]
  reg [21:0] tag_1_10; // @[playground/src/noop/dcache.scala 88:26]
  reg [21:0] tag_1_11; // @[playground/src/noop/dcache.scala 88:26]
  reg [21:0] tag_1_12; // @[playground/src/noop/dcache.scala 88:26]
  reg [21:0] tag_1_13; // @[playground/src/noop/dcache.scala 88:26]
  reg [21:0] tag_1_14; // @[playground/src/noop/dcache.scala 88:26]
  reg [21:0] tag_1_15; // @[playground/src/noop/dcache.scala 88:26]
  reg [21:0] tag_2_0; // @[playground/src/noop/dcache.scala 88:26]
  reg [21:0] tag_2_1; // @[playground/src/noop/dcache.scala 88:26]
  reg [21:0] tag_2_2; // @[playground/src/noop/dcache.scala 88:26]
  reg [21:0] tag_2_3; // @[playground/src/noop/dcache.scala 88:26]
  reg [21:0] tag_2_4; // @[playground/src/noop/dcache.scala 88:26]
  reg [21:0] tag_2_5; // @[playground/src/noop/dcache.scala 88:26]
  reg [21:0] tag_2_6; // @[playground/src/noop/dcache.scala 88:26]
  reg [21:0] tag_2_7; // @[playground/src/noop/dcache.scala 88:26]
  reg [21:0] tag_2_8; // @[playground/src/noop/dcache.scala 88:26]
  reg [21:0] tag_2_9; // @[playground/src/noop/dcache.scala 88:26]
  reg [21:0] tag_2_10; // @[playground/src/noop/dcache.scala 88:26]
  reg [21:0] tag_2_11; // @[playground/src/noop/dcache.scala 88:26]
  reg [21:0] tag_2_12; // @[playground/src/noop/dcache.scala 88:26]
  reg [21:0] tag_2_13; // @[playground/src/noop/dcache.scala 88:26]
  reg [21:0] tag_2_14; // @[playground/src/noop/dcache.scala 88:26]
  reg [21:0] tag_2_15; // @[playground/src/noop/dcache.scala 88:26]
  reg [21:0] tag_3_0; // @[playground/src/noop/dcache.scala 88:26]
  reg [21:0] tag_3_1; // @[playground/src/noop/dcache.scala 88:26]
  reg [21:0] tag_3_2; // @[playground/src/noop/dcache.scala 88:26]
  reg [21:0] tag_3_3; // @[playground/src/noop/dcache.scala 88:26]
  reg [21:0] tag_3_4; // @[playground/src/noop/dcache.scala 88:26]
  reg [21:0] tag_3_5; // @[playground/src/noop/dcache.scala 88:26]
  reg [21:0] tag_3_6; // @[playground/src/noop/dcache.scala 88:26]
  reg [21:0] tag_3_7; // @[playground/src/noop/dcache.scala 88:26]
  reg [21:0] tag_3_8; // @[playground/src/noop/dcache.scala 88:26]
  reg [21:0] tag_3_9; // @[playground/src/noop/dcache.scala 88:26]
  reg [21:0] tag_3_10; // @[playground/src/noop/dcache.scala 88:26]
  reg [21:0] tag_3_11; // @[playground/src/noop/dcache.scala 88:26]
  reg [21:0] tag_3_12; // @[playground/src/noop/dcache.scala 88:26]
  reg [21:0] tag_3_13; // @[playground/src/noop/dcache.scala 88:26]
  reg [21:0] tag_3_14; // @[playground/src/noop/dcache.scala 88:26]
  reg [21:0] tag_3_15; // @[playground/src/noop/dcache.scala 88:26]
  reg  valid_0_0; // @[playground/src/noop/dcache.scala 89:26]
  reg  valid_0_1; // @[playground/src/noop/dcache.scala 89:26]
  reg  valid_0_2; // @[playground/src/noop/dcache.scala 89:26]
  reg  valid_0_3; // @[playground/src/noop/dcache.scala 89:26]
  reg  valid_0_4; // @[playground/src/noop/dcache.scala 89:26]
  reg  valid_0_5; // @[playground/src/noop/dcache.scala 89:26]
  reg  valid_0_6; // @[playground/src/noop/dcache.scala 89:26]
  reg  valid_0_7; // @[playground/src/noop/dcache.scala 89:26]
  reg  valid_0_8; // @[playground/src/noop/dcache.scala 89:26]
  reg  valid_0_9; // @[playground/src/noop/dcache.scala 89:26]
  reg  valid_0_10; // @[playground/src/noop/dcache.scala 89:26]
  reg  valid_0_11; // @[playground/src/noop/dcache.scala 89:26]
  reg  valid_0_12; // @[playground/src/noop/dcache.scala 89:26]
  reg  valid_0_13; // @[playground/src/noop/dcache.scala 89:26]
  reg  valid_0_14; // @[playground/src/noop/dcache.scala 89:26]
  reg  valid_0_15; // @[playground/src/noop/dcache.scala 89:26]
  reg  valid_1_0; // @[playground/src/noop/dcache.scala 89:26]
  reg  valid_1_1; // @[playground/src/noop/dcache.scala 89:26]
  reg  valid_1_2; // @[playground/src/noop/dcache.scala 89:26]
  reg  valid_1_3; // @[playground/src/noop/dcache.scala 89:26]
  reg  valid_1_4; // @[playground/src/noop/dcache.scala 89:26]
  reg  valid_1_5; // @[playground/src/noop/dcache.scala 89:26]
  reg  valid_1_6; // @[playground/src/noop/dcache.scala 89:26]
  reg  valid_1_7; // @[playground/src/noop/dcache.scala 89:26]
  reg  valid_1_8; // @[playground/src/noop/dcache.scala 89:26]
  reg  valid_1_9; // @[playground/src/noop/dcache.scala 89:26]
  reg  valid_1_10; // @[playground/src/noop/dcache.scala 89:26]
  reg  valid_1_11; // @[playground/src/noop/dcache.scala 89:26]
  reg  valid_1_12; // @[playground/src/noop/dcache.scala 89:26]
  reg  valid_1_13; // @[playground/src/noop/dcache.scala 89:26]
  reg  valid_1_14; // @[playground/src/noop/dcache.scala 89:26]
  reg  valid_1_15; // @[playground/src/noop/dcache.scala 89:26]
  reg  valid_2_0; // @[playground/src/noop/dcache.scala 89:26]
  reg  valid_2_1; // @[playground/src/noop/dcache.scala 89:26]
  reg  valid_2_2; // @[playground/src/noop/dcache.scala 89:26]
  reg  valid_2_3; // @[playground/src/noop/dcache.scala 89:26]
  reg  valid_2_4; // @[playground/src/noop/dcache.scala 89:26]
  reg  valid_2_5; // @[playground/src/noop/dcache.scala 89:26]
  reg  valid_2_6; // @[playground/src/noop/dcache.scala 89:26]
  reg  valid_2_7; // @[playground/src/noop/dcache.scala 89:26]
  reg  valid_2_8; // @[playground/src/noop/dcache.scala 89:26]
  reg  valid_2_9; // @[playground/src/noop/dcache.scala 89:26]
  reg  valid_2_10; // @[playground/src/noop/dcache.scala 89:26]
  reg  valid_2_11; // @[playground/src/noop/dcache.scala 89:26]
  reg  valid_2_12; // @[playground/src/noop/dcache.scala 89:26]
  reg  valid_2_13; // @[playground/src/noop/dcache.scala 89:26]
  reg  valid_2_14; // @[playground/src/noop/dcache.scala 89:26]
  reg  valid_2_15; // @[playground/src/noop/dcache.scala 89:26]
  reg  valid_3_0; // @[playground/src/noop/dcache.scala 89:26]
  reg  valid_3_1; // @[playground/src/noop/dcache.scala 89:26]
  reg  valid_3_2; // @[playground/src/noop/dcache.scala 89:26]
  reg  valid_3_3; // @[playground/src/noop/dcache.scala 89:26]
  reg  valid_3_4; // @[playground/src/noop/dcache.scala 89:26]
  reg  valid_3_5; // @[playground/src/noop/dcache.scala 89:26]
  reg  valid_3_6; // @[playground/src/noop/dcache.scala 89:26]
  reg  valid_3_7; // @[playground/src/noop/dcache.scala 89:26]
  reg  valid_3_8; // @[playground/src/noop/dcache.scala 89:26]
  reg  valid_3_9; // @[playground/src/noop/dcache.scala 89:26]
  reg  valid_3_10; // @[playground/src/noop/dcache.scala 89:26]
  reg  valid_3_11; // @[playground/src/noop/dcache.scala 89:26]
  reg  valid_3_12; // @[playground/src/noop/dcache.scala 89:26]
  reg  valid_3_13; // @[playground/src/noop/dcache.scala 89:26]
  reg  valid_3_14; // @[playground/src/noop/dcache.scala 89:26]
  reg  valid_3_15; // @[playground/src/noop/dcache.scala 89:26]
  reg  dirty_0_0; // @[playground/src/noop/dcache.scala 90:26]
  reg  dirty_0_1; // @[playground/src/noop/dcache.scala 90:26]
  reg  dirty_0_2; // @[playground/src/noop/dcache.scala 90:26]
  reg  dirty_0_3; // @[playground/src/noop/dcache.scala 90:26]
  reg  dirty_0_4; // @[playground/src/noop/dcache.scala 90:26]
  reg  dirty_0_5; // @[playground/src/noop/dcache.scala 90:26]
  reg  dirty_0_6; // @[playground/src/noop/dcache.scala 90:26]
  reg  dirty_0_7; // @[playground/src/noop/dcache.scala 90:26]
  reg  dirty_0_8; // @[playground/src/noop/dcache.scala 90:26]
  reg  dirty_0_9; // @[playground/src/noop/dcache.scala 90:26]
  reg  dirty_0_10; // @[playground/src/noop/dcache.scala 90:26]
  reg  dirty_0_11; // @[playground/src/noop/dcache.scala 90:26]
  reg  dirty_0_12; // @[playground/src/noop/dcache.scala 90:26]
  reg  dirty_0_13; // @[playground/src/noop/dcache.scala 90:26]
  reg  dirty_0_14; // @[playground/src/noop/dcache.scala 90:26]
  reg  dirty_0_15; // @[playground/src/noop/dcache.scala 90:26]
  reg  dirty_1_0; // @[playground/src/noop/dcache.scala 90:26]
  reg  dirty_1_1; // @[playground/src/noop/dcache.scala 90:26]
  reg  dirty_1_2; // @[playground/src/noop/dcache.scala 90:26]
  reg  dirty_1_3; // @[playground/src/noop/dcache.scala 90:26]
  reg  dirty_1_4; // @[playground/src/noop/dcache.scala 90:26]
  reg  dirty_1_5; // @[playground/src/noop/dcache.scala 90:26]
  reg  dirty_1_6; // @[playground/src/noop/dcache.scala 90:26]
  reg  dirty_1_7; // @[playground/src/noop/dcache.scala 90:26]
  reg  dirty_1_8; // @[playground/src/noop/dcache.scala 90:26]
  reg  dirty_1_9; // @[playground/src/noop/dcache.scala 90:26]
  reg  dirty_1_10; // @[playground/src/noop/dcache.scala 90:26]
  reg  dirty_1_11; // @[playground/src/noop/dcache.scala 90:26]
  reg  dirty_1_12; // @[playground/src/noop/dcache.scala 90:26]
  reg  dirty_1_13; // @[playground/src/noop/dcache.scala 90:26]
  reg  dirty_1_14; // @[playground/src/noop/dcache.scala 90:26]
  reg  dirty_1_15; // @[playground/src/noop/dcache.scala 90:26]
  reg  dirty_2_0; // @[playground/src/noop/dcache.scala 90:26]
  reg  dirty_2_1; // @[playground/src/noop/dcache.scala 90:26]
  reg  dirty_2_2; // @[playground/src/noop/dcache.scala 90:26]
  reg  dirty_2_3; // @[playground/src/noop/dcache.scala 90:26]
  reg  dirty_2_4; // @[playground/src/noop/dcache.scala 90:26]
  reg  dirty_2_5; // @[playground/src/noop/dcache.scala 90:26]
  reg  dirty_2_6; // @[playground/src/noop/dcache.scala 90:26]
  reg  dirty_2_7; // @[playground/src/noop/dcache.scala 90:26]
  reg  dirty_2_8; // @[playground/src/noop/dcache.scala 90:26]
  reg  dirty_2_9; // @[playground/src/noop/dcache.scala 90:26]
  reg  dirty_2_10; // @[playground/src/noop/dcache.scala 90:26]
  reg  dirty_2_11; // @[playground/src/noop/dcache.scala 90:26]
  reg  dirty_2_12; // @[playground/src/noop/dcache.scala 90:26]
  reg  dirty_2_13; // @[playground/src/noop/dcache.scala 90:26]
  reg  dirty_2_14; // @[playground/src/noop/dcache.scala 90:26]
  reg  dirty_2_15; // @[playground/src/noop/dcache.scala 90:26]
  reg  dirty_3_0; // @[playground/src/noop/dcache.scala 90:26]
  reg  dirty_3_1; // @[playground/src/noop/dcache.scala 90:26]
  reg  dirty_3_2; // @[playground/src/noop/dcache.scala 90:26]
  reg  dirty_3_3; // @[playground/src/noop/dcache.scala 90:26]
  reg  dirty_3_4; // @[playground/src/noop/dcache.scala 90:26]
  reg  dirty_3_5; // @[playground/src/noop/dcache.scala 90:26]
  reg  dirty_3_6; // @[playground/src/noop/dcache.scala 90:26]
  reg  dirty_3_7; // @[playground/src/noop/dcache.scala 90:26]
  reg  dirty_3_8; // @[playground/src/noop/dcache.scala 90:26]
  reg  dirty_3_9; // @[playground/src/noop/dcache.scala 90:26]
  reg  dirty_3_10; // @[playground/src/noop/dcache.scala 90:26]
  reg  dirty_3_11; // @[playground/src/noop/dcache.scala 90:26]
  reg  dirty_3_12; // @[playground/src/noop/dcache.scala 90:26]
  reg  dirty_3_13; // @[playground/src/noop/dcache.scala 90:26]
  reg  dirty_3_14; // @[playground/src/noop/dcache.scala 90:26]
  reg  dirty_3_15; // @[playground/src/noop/dcache.scala 90:26]
  reg  wait_r; // @[playground/src/noop/dcache.scala 95:30]
  reg  valid_r; // @[playground/src/noop/dcache.scala 96:30]
  reg  flush_r; // @[playground/src/noop/dcache.scala 97:30]
  reg [4:0] mode_r; // @[playground/src/noop/dcache.scala 98:30]
  reg [63:0] wdata_r; // @[playground/src/noop/dcache.scala 99:30]
  reg [4:0] amo_r; // @[playground/src/noop/dcache.scala 100:30]
  wire  _valid_in_T = io_dcRW_dc_mode != 5'h0; // @[playground/src/noop/dcache.scala 102:40]
  wire  valid_in = io_dcRW_dc_mode != 5'h0 & ~io_flush; // @[playground/src/noop/dcache.scala 102:54]
  wire  hs_in = _valid_in_T & io_dcRW_ready; // @[playground/src/noop/dcache.scala 103:52]
  wire  _io_dcRW_ready_T = ~wait_r; // @[playground/src/noop/dcache.scala 104:34]
  reg [31:0] addr_r; // @[playground/src/noop/dcache.scala 107:34]
  wire [31:0] cur_addr = hs_in ? io_dcRW_addr : addr_r; // @[playground/src/noop/dcache.scala 108:30]
  reg [1:0] matchWay_r; // @[playground/src/noop/dcache.scala 109:34]
  reg [2:0] offset; // @[playground/src/noop/dcache.scala 110:34]
  reg [63:0] rdatabuf; // @[playground/src/noop/dcache.scala 111:34]
  wire [3:0] blockIdx = cur_addr[9:6]; // @[playground/src/noop/dcache.scala 112:35]
  reg [3:0] blockIdx_r; // @[playground/src/noop/dcache.scala 113:34]
  wire [21:0] cur_tag = cur_addr[31:10]; // @[playground/src/noop/dcache.scala 114:35]
  wire [21:0] _GEN_1 = 4'h1 == blockIdx ? tag_0_1 : tag_0_0; // @[playground/src/noop/dcache.scala 115:{85,85}]
  wire [21:0] _GEN_2 = 4'h2 == blockIdx ? tag_0_2 : _GEN_1; // @[playground/src/noop/dcache.scala 115:{85,85}]
  wire [21:0] _GEN_3 = 4'h3 == blockIdx ? tag_0_3 : _GEN_2; // @[playground/src/noop/dcache.scala 115:{85,85}]
  wire [21:0] _GEN_4 = 4'h4 == blockIdx ? tag_0_4 : _GEN_3; // @[playground/src/noop/dcache.scala 115:{85,85}]
  wire [21:0] _GEN_5 = 4'h5 == blockIdx ? tag_0_5 : _GEN_4; // @[playground/src/noop/dcache.scala 115:{85,85}]
  wire [21:0] _GEN_6 = 4'h6 == blockIdx ? tag_0_6 : _GEN_5; // @[playground/src/noop/dcache.scala 115:{85,85}]
  wire [21:0] _GEN_7 = 4'h7 == blockIdx ? tag_0_7 : _GEN_6; // @[playground/src/noop/dcache.scala 115:{85,85}]
  wire [21:0] _GEN_8 = 4'h8 == blockIdx ? tag_0_8 : _GEN_7; // @[playground/src/noop/dcache.scala 115:{85,85}]
  wire [21:0] _GEN_9 = 4'h9 == blockIdx ? tag_0_9 : _GEN_8; // @[playground/src/noop/dcache.scala 115:{85,85}]
  wire [21:0] _GEN_10 = 4'ha == blockIdx ? tag_0_10 : _GEN_9; // @[playground/src/noop/dcache.scala 115:{85,85}]
  wire [21:0] _GEN_11 = 4'hb == blockIdx ? tag_0_11 : _GEN_10; // @[playground/src/noop/dcache.scala 115:{85,85}]
  wire [21:0] _GEN_12 = 4'hc == blockIdx ? tag_0_12 : _GEN_11; // @[playground/src/noop/dcache.scala 115:{85,85}]
  wire [21:0] _GEN_13 = 4'hd == blockIdx ? tag_0_13 : _GEN_12; // @[playground/src/noop/dcache.scala 115:{85,85}]
  wire [21:0] _GEN_14 = 4'he == blockIdx ? tag_0_14 : _GEN_13; // @[playground/src/noop/dcache.scala 115:{85,85}]
  wire [21:0] _GEN_15 = 4'hf == blockIdx ? tag_0_15 : _GEN_14; // @[playground/src/noop/dcache.scala 115:{85,85}]
  wire  _GEN_17 = 4'h1 == blockIdx ? valid_0_1 : valid_0_0; // @[playground/src/noop/dcache.scala 115:{97,97}]
  wire  _GEN_18 = 4'h2 == blockIdx ? valid_0_2 : _GEN_17; // @[playground/src/noop/dcache.scala 115:{97,97}]
  wire  _GEN_19 = 4'h3 == blockIdx ? valid_0_3 : _GEN_18; // @[playground/src/noop/dcache.scala 115:{97,97}]
  wire  _GEN_20 = 4'h4 == blockIdx ? valid_0_4 : _GEN_19; // @[playground/src/noop/dcache.scala 115:{97,97}]
  wire  _GEN_21 = 4'h5 == blockIdx ? valid_0_5 : _GEN_20; // @[playground/src/noop/dcache.scala 115:{97,97}]
  wire  _GEN_22 = 4'h6 == blockIdx ? valid_0_6 : _GEN_21; // @[playground/src/noop/dcache.scala 115:{97,97}]
  wire  _GEN_23 = 4'h7 == blockIdx ? valid_0_7 : _GEN_22; // @[playground/src/noop/dcache.scala 115:{97,97}]
  wire  _GEN_24 = 4'h8 == blockIdx ? valid_0_8 : _GEN_23; // @[playground/src/noop/dcache.scala 115:{97,97}]
  wire  _GEN_25 = 4'h9 == blockIdx ? valid_0_9 : _GEN_24; // @[playground/src/noop/dcache.scala 115:{97,97}]
  wire  _GEN_26 = 4'ha == blockIdx ? valid_0_10 : _GEN_25; // @[playground/src/noop/dcache.scala 115:{97,97}]
  wire  _GEN_27 = 4'hb == blockIdx ? valid_0_11 : _GEN_26; // @[playground/src/noop/dcache.scala 115:{97,97}]
  wire  _GEN_28 = 4'hc == blockIdx ? valid_0_12 : _GEN_27; // @[playground/src/noop/dcache.scala 115:{97,97}]
  wire  _GEN_29 = 4'hd == blockIdx ? valid_0_13 : _GEN_28; // @[playground/src/noop/dcache.scala 115:{97,97}]
  wire  _GEN_30 = 4'he == blockIdx ? valid_0_14 : _GEN_29; // @[playground/src/noop/dcache.scala 115:{97,97}]
  wire  _GEN_31 = 4'hf == blockIdx ? valid_0_15 : _GEN_30; // @[playground/src/noop/dcache.scala 115:{97,97}]
  wire  cache_hit_vec_0 = _GEN_15 == cur_tag & _GEN_31; // @[playground/src/noop/dcache.scala 115:97]
  wire [21:0] _GEN_33 = 4'h1 == blockIdx ? tag_1_1 : tag_1_0; // @[playground/src/noop/dcache.scala 115:{85,85}]
  wire [21:0] _GEN_34 = 4'h2 == blockIdx ? tag_1_2 : _GEN_33; // @[playground/src/noop/dcache.scala 115:{85,85}]
  wire [21:0] _GEN_35 = 4'h3 == blockIdx ? tag_1_3 : _GEN_34; // @[playground/src/noop/dcache.scala 115:{85,85}]
  wire [21:0] _GEN_36 = 4'h4 == blockIdx ? tag_1_4 : _GEN_35; // @[playground/src/noop/dcache.scala 115:{85,85}]
  wire [21:0] _GEN_37 = 4'h5 == blockIdx ? tag_1_5 : _GEN_36; // @[playground/src/noop/dcache.scala 115:{85,85}]
  wire [21:0] _GEN_38 = 4'h6 == blockIdx ? tag_1_6 : _GEN_37; // @[playground/src/noop/dcache.scala 115:{85,85}]
  wire [21:0] _GEN_39 = 4'h7 == blockIdx ? tag_1_7 : _GEN_38; // @[playground/src/noop/dcache.scala 115:{85,85}]
  wire [21:0] _GEN_40 = 4'h8 == blockIdx ? tag_1_8 : _GEN_39; // @[playground/src/noop/dcache.scala 115:{85,85}]
  wire [21:0] _GEN_41 = 4'h9 == blockIdx ? tag_1_9 : _GEN_40; // @[playground/src/noop/dcache.scala 115:{85,85}]
  wire [21:0] _GEN_42 = 4'ha == blockIdx ? tag_1_10 : _GEN_41; // @[playground/src/noop/dcache.scala 115:{85,85}]
  wire [21:0] _GEN_43 = 4'hb == blockIdx ? tag_1_11 : _GEN_42; // @[playground/src/noop/dcache.scala 115:{85,85}]
  wire [21:0] _GEN_44 = 4'hc == blockIdx ? tag_1_12 : _GEN_43; // @[playground/src/noop/dcache.scala 115:{85,85}]
  wire [21:0] _GEN_45 = 4'hd == blockIdx ? tag_1_13 : _GEN_44; // @[playground/src/noop/dcache.scala 115:{85,85}]
  wire [21:0] _GEN_46 = 4'he == blockIdx ? tag_1_14 : _GEN_45; // @[playground/src/noop/dcache.scala 115:{85,85}]
  wire [21:0] _GEN_47 = 4'hf == blockIdx ? tag_1_15 : _GEN_46; // @[playground/src/noop/dcache.scala 115:{85,85}]
  wire  _GEN_49 = 4'h1 == blockIdx ? valid_1_1 : valid_1_0; // @[playground/src/noop/dcache.scala 115:{97,97}]
  wire  _GEN_50 = 4'h2 == blockIdx ? valid_1_2 : _GEN_49; // @[playground/src/noop/dcache.scala 115:{97,97}]
  wire  _GEN_51 = 4'h3 == blockIdx ? valid_1_3 : _GEN_50; // @[playground/src/noop/dcache.scala 115:{97,97}]
  wire  _GEN_52 = 4'h4 == blockIdx ? valid_1_4 : _GEN_51; // @[playground/src/noop/dcache.scala 115:{97,97}]
  wire  _GEN_53 = 4'h5 == blockIdx ? valid_1_5 : _GEN_52; // @[playground/src/noop/dcache.scala 115:{97,97}]
  wire  _GEN_54 = 4'h6 == blockIdx ? valid_1_6 : _GEN_53; // @[playground/src/noop/dcache.scala 115:{97,97}]
  wire  _GEN_55 = 4'h7 == blockIdx ? valid_1_7 : _GEN_54; // @[playground/src/noop/dcache.scala 115:{97,97}]
  wire  _GEN_56 = 4'h8 == blockIdx ? valid_1_8 : _GEN_55; // @[playground/src/noop/dcache.scala 115:{97,97}]
  wire  _GEN_57 = 4'h9 == blockIdx ? valid_1_9 : _GEN_56; // @[playground/src/noop/dcache.scala 115:{97,97}]
  wire  _GEN_58 = 4'ha == blockIdx ? valid_1_10 : _GEN_57; // @[playground/src/noop/dcache.scala 115:{97,97}]
  wire  _GEN_59 = 4'hb == blockIdx ? valid_1_11 : _GEN_58; // @[playground/src/noop/dcache.scala 115:{97,97}]
  wire  _GEN_60 = 4'hc == blockIdx ? valid_1_12 : _GEN_59; // @[playground/src/noop/dcache.scala 115:{97,97}]
  wire  _GEN_61 = 4'hd == blockIdx ? valid_1_13 : _GEN_60; // @[playground/src/noop/dcache.scala 115:{97,97}]
  wire  _GEN_62 = 4'he == blockIdx ? valid_1_14 : _GEN_61; // @[playground/src/noop/dcache.scala 115:{97,97}]
  wire  _GEN_63 = 4'hf == blockIdx ? valid_1_15 : _GEN_62; // @[playground/src/noop/dcache.scala 115:{97,97}]
  wire  cache_hit_vec_1 = _GEN_47 == cur_tag & _GEN_63; // @[playground/src/noop/dcache.scala 115:97]
  wire [21:0] _GEN_65 = 4'h1 == blockIdx ? tag_2_1 : tag_2_0; // @[playground/src/noop/dcache.scala 115:{85,85}]
  wire [21:0] _GEN_66 = 4'h2 == blockIdx ? tag_2_2 : _GEN_65; // @[playground/src/noop/dcache.scala 115:{85,85}]
  wire [21:0] _GEN_67 = 4'h3 == blockIdx ? tag_2_3 : _GEN_66; // @[playground/src/noop/dcache.scala 115:{85,85}]
  wire [21:0] _GEN_68 = 4'h4 == blockIdx ? tag_2_4 : _GEN_67; // @[playground/src/noop/dcache.scala 115:{85,85}]
  wire [21:0] _GEN_69 = 4'h5 == blockIdx ? tag_2_5 : _GEN_68; // @[playground/src/noop/dcache.scala 115:{85,85}]
  wire [21:0] _GEN_70 = 4'h6 == blockIdx ? tag_2_6 : _GEN_69; // @[playground/src/noop/dcache.scala 115:{85,85}]
  wire [21:0] _GEN_71 = 4'h7 == blockIdx ? tag_2_7 : _GEN_70; // @[playground/src/noop/dcache.scala 115:{85,85}]
  wire [21:0] _GEN_72 = 4'h8 == blockIdx ? tag_2_8 : _GEN_71; // @[playground/src/noop/dcache.scala 115:{85,85}]
  wire [21:0] _GEN_73 = 4'h9 == blockIdx ? tag_2_9 : _GEN_72; // @[playground/src/noop/dcache.scala 115:{85,85}]
  wire [21:0] _GEN_74 = 4'ha == blockIdx ? tag_2_10 : _GEN_73; // @[playground/src/noop/dcache.scala 115:{85,85}]
  wire [21:0] _GEN_75 = 4'hb == blockIdx ? tag_2_11 : _GEN_74; // @[playground/src/noop/dcache.scala 115:{85,85}]
  wire [21:0] _GEN_76 = 4'hc == blockIdx ? tag_2_12 : _GEN_75; // @[playground/src/noop/dcache.scala 115:{85,85}]
  wire [21:0] _GEN_77 = 4'hd == blockIdx ? tag_2_13 : _GEN_76; // @[playground/src/noop/dcache.scala 115:{85,85}]
  wire [21:0] _GEN_78 = 4'he == blockIdx ? tag_2_14 : _GEN_77; // @[playground/src/noop/dcache.scala 115:{85,85}]
  wire [21:0] _GEN_79 = 4'hf == blockIdx ? tag_2_15 : _GEN_78; // @[playground/src/noop/dcache.scala 115:{85,85}]
  wire  _GEN_81 = 4'h1 == blockIdx ? valid_2_1 : valid_2_0; // @[playground/src/noop/dcache.scala 115:{97,97}]
  wire  _GEN_82 = 4'h2 == blockIdx ? valid_2_2 : _GEN_81; // @[playground/src/noop/dcache.scala 115:{97,97}]
  wire  _GEN_83 = 4'h3 == blockIdx ? valid_2_3 : _GEN_82; // @[playground/src/noop/dcache.scala 115:{97,97}]
  wire  _GEN_84 = 4'h4 == blockIdx ? valid_2_4 : _GEN_83; // @[playground/src/noop/dcache.scala 115:{97,97}]
  wire  _GEN_85 = 4'h5 == blockIdx ? valid_2_5 : _GEN_84; // @[playground/src/noop/dcache.scala 115:{97,97}]
  wire  _GEN_86 = 4'h6 == blockIdx ? valid_2_6 : _GEN_85; // @[playground/src/noop/dcache.scala 115:{97,97}]
  wire  _GEN_87 = 4'h7 == blockIdx ? valid_2_7 : _GEN_86; // @[playground/src/noop/dcache.scala 115:{97,97}]
  wire  _GEN_88 = 4'h8 == blockIdx ? valid_2_8 : _GEN_87; // @[playground/src/noop/dcache.scala 115:{97,97}]
  wire  _GEN_89 = 4'h9 == blockIdx ? valid_2_9 : _GEN_88; // @[playground/src/noop/dcache.scala 115:{97,97}]
  wire  _GEN_90 = 4'ha == blockIdx ? valid_2_10 : _GEN_89; // @[playground/src/noop/dcache.scala 115:{97,97}]
  wire  _GEN_91 = 4'hb == blockIdx ? valid_2_11 : _GEN_90; // @[playground/src/noop/dcache.scala 115:{97,97}]
  wire  _GEN_92 = 4'hc == blockIdx ? valid_2_12 : _GEN_91; // @[playground/src/noop/dcache.scala 115:{97,97}]
  wire  _GEN_93 = 4'hd == blockIdx ? valid_2_13 : _GEN_92; // @[playground/src/noop/dcache.scala 115:{97,97}]
  wire  _GEN_94 = 4'he == blockIdx ? valid_2_14 : _GEN_93; // @[playground/src/noop/dcache.scala 115:{97,97}]
  wire  _GEN_95 = 4'hf == blockIdx ? valid_2_15 : _GEN_94; // @[playground/src/noop/dcache.scala 115:{97,97}]
  wire  cache_hit_vec_2 = _GEN_79 == cur_tag & _GEN_95; // @[playground/src/noop/dcache.scala 115:97]
  wire [21:0] _GEN_97 = 4'h1 == blockIdx ? tag_3_1 : tag_3_0; // @[playground/src/noop/dcache.scala 115:{85,85}]
  wire [21:0] _GEN_98 = 4'h2 == blockIdx ? tag_3_2 : _GEN_97; // @[playground/src/noop/dcache.scala 115:{85,85}]
  wire [21:0] _GEN_99 = 4'h3 == blockIdx ? tag_3_3 : _GEN_98; // @[playground/src/noop/dcache.scala 115:{85,85}]
  wire [21:0] _GEN_100 = 4'h4 == blockIdx ? tag_3_4 : _GEN_99; // @[playground/src/noop/dcache.scala 115:{85,85}]
  wire [21:0] _GEN_101 = 4'h5 == blockIdx ? tag_3_5 : _GEN_100; // @[playground/src/noop/dcache.scala 115:{85,85}]
  wire [21:0] _GEN_102 = 4'h6 == blockIdx ? tag_3_6 : _GEN_101; // @[playground/src/noop/dcache.scala 115:{85,85}]
  wire [21:0] _GEN_103 = 4'h7 == blockIdx ? tag_3_7 : _GEN_102; // @[playground/src/noop/dcache.scala 115:{85,85}]
  wire [21:0] _GEN_104 = 4'h8 == blockIdx ? tag_3_8 : _GEN_103; // @[playground/src/noop/dcache.scala 115:{85,85}]
  wire [21:0] _GEN_105 = 4'h9 == blockIdx ? tag_3_9 : _GEN_104; // @[playground/src/noop/dcache.scala 115:{85,85}]
  wire [21:0] _GEN_106 = 4'ha == blockIdx ? tag_3_10 : _GEN_105; // @[playground/src/noop/dcache.scala 115:{85,85}]
  wire [21:0] _GEN_107 = 4'hb == blockIdx ? tag_3_11 : _GEN_106; // @[playground/src/noop/dcache.scala 115:{85,85}]
  wire [21:0] _GEN_108 = 4'hc == blockIdx ? tag_3_12 : _GEN_107; // @[playground/src/noop/dcache.scala 115:{85,85}]
  wire [21:0] _GEN_109 = 4'hd == blockIdx ? tag_3_13 : _GEN_108; // @[playground/src/noop/dcache.scala 115:{85,85}]
  wire [21:0] _GEN_110 = 4'he == blockIdx ? tag_3_14 : _GEN_109; // @[playground/src/noop/dcache.scala 115:{85,85}]
  wire [21:0] _GEN_111 = 4'hf == blockIdx ? tag_3_15 : _GEN_110; // @[playground/src/noop/dcache.scala 115:{85,85}]
  wire  _GEN_113 = 4'h1 == blockIdx ? valid_3_1 : valid_3_0; // @[playground/src/noop/dcache.scala 115:{97,97}]
  wire  _GEN_114 = 4'h2 == blockIdx ? valid_3_2 : _GEN_113; // @[playground/src/noop/dcache.scala 115:{97,97}]
  wire  _GEN_115 = 4'h3 == blockIdx ? valid_3_3 : _GEN_114; // @[playground/src/noop/dcache.scala 115:{97,97}]
  wire  _GEN_116 = 4'h4 == blockIdx ? valid_3_4 : _GEN_115; // @[playground/src/noop/dcache.scala 115:{97,97}]
  wire  _GEN_117 = 4'h5 == blockIdx ? valid_3_5 : _GEN_116; // @[playground/src/noop/dcache.scala 115:{97,97}]
  wire  _GEN_118 = 4'h6 == blockIdx ? valid_3_6 : _GEN_117; // @[playground/src/noop/dcache.scala 115:{97,97}]
  wire  _GEN_119 = 4'h7 == blockIdx ? valid_3_7 : _GEN_118; // @[playground/src/noop/dcache.scala 115:{97,97}]
  wire  _GEN_120 = 4'h8 == blockIdx ? valid_3_8 : _GEN_119; // @[playground/src/noop/dcache.scala 115:{97,97}]
  wire  _GEN_121 = 4'h9 == blockIdx ? valid_3_9 : _GEN_120; // @[playground/src/noop/dcache.scala 115:{97,97}]
  wire  _GEN_122 = 4'ha == blockIdx ? valid_3_10 : _GEN_121; // @[playground/src/noop/dcache.scala 115:{97,97}]
  wire  _GEN_123 = 4'hb == blockIdx ? valid_3_11 : _GEN_122; // @[playground/src/noop/dcache.scala 115:{97,97}]
  wire  _GEN_124 = 4'hc == blockIdx ? valid_3_12 : _GEN_123; // @[playground/src/noop/dcache.scala 115:{97,97}]
  wire  _GEN_125 = 4'hd == blockIdx ? valid_3_13 : _GEN_124; // @[playground/src/noop/dcache.scala 115:{97,97}]
  wire  _GEN_126 = 4'he == blockIdx ? valid_3_14 : _GEN_125; // @[playground/src/noop/dcache.scala 115:{97,97}]
  wire  _GEN_127 = 4'hf == blockIdx ? valid_3_15 : _GEN_126; // @[playground/src/noop/dcache.scala 115:{97,97}]
  wire  cache_hit_vec_3 = _GEN_111 == cur_tag & _GEN_127; // @[playground/src/noop/dcache.scala 115:97]
  wire [3:0] _cacheHit_T = {cache_hit_vec_3,cache_hit_vec_2,cache_hit_vec_1,cache_hit_vec_0}; // @[playground/src/noop/dcache.scala 116:41]
  wire  cacheHit = |_cacheHit_T; // @[playground/src/noop/dcache.scala 116:48]
  wire [1:0] matchWay_hi_1 = _cacheHit_T[3:2]; // @[src/main/scala/chisel3/util/OneHot.scala 30:18]
  wire [1:0] matchWay_lo_1 = _cacheHit_T[1:0]; // @[src/main/scala/chisel3/util/OneHot.scala 31:18]
  wire [1:0] _matchWay_T_2 = matchWay_hi_1 | matchWay_lo_1; // @[src/main/scala/chisel3/util/OneHot.scala 32:28]
  wire [1:0] _matchWay_T_4 = {|matchWay_hi_1,_matchWay_T_2[1]}; // @[src/main/scala/chisel3/util/OneHot.scala 32:10]
  wire [1:0] _matchWay_T_5 = {matchWay_prng_io_out_1,matchWay_prng_io_out_0}; // @[src/main/scala/chisel3/util/random/PRNG.scala 95:17]
  wire [1:0] _matchWay_T_6 = hs_in ? _matchWay_T_5 : matchWay_r; // @[playground/src/noop/dcache.scala 117:69]
  wire [1:0] matchWay = cacheHit ? _matchWay_T_4 : _matchWay_T_6; // @[playground/src/noop/dcache.scala 117:30]
  wire [1:0] _GEN_129 = hs_in ? matchWay : matchWay_r; // @[playground/src/noop/dcache.scala 119:16 121:20 109:34]
  wire [4:0] _GEN_130 = hs_in ? io_dcRW_dc_mode : mode_r; // @[playground/src/noop/dcache.scala 119:16 122:17 98:30]
  wire [63:0] _GEN_131 = hs_in ? io_dcRW_wdata : wdata_r; // @[playground/src/noop/dcache.scala 119:16 123:17 99:30]
  wire [3:0] _GEN_133 = hs_in ? io_dcRW_addr[9:6] : blockIdx_r; // @[playground/src/noop/dcache.scala 119:16 125:20 113:34]
  wire  _GEN_134 = io_flush | flush_r; // @[playground/src/noop/dcache.scala 128:19 129:17 97:30]
  wire  _GEN_136 = valid_0_0 & dirty_0_0 ? 1'h0 : 1'h1; // @[playground/src/noop/dcache.scala 137:45 140:28 134:52]
  wire  _T_1 = valid_0_1 & dirty_0_1; // @[playground/src/noop/dcache.scala 137:30]
  wire  _GEN_139 = valid_0_1 & dirty_0_1 ? 1'h0 : _GEN_136; // @[playground/src/noop/dcache.scala 137:45 140:28]
  wire [1:0] _GEN_141 = valid_0_2 & dirty_0_2 ? 2'h2 : {{1'd0}, _T_1}; // @[playground/src/noop/dcache.scala 137:45 139:27]
  wire  _GEN_142 = valid_0_2 & dirty_0_2 ? 1'h0 : _GEN_139; // @[playground/src/noop/dcache.scala 137:45 140:28]
  wire [1:0] _GEN_144 = valid_0_3 & dirty_0_3 ? 2'h3 : _GEN_141; // @[playground/src/noop/dcache.scala 137:45 139:27]
  wire  _GEN_145 = valid_0_3 & dirty_0_3 ? 1'h0 : _GEN_142; // @[playground/src/noop/dcache.scala 137:45 140:28]
  wire [2:0] _GEN_147 = valid_0_4 & dirty_0_4 ? 3'h4 : {{1'd0}, _GEN_144}; // @[playground/src/noop/dcache.scala 137:45 139:27]
  wire  _GEN_148 = valid_0_4 & dirty_0_4 ? 1'h0 : _GEN_145; // @[playground/src/noop/dcache.scala 137:45 140:28]
  wire [2:0] _GEN_150 = valid_0_5 & dirty_0_5 ? 3'h5 : _GEN_147; // @[playground/src/noop/dcache.scala 137:45 139:27]
  wire  _GEN_151 = valid_0_5 & dirty_0_5 ? 1'h0 : _GEN_148; // @[playground/src/noop/dcache.scala 137:45 140:28]
  wire [2:0] _GEN_153 = valid_0_6 & dirty_0_6 ? 3'h6 : _GEN_150; // @[playground/src/noop/dcache.scala 137:45 139:27]
  wire  _GEN_154 = valid_0_6 & dirty_0_6 ? 1'h0 : _GEN_151; // @[playground/src/noop/dcache.scala 137:45 140:28]
  wire [2:0] _GEN_156 = valid_0_7 & dirty_0_7 ? 3'h7 : _GEN_153; // @[playground/src/noop/dcache.scala 137:45 139:27]
  wire  _GEN_157 = valid_0_7 & dirty_0_7 ? 1'h0 : _GEN_154; // @[playground/src/noop/dcache.scala 137:45 140:28]
  wire [3:0] _GEN_159 = valid_0_8 & dirty_0_8 ? 4'h8 : {{1'd0}, _GEN_156}; // @[playground/src/noop/dcache.scala 137:45 139:27]
  wire  _GEN_160 = valid_0_8 & dirty_0_8 ? 1'h0 : _GEN_157; // @[playground/src/noop/dcache.scala 137:45 140:28]
  wire [3:0] _GEN_162 = valid_0_9 & dirty_0_9 ? 4'h9 : _GEN_159; // @[playground/src/noop/dcache.scala 137:45 139:27]
  wire  _GEN_163 = valid_0_9 & dirty_0_9 ? 1'h0 : _GEN_160; // @[playground/src/noop/dcache.scala 137:45 140:28]
  wire [3:0] _GEN_165 = valid_0_10 & dirty_0_10 ? 4'ha : _GEN_162; // @[playground/src/noop/dcache.scala 137:45 139:27]
  wire  _GEN_166 = valid_0_10 & dirty_0_10 ? 1'h0 : _GEN_163; // @[playground/src/noop/dcache.scala 137:45 140:28]
  wire [3:0] _GEN_168 = valid_0_11 & dirty_0_11 ? 4'hb : _GEN_165; // @[playground/src/noop/dcache.scala 137:45 139:27]
  wire  _GEN_169 = valid_0_11 & dirty_0_11 ? 1'h0 : _GEN_166; // @[playground/src/noop/dcache.scala 137:45 140:28]
  wire [3:0] _GEN_171 = valid_0_12 & dirty_0_12 ? 4'hc : _GEN_168; // @[playground/src/noop/dcache.scala 137:45 139:27]
  wire  _GEN_172 = valid_0_12 & dirty_0_12 ? 1'h0 : _GEN_169; // @[playground/src/noop/dcache.scala 137:45 140:28]
  wire [3:0] _GEN_174 = valid_0_13 & dirty_0_13 ? 4'hd : _GEN_171; // @[playground/src/noop/dcache.scala 137:45 139:27]
  wire  _GEN_175 = valid_0_13 & dirty_0_13 ? 1'h0 : _GEN_172; // @[playground/src/noop/dcache.scala 137:45 140:28]
  wire [3:0] _GEN_177 = valid_0_14 & dirty_0_14 ? 4'he : _GEN_174; // @[playground/src/noop/dcache.scala 137:45 139:27]
  wire  _GEN_178 = valid_0_14 & dirty_0_14 ? 1'h0 : _GEN_175; // @[playground/src/noop/dcache.scala 137:45 140:28]
  wire [3:0] _GEN_180 = valid_0_15 & dirty_0_15 ? 4'hf : _GEN_177; // @[playground/src/noop/dcache.scala 137:45 139:27]
  wire  _GEN_181 = valid_0_15 & dirty_0_15 ? 1'h0 : _GEN_178; // @[playground/src/noop/dcache.scala 137:45 140:28]
  wire [3:0] _GEN_183 = valid_1_0 & dirty_1_0 ? 4'h0 : _GEN_180; // @[playground/src/noop/dcache.scala 137:45 139:27]
  wire  _GEN_184 = valid_1_0 & dirty_1_0 ? 1'h0 : _GEN_181; // @[playground/src/noop/dcache.scala 137:45 140:28]
  wire [3:0] _GEN_186 = valid_1_1 & dirty_1_1 ? 4'h1 : _GEN_183; // @[playground/src/noop/dcache.scala 137:45 139:27]
  wire  _GEN_187 = valid_1_1 & dirty_1_1 ? 1'h0 : _GEN_184; // @[playground/src/noop/dcache.scala 137:45 140:28]
  wire [3:0] _GEN_189 = valid_1_2 & dirty_1_2 ? 4'h2 : _GEN_186; // @[playground/src/noop/dcache.scala 137:45 139:27]
  wire  _GEN_190 = valid_1_2 & dirty_1_2 ? 1'h0 : _GEN_187; // @[playground/src/noop/dcache.scala 137:45 140:28]
  wire [3:0] _GEN_192 = valid_1_3 & dirty_1_3 ? 4'h3 : _GEN_189; // @[playground/src/noop/dcache.scala 137:45 139:27]
  wire  _GEN_193 = valid_1_3 & dirty_1_3 ? 1'h0 : _GEN_190; // @[playground/src/noop/dcache.scala 137:45 140:28]
  wire [3:0] _GEN_195 = valid_1_4 & dirty_1_4 ? 4'h4 : _GEN_192; // @[playground/src/noop/dcache.scala 137:45 139:27]
  wire  _GEN_196 = valid_1_4 & dirty_1_4 ? 1'h0 : _GEN_193; // @[playground/src/noop/dcache.scala 137:45 140:28]
  wire [3:0] _GEN_198 = valid_1_5 & dirty_1_5 ? 4'h5 : _GEN_195; // @[playground/src/noop/dcache.scala 137:45 139:27]
  wire  _GEN_199 = valid_1_5 & dirty_1_5 ? 1'h0 : _GEN_196; // @[playground/src/noop/dcache.scala 137:45 140:28]
  wire [3:0] _GEN_201 = valid_1_6 & dirty_1_6 ? 4'h6 : _GEN_198; // @[playground/src/noop/dcache.scala 137:45 139:27]
  wire  _GEN_202 = valid_1_6 & dirty_1_6 ? 1'h0 : _GEN_199; // @[playground/src/noop/dcache.scala 137:45 140:28]
  wire [3:0] _GEN_204 = valid_1_7 & dirty_1_7 ? 4'h7 : _GEN_201; // @[playground/src/noop/dcache.scala 137:45 139:27]
  wire  _GEN_205 = valid_1_7 & dirty_1_7 ? 1'h0 : _GEN_202; // @[playground/src/noop/dcache.scala 137:45 140:28]
  wire [3:0] _GEN_207 = valid_1_8 & dirty_1_8 ? 4'h8 : _GEN_204; // @[playground/src/noop/dcache.scala 137:45 139:27]
  wire  _GEN_208 = valid_1_8 & dirty_1_8 ? 1'h0 : _GEN_205; // @[playground/src/noop/dcache.scala 137:45 140:28]
  wire [3:0] _GEN_210 = valid_1_9 & dirty_1_9 ? 4'h9 : _GEN_207; // @[playground/src/noop/dcache.scala 137:45 139:27]
  wire  _GEN_211 = valid_1_9 & dirty_1_9 ? 1'h0 : _GEN_208; // @[playground/src/noop/dcache.scala 137:45 140:28]
  wire [3:0] _GEN_213 = valid_1_10 & dirty_1_10 ? 4'ha : _GEN_210; // @[playground/src/noop/dcache.scala 137:45 139:27]
  wire  _GEN_214 = valid_1_10 & dirty_1_10 ? 1'h0 : _GEN_211; // @[playground/src/noop/dcache.scala 137:45 140:28]
  wire [3:0] _GEN_216 = valid_1_11 & dirty_1_11 ? 4'hb : _GEN_213; // @[playground/src/noop/dcache.scala 137:45 139:27]
  wire  _GEN_217 = valid_1_11 & dirty_1_11 ? 1'h0 : _GEN_214; // @[playground/src/noop/dcache.scala 137:45 140:28]
  wire [3:0] _GEN_219 = valid_1_12 & dirty_1_12 ? 4'hc : _GEN_216; // @[playground/src/noop/dcache.scala 137:45 139:27]
  wire  _GEN_220 = valid_1_12 & dirty_1_12 ? 1'h0 : _GEN_217; // @[playground/src/noop/dcache.scala 137:45 140:28]
  wire [3:0] _GEN_222 = valid_1_13 & dirty_1_13 ? 4'hd : _GEN_219; // @[playground/src/noop/dcache.scala 137:45 139:27]
  wire  _GEN_223 = valid_1_13 & dirty_1_13 ? 1'h0 : _GEN_220; // @[playground/src/noop/dcache.scala 137:45 140:28]
  wire  _GEN_224 = valid_1_14 & dirty_1_14 | (valid_1_13 & dirty_1_13 | (valid_1_12 & dirty_1_12 | (valid_1_11 &
    dirty_1_11 | (valid_1_10 & dirty_1_10 | (valid_1_9 & dirty_1_9 | (valid_1_8 & dirty_1_8 | (valid_1_7 & dirty_1_7 | (
    valid_1_6 & dirty_1_6 | (valid_1_5 & dirty_1_5 | (valid_1_4 & dirty_1_4 | (valid_1_3 & dirty_1_3 | (valid_1_2 &
    dirty_1_2 | (valid_1_1 & dirty_1_1 | valid_1_0 & dirty_1_0))))))))))))); // @[playground/src/noop/dcache.scala 137:45 138:27]
  wire [3:0] _GEN_225 = valid_1_14 & dirty_1_14 ? 4'he : _GEN_222; // @[playground/src/noop/dcache.scala 137:45 139:27]
  wire  _GEN_226 = valid_1_14 & dirty_1_14 ? 1'h0 : _GEN_223; // @[playground/src/noop/dcache.scala 137:45 140:28]
  wire  _GEN_227 = valid_1_15 & dirty_1_15 | _GEN_224; // @[playground/src/noop/dcache.scala 137:45 138:27]
  wire [3:0] _GEN_228 = valid_1_15 & dirty_1_15 ? 4'hf : _GEN_225; // @[playground/src/noop/dcache.scala 137:45 139:27]
  wire  _GEN_229 = valid_1_15 & dirty_1_15 ? 1'h0 : _GEN_226; // @[playground/src/noop/dcache.scala 137:45 140:28]
  wire [1:0] _GEN_230 = valid_2_0 & dirty_2_0 ? 2'h2 : {{1'd0}, _GEN_227}; // @[playground/src/noop/dcache.scala 137:45 138:27]
  wire [3:0] _GEN_231 = valid_2_0 & dirty_2_0 ? 4'h0 : _GEN_228; // @[playground/src/noop/dcache.scala 137:45 139:27]
  wire  _GEN_232 = valid_2_0 & dirty_2_0 ? 1'h0 : _GEN_229; // @[playground/src/noop/dcache.scala 137:45 140:28]
  wire [1:0] _GEN_233 = valid_2_1 & dirty_2_1 ? 2'h2 : _GEN_230; // @[playground/src/noop/dcache.scala 137:45 138:27]
  wire [3:0] _GEN_234 = valid_2_1 & dirty_2_1 ? 4'h1 : _GEN_231; // @[playground/src/noop/dcache.scala 137:45 139:27]
  wire  _GEN_235 = valid_2_1 & dirty_2_1 ? 1'h0 : _GEN_232; // @[playground/src/noop/dcache.scala 137:45 140:28]
  wire [1:0] _GEN_236 = valid_2_2 & dirty_2_2 ? 2'h2 : _GEN_233; // @[playground/src/noop/dcache.scala 137:45 138:27]
  wire [3:0] _GEN_237 = valid_2_2 & dirty_2_2 ? 4'h2 : _GEN_234; // @[playground/src/noop/dcache.scala 137:45 139:27]
  wire  _GEN_238 = valid_2_2 & dirty_2_2 ? 1'h0 : _GEN_235; // @[playground/src/noop/dcache.scala 137:45 140:28]
  wire [1:0] _GEN_239 = valid_2_3 & dirty_2_3 ? 2'h2 : _GEN_236; // @[playground/src/noop/dcache.scala 137:45 138:27]
  wire [3:0] _GEN_240 = valid_2_3 & dirty_2_3 ? 4'h3 : _GEN_237; // @[playground/src/noop/dcache.scala 137:45 139:27]
  wire  _GEN_241 = valid_2_3 & dirty_2_3 ? 1'h0 : _GEN_238; // @[playground/src/noop/dcache.scala 137:45 140:28]
  wire [1:0] _GEN_242 = valid_2_4 & dirty_2_4 ? 2'h2 : _GEN_239; // @[playground/src/noop/dcache.scala 137:45 138:27]
  wire [3:0] _GEN_243 = valid_2_4 & dirty_2_4 ? 4'h4 : _GEN_240; // @[playground/src/noop/dcache.scala 137:45 139:27]
  wire  _GEN_244 = valid_2_4 & dirty_2_4 ? 1'h0 : _GEN_241; // @[playground/src/noop/dcache.scala 137:45 140:28]
  wire [1:0] _GEN_245 = valid_2_5 & dirty_2_5 ? 2'h2 : _GEN_242; // @[playground/src/noop/dcache.scala 137:45 138:27]
  wire [3:0] _GEN_246 = valid_2_5 & dirty_2_5 ? 4'h5 : _GEN_243; // @[playground/src/noop/dcache.scala 137:45 139:27]
  wire  _GEN_247 = valid_2_5 & dirty_2_5 ? 1'h0 : _GEN_244; // @[playground/src/noop/dcache.scala 137:45 140:28]
  wire [1:0] _GEN_248 = valid_2_6 & dirty_2_6 ? 2'h2 : _GEN_245; // @[playground/src/noop/dcache.scala 137:45 138:27]
  wire [3:0] _GEN_249 = valid_2_6 & dirty_2_6 ? 4'h6 : _GEN_246; // @[playground/src/noop/dcache.scala 137:45 139:27]
  wire  _GEN_250 = valid_2_6 & dirty_2_6 ? 1'h0 : _GEN_247; // @[playground/src/noop/dcache.scala 137:45 140:28]
  wire [1:0] _GEN_251 = valid_2_7 & dirty_2_7 ? 2'h2 : _GEN_248; // @[playground/src/noop/dcache.scala 137:45 138:27]
  wire [3:0] _GEN_252 = valid_2_7 & dirty_2_7 ? 4'h7 : _GEN_249; // @[playground/src/noop/dcache.scala 137:45 139:27]
  wire  _GEN_253 = valid_2_7 & dirty_2_7 ? 1'h0 : _GEN_250; // @[playground/src/noop/dcache.scala 137:45 140:28]
  wire [1:0] _GEN_254 = valid_2_8 & dirty_2_8 ? 2'h2 : _GEN_251; // @[playground/src/noop/dcache.scala 137:45 138:27]
  wire [3:0] _GEN_255 = valid_2_8 & dirty_2_8 ? 4'h8 : _GEN_252; // @[playground/src/noop/dcache.scala 137:45 139:27]
  wire  _GEN_256 = valid_2_8 & dirty_2_8 ? 1'h0 : _GEN_253; // @[playground/src/noop/dcache.scala 137:45 140:28]
  wire [1:0] _GEN_257 = valid_2_9 & dirty_2_9 ? 2'h2 : _GEN_254; // @[playground/src/noop/dcache.scala 137:45 138:27]
  wire [3:0] _GEN_258 = valid_2_9 & dirty_2_9 ? 4'h9 : _GEN_255; // @[playground/src/noop/dcache.scala 137:45 139:27]
  wire  _GEN_259 = valid_2_9 & dirty_2_9 ? 1'h0 : _GEN_256; // @[playground/src/noop/dcache.scala 137:45 140:28]
  wire [1:0] _GEN_260 = valid_2_10 & dirty_2_10 ? 2'h2 : _GEN_257; // @[playground/src/noop/dcache.scala 137:45 138:27]
  wire [3:0] _GEN_261 = valid_2_10 & dirty_2_10 ? 4'ha : _GEN_258; // @[playground/src/noop/dcache.scala 137:45 139:27]
  wire  _GEN_262 = valid_2_10 & dirty_2_10 ? 1'h0 : _GEN_259; // @[playground/src/noop/dcache.scala 137:45 140:28]
  wire [1:0] _GEN_263 = valid_2_11 & dirty_2_11 ? 2'h2 : _GEN_260; // @[playground/src/noop/dcache.scala 137:45 138:27]
  wire [3:0] _GEN_264 = valid_2_11 & dirty_2_11 ? 4'hb : _GEN_261; // @[playground/src/noop/dcache.scala 137:45 139:27]
  wire  _GEN_265 = valid_2_11 & dirty_2_11 ? 1'h0 : _GEN_262; // @[playground/src/noop/dcache.scala 137:45 140:28]
  wire [1:0] _GEN_266 = valid_2_12 & dirty_2_12 ? 2'h2 : _GEN_263; // @[playground/src/noop/dcache.scala 137:45 138:27]
  wire [3:0] _GEN_267 = valid_2_12 & dirty_2_12 ? 4'hc : _GEN_264; // @[playground/src/noop/dcache.scala 137:45 139:27]
  wire  _GEN_268 = valid_2_12 & dirty_2_12 ? 1'h0 : _GEN_265; // @[playground/src/noop/dcache.scala 137:45 140:28]
  wire [1:0] _GEN_269 = valid_2_13 & dirty_2_13 ? 2'h2 : _GEN_266; // @[playground/src/noop/dcache.scala 137:45 138:27]
  wire [3:0] _GEN_270 = valid_2_13 & dirty_2_13 ? 4'hd : _GEN_267; // @[playground/src/noop/dcache.scala 137:45 139:27]
  wire  _GEN_271 = valid_2_13 & dirty_2_13 ? 1'h0 : _GEN_268; // @[playground/src/noop/dcache.scala 137:45 140:28]
  wire [1:0] _GEN_272 = valid_2_14 & dirty_2_14 ? 2'h2 : _GEN_269; // @[playground/src/noop/dcache.scala 137:45 138:27]
  wire [3:0] _GEN_273 = valid_2_14 & dirty_2_14 ? 4'he : _GEN_270; // @[playground/src/noop/dcache.scala 137:45 139:27]
  wire  _GEN_274 = valid_2_14 & dirty_2_14 ? 1'h0 : _GEN_271; // @[playground/src/noop/dcache.scala 137:45 140:28]
  wire [1:0] _GEN_275 = valid_2_15 & dirty_2_15 ? 2'h2 : _GEN_272; // @[playground/src/noop/dcache.scala 137:45 138:27]
  wire [3:0] _GEN_276 = valid_2_15 & dirty_2_15 ? 4'hf : _GEN_273; // @[playground/src/noop/dcache.scala 137:45 139:27]
  wire  _GEN_277 = valid_2_15 & dirty_2_15 ? 1'h0 : _GEN_274; // @[playground/src/noop/dcache.scala 137:45 140:28]
  wire [1:0] _GEN_278 = valid_3_0 & dirty_3_0 ? 2'h3 : _GEN_275; // @[playground/src/noop/dcache.scala 137:45 138:27]
  wire [3:0] _GEN_279 = valid_3_0 & dirty_3_0 ? 4'h0 : _GEN_276; // @[playground/src/noop/dcache.scala 137:45 139:27]
  wire  _GEN_280 = valid_3_0 & dirty_3_0 ? 1'h0 : _GEN_277; // @[playground/src/noop/dcache.scala 137:45 140:28]
  wire [1:0] _GEN_281 = valid_3_1 & dirty_3_1 ? 2'h3 : _GEN_278; // @[playground/src/noop/dcache.scala 137:45 138:27]
  wire [3:0] _GEN_282 = valid_3_1 & dirty_3_1 ? 4'h1 : _GEN_279; // @[playground/src/noop/dcache.scala 137:45 139:27]
  wire  _GEN_283 = valid_3_1 & dirty_3_1 ? 1'h0 : _GEN_280; // @[playground/src/noop/dcache.scala 137:45 140:28]
  wire [1:0] _GEN_284 = valid_3_2 & dirty_3_2 ? 2'h3 : _GEN_281; // @[playground/src/noop/dcache.scala 137:45 138:27]
  wire [3:0] _GEN_285 = valid_3_2 & dirty_3_2 ? 4'h2 : _GEN_282; // @[playground/src/noop/dcache.scala 137:45 139:27]
  wire  _GEN_286 = valid_3_2 & dirty_3_2 ? 1'h0 : _GEN_283; // @[playground/src/noop/dcache.scala 137:45 140:28]
  wire [1:0] _GEN_287 = valid_3_3 & dirty_3_3 ? 2'h3 : _GEN_284; // @[playground/src/noop/dcache.scala 137:45 138:27]
  wire [3:0] _GEN_288 = valid_3_3 & dirty_3_3 ? 4'h3 : _GEN_285; // @[playground/src/noop/dcache.scala 137:45 139:27]
  wire  _GEN_289 = valid_3_3 & dirty_3_3 ? 1'h0 : _GEN_286; // @[playground/src/noop/dcache.scala 137:45 140:28]
  wire [1:0] _GEN_290 = valid_3_4 & dirty_3_4 ? 2'h3 : _GEN_287; // @[playground/src/noop/dcache.scala 137:45 138:27]
  wire [3:0] _GEN_291 = valid_3_4 & dirty_3_4 ? 4'h4 : _GEN_288; // @[playground/src/noop/dcache.scala 137:45 139:27]
  wire  _GEN_292 = valid_3_4 & dirty_3_4 ? 1'h0 : _GEN_289; // @[playground/src/noop/dcache.scala 137:45 140:28]
  wire [1:0] _GEN_293 = valid_3_5 & dirty_3_5 ? 2'h3 : _GEN_290; // @[playground/src/noop/dcache.scala 137:45 138:27]
  wire [3:0] _GEN_294 = valid_3_5 & dirty_3_5 ? 4'h5 : _GEN_291; // @[playground/src/noop/dcache.scala 137:45 139:27]
  wire  _GEN_295 = valid_3_5 & dirty_3_5 ? 1'h0 : _GEN_292; // @[playground/src/noop/dcache.scala 137:45 140:28]
  wire [1:0] _GEN_296 = valid_3_6 & dirty_3_6 ? 2'h3 : _GEN_293; // @[playground/src/noop/dcache.scala 137:45 138:27]
  wire [3:0] _GEN_297 = valid_3_6 & dirty_3_6 ? 4'h6 : _GEN_294; // @[playground/src/noop/dcache.scala 137:45 139:27]
  wire  _GEN_298 = valid_3_6 & dirty_3_6 ? 1'h0 : _GEN_295; // @[playground/src/noop/dcache.scala 137:45 140:28]
  wire [1:0] _GEN_299 = valid_3_7 & dirty_3_7 ? 2'h3 : _GEN_296; // @[playground/src/noop/dcache.scala 137:45 138:27]
  wire [3:0] _GEN_300 = valid_3_7 & dirty_3_7 ? 4'h7 : _GEN_297; // @[playground/src/noop/dcache.scala 137:45 139:27]
  wire  _GEN_301 = valid_3_7 & dirty_3_7 ? 1'h0 : _GEN_298; // @[playground/src/noop/dcache.scala 137:45 140:28]
  wire [1:0] _GEN_302 = valid_3_8 & dirty_3_8 ? 2'h3 : _GEN_299; // @[playground/src/noop/dcache.scala 137:45 138:27]
  wire [3:0] _GEN_303 = valid_3_8 & dirty_3_8 ? 4'h8 : _GEN_300; // @[playground/src/noop/dcache.scala 137:45 139:27]
  wire  _GEN_304 = valid_3_8 & dirty_3_8 ? 1'h0 : _GEN_301; // @[playground/src/noop/dcache.scala 137:45 140:28]
  wire [1:0] _GEN_305 = valid_3_9 & dirty_3_9 ? 2'h3 : _GEN_302; // @[playground/src/noop/dcache.scala 137:45 138:27]
  wire [3:0] _GEN_306 = valid_3_9 & dirty_3_9 ? 4'h9 : _GEN_303; // @[playground/src/noop/dcache.scala 137:45 139:27]
  wire  _GEN_307 = valid_3_9 & dirty_3_9 ? 1'h0 : _GEN_304; // @[playground/src/noop/dcache.scala 137:45 140:28]
  wire [1:0] _GEN_308 = valid_3_10 & dirty_3_10 ? 2'h3 : _GEN_305; // @[playground/src/noop/dcache.scala 137:45 138:27]
  wire [3:0] _GEN_309 = valid_3_10 & dirty_3_10 ? 4'ha : _GEN_306; // @[playground/src/noop/dcache.scala 137:45 139:27]
  wire  _GEN_310 = valid_3_10 & dirty_3_10 ? 1'h0 : _GEN_307; // @[playground/src/noop/dcache.scala 137:45 140:28]
  wire [1:0] _GEN_311 = valid_3_11 & dirty_3_11 ? 2'h3 : _GEN_308; // @[playground/src/noop/dcache.scala 137:45 138:27]
  wire [3:0] _GEN_312 = valid_3_11 & dirty_3_11 ? 4'hb : _GEN_309; // @[playground/src/noop/dcache.scala 137:45 139:27]
  wire  _GEN_313 = valid_3_11 & dirty_3_11 ? 1'h0 : _GEN_310; // @[playground/src/noop/dcache.scala 137:45 140:28]
  wire [1:0] _GEN_314 = valid_3_12 & dirty_3_12 ? 2'h3 : _GEN_311; // @[playground/src/noop/dcache.scala 137:45 138:27]
  wire [3:0] _GEN_315 = valid_3_12 & dirty_3_12 ? 4'hc : _GEN_312; // @[playground/src/noop/dcache.scala 137:45 139:27]
  wire  _GEN_316 = valid_3_12 & dirty_3_12 ? 1'h0 : _GEN_313; // @[playground/src/noop/dcache.scala 137:45 140:28]
  wire [1:0] _GEN_317 = valid_3_13 & dirty_3_13 ? 2'h3 : _GEN_314; // @[playground/src/noop/dcache.scala 137:45 138:27]
  wire [3:0] _GEN_318 = valid_3_13 & dirty_3_13 ? 4'hd : _GEN_315; // @[playground/src/noop/dcache.scala 137:45 139:27]
  wire  _GEN_319 = valid_3_13 & dirty_3_13 ? 1'h0 : _GEN_316; // @[playground/src/noop/dcache.scala 137:45 140:28]
  wire [1:0] _GEN_320 = valid_3_14 & dirty_3_14 ? 2'h3 : _GEN_317; // @[playground/src/noop/dcache.scala 137:45 138:27]
  wire [3:0] _GEN_321 = valid_3_14 & dirty_3_14 ? 4'he : _GEN_318; // @[playground/src/noop/dcache.scala 137:45 139:27]
  wire  _GEN_322 = valid_3_14 & dirty_3_14 ? 1'h0 : _GEN_319; // @[playground/src/noop/dcache.scala 137:45 140:28]
  wire [1:0] flush_way = valid_3_15 & dirty_3_15 ? 2'h3 : _GEN_320; // @[playground/src/noop/dcache.scala 137:45 138:27]
  wire [3:0] flush_idx = valid_3_15 & dirty_3_15 ? 4'hf : _GEN_321; // @[playground/src/noop/dcache.scala 137:45 139:27]
  wire  flush_done = valid_3_15 & dirty_3_15 ? 1'h0 : _GEN_322; // @[playground/src/noop/dcache.scala 137:45 140:28]
  wire [5:0] cur_ram_addr = cur_addr[9:4]; // @[playground/src/noop/dcache.scala 145:35]
  wire [5:0] _cur_axi_addr_T_1 = {flush_idx,offset[2:1]}; // @[playground/src/noop/dcache.scala 146:43]
  wire [5:0] _cur_axi_addr_T_4 = {blockIdx,offset[2:1]}; // @[playground/src/noop/dcache.scala 146:72]
  wire [5:0] cur_axi_addr = flush_r ? _cur_axi_addr_T_1 : _cur_axi_addr_T_4; // @[playground/src/noop/dcache.scala 146:30]
  wire [3:0] pre_blockIdx = addr_r[9:6]; // @[playground/src/noop/dcache.scala 149:33]
  wire [21:0] pre_tag = addr_r[31:10]; // @[playground/src/noop/dcache.scala 150:29]
  reg [2:0] state; // @[playground/src/noop/dcache.scala 152:24]
  wire [6:0] _rdata64_T_1 = {addr_r[3:0],3'h0}; // @[playground/src/noop/dcache.scala 153:48]
  wire [127:0] data_0_rdata = Ram_bw_io_rdata; // @[playground/src/noop/dcache.scala 91:{26,26}]
  wire [127:0] data_1_rdata = Ram_bw_1_io_rdata; // @[playground/src/noop/dcache.scala 91:{26,26}]
  wire [127:0] _GEN_327 = 2'h1 == matchWay_r ? data_1_rdata : data_0_rdata; // @[playground/src/noop/dcache.scala 153:{42,42}]
  wire [127:0] data_2_rdata = Ram_bw_2_io_rdata; // @[playground/src/noop/dcache.scala 91:{26,26}]
  wire [127:0] _GEN_328 = 2'h2 == matchWay_r ? data_2_rdata : _GEN_327; // @[playground/src/noop/dcache.scala 153:{42,42}]
  wire [127:0] data_3_rdata = Ram_bw_3_io_rdata; // @[playground/src/noop/dcache.scala 91:{26,26}]
  wire [127:0] _GEN_329 = 2'h3 == matchWay_r ? data_3_rdata : _GEN_328; // @[playground/src/noop/dcache.scala 153:{42,42}]
  wire [127:0] rdata64 = _GEN_329 >> _rdata64_T_1; // @[playground/src/noop/dcache.scala 153:42]
  wire [55:0] _io_dcRW_rdata_T_2 = rdata64[7] ? 56'hffffffffffffff : 56'h0; // @[playground/src/noop/common.scala 296:33]
  wire [63:0] _io_dcRW_rdata_T_4 = {_io_dcRW_rdata_T_2,rdata64[7:0]}; // @[playground/src/noop/common.scala 296:28]
  wire [47:0] _io_dcRW_rdata_T_8 = rdata64[15] ? 48'hffffffffffff : 48'h0; // @[playground/src/noop/common.scala 298:33]
  wire [63:0] _io_dcRW_rdata_T_10 = {_io_dcRW_rdata_T_8,rdata64[15:0]}; // @[playground/src/noop/common.scala 298:28]
  wire [31:0] _io_dcRW_rdata_T_14 = rdata64[31] ? 32'hffffffff : 32'h0; // @[playground/src/noop/common.scala 300:33]
  wire [63:0] _io_dcRW_rdata_T_16 = {_io_dcRW_rdata_T_14,rdata64[31:0]}; // @[playground/src/noop/common.scala 300:28]
  wire [63:0] _io_dcRW_rdata_T_24 = 5'h4 == mode_r ? _io_dcRW_rdata_T_4 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 81:58]
  wire [63:0] _io_dcRW_rdata_T_26 = 5'h14 == mode_r ? {{56'd0}, rdata64[7:0]} : _io_dcRW_rdata_T_24; // @[src/main/scala/chisel3/util/Mux.scala 81:58]
  wire [63:0] _io_dcRW_rdata_T_28 = 5'h5 == mode_r ? _io_dcRW_rdata_T_10 : _io_dcRW_rdata_T_26; // @[src/main/scala/chisel3/util/Mux.scala 81:58]
  wire [63:0] _io_dcRW_rdata_T_30 = 5'h15 == mode_r ? {{48'd0}, rdata64[15:0]} : _io_dcRW_rdata_T_28; // @[src/main/scala/chisel3/util/Mux.scala 81:58]
  wire [63:0] _io_dcRW_rdata_T_32 = 5'h6 == mode_r ? _io_dcRW_rdata_T_16 : _io_dcRW_rdata_T_30; // @[src/main/scala/chisel3/util/Mux.scala 81:58]
  wire [63:0] _io_dcRW_rdata_T_34 = 5'h16 == mode_r ? {{32'd0}, rdata64[31:0]} : _io_dcRW_rdata_T_32; // @[src/main/scala/chisel3/util/Mux.scala 81:58]
  wire [127:0] _io_dcRW_rdata_T_36 = 5'h7 == mode_r ? rdata64 : {{64'd0}, _io_dcRW_rdata_T_34}; // @[src/main/scala/chisel3/util/Mux.scala 81:58]
  wire [127:0] _io_dcRW_rdata_T_38 = 5'he == mode_r ? {{64'd0}, _io_dcRW_rdata_T_16} : _io_dcRW_rdata_T_36; // @[src/main/scala/chisel3/util/Mux.scala 81:58]
  wire [127:0] _io_dcRW_rdata_T_40 = 5'hf == mode_r ? rdata64 : _io_dcRW_rdata_T_38; // @[src/main/scala/chisel3/util/Mux.scala 81:58]
  wire [1:0] cur_mode_sl = _GEN_130[3:2]; // @[playground/src/noop/dcache.scala 155:31]
  wire [63:0] _amo_rdata_ans_T_17 = 2'h2 == mode_r[1:0] ? _io_dcRW_rdata_T_16 : rdata64[63:0]; // @[src/main/scala/chisel3/util/Mux.scala 81:58]
  wire [63:0] _amo_rdata_ans_T_19 = 2'h1 == mode_r[1:0] ? _io_dcRW_rdata_T_10 : _amo_rdata_ans_T_17; // @[src/main/scala/chisel3/util/Mux.scala 81:58]
  wire [63:0] amo_rdata = 2'h0 == mode_r[1:0] ? _io_dcRW_rdata_T_4 : _amo_rdata_ans_T_19; // @[src/main/scala/chisel3/util/Mux.scala 81:58]
  wire [31:0] _amo_imm_ans_T_3 = wdata_r[31] ? 32'hffffffff : 32'h0; // @[playground/src/noop/common.scala 319:28]
  wire [63:0] _amo_imm_ans_T_5 = {_amo_imm_ans_T_3,wdata_r[31:0]}; // @[playground/src/noop/common.scala 319:23]
  wire [47:0] _amo_imm_ans_T_8 = wdata_r[15] ? 48'hffffffffffff : 48'h0; // @[playground/src/noop/common.scala 320:28]
  wire [63:0] _amo_imm_ans_T_10 = {_amo_imm_ans_T_8,wdata_r[15:0]}; // @[playground/src/noop/common.scala 320:23]
  wire [55:0] _amo_imm_ans_T_13 = wdata_r[7] ? 56'hffffffffffffff : 56'h0; // @[playground/src/noop/common.scala 321:28]
  wire [63:0] _amo_imm_ans_T_15 = {_amo_imm_ans_T_13,wdata_r[7:0]}; // @[playground/src/noop/common.scala 321:23]
  wire [63:0] _amo_imm_ans_T_17 = 2'h2 == mode_r[1:0] ? _amo_imm_ans_T_5 : wdata_r; // @[src/main/scala/chisel3/util/Mux.scala 81:58]
  wire [63:0] _amo_imm_ans_T_19 = 2'h1 == mode_r[1:0] ? _amo_imm_ans_T_10 : _amo_imm_ans_T_17; // @[src/main/scala/chisel3/util/Mux.scala 81:58]
  wire [63:0] amo_imm = 2'h0 == mode_r[1:0] ? _amo_imm_ans_T_15 : _amo_imm_ans_T_19; // @[src/main/scala/chisel3/util/Mux.scala 81:58]
  wire [63:0] _amo_alu_T_1 = amo_imm + amo_rdata; // @[playground/src/noop/dcache.scala 165:29]
  wire [63:0] _amo_alu_T_2 = amo_imm ^ amo_rdata; // @[playground/src/noop/dcache.scala 166:29]
  wire [63:0] _amo_alu_T_3 = amo_imm & amo_rdata; // @[playground/src/noop/dcache.scala 167:29]
  wire [63:0] _amo_alu_T_4 = amo_imm | amo_rdata; // @[playground/src/noop/dcache.scala 168:29]
  wire [63:0] _amo_alu_T_5 = 2'h0 == mode_r[1:0] ? _amo_imm_ans_T_15 : _amo_imm_ans_T_19; // @[playground/src/noop/dcache.scala 169:32]
  wire [63:0] _amo_alu_T_6 = 2'h0 == mode_r[1:0] ? _io_dcRW_rdata_T_4 : _amo_rdata_ans_T_19; // @[playground/src/noop/dcache.scala 169:51]
  wire  _amo_alu_T_7 = $signed(_amo_alu_T_5) > $signed(_amo_alu_T_6); // @[playground/src/noop/dcache.scala 169:39]
  wire [63:0] _amo_alu_T_8 = $signed(_amo_alu_T_5) > $signed(_amo_alu_T_6) ? amo_rdata : amo_imm; // @[playground/src/noop/dcache.scala 169:23]
  wire [63:0] _amo_alu_T_12 = _amo_alu_T_7 ? amo_imm : amo_rdata; // @[playground/src/noop/dcache.scala 170:23]
  wire  _amo_alu_T_13 = amo_imm > amo_rdata; // @[playground/src/noop/dcache.scala 171:32]
  wire [63:0] _amo_alu_T_14 = amo_imm > amo_rdata ? amo_rdata : amo_imm; // @[playground/src/noop/dcache.scala 171:23]
  wire [63:0] _amo_alu_T_16 = _amo_alu_T_13 ? amo_imm : amo_rdata; // @[playground/src/noop/dcache.scala 172:23]
  wire [63:0] _amo_alu_T_18 = 5'h1 == amo_r ? amo_imm : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 81:58]
  wire [63:0] _amo_alu_T_20 = 5'h0 == amo_r ? _amo_alu_T_1 : _amo_alu_T_18; // @[src/main/scala/chisel3/util/Mux.scala 81:58]
  wire [63:0] _amo_alu_T_22 = 5'h4 == amo_r ? _amo_alu_T_2 : _amo_alu_T_20; // @[src/main/scala/chisel3/util/Mux.scala 81:58]
  wire [63:0] _amo_alu_T_24 = 5'hc == amo_r ? _amo_alu_T_3 : _amo_alu_T_22; // @[src/main/scala/chisel3/util/Mux.scala 81:58]
  wire [63:0] _amo_alu_T_26 = 5'h8 == amo_r ? _amo_alu_T_4 : _amo_alu_T_24; // @[src/main/scala/chisel3/util/Mux.scala 81:58]
  wire [63:0] _amo_alu_T_28 = 5'h10 == amo_r ? _amo_alu_T_8 : _amo_alu_T_26; // @[src/main/scala/chisel3/util/Mux.scala 81:58]
  wire [63:0] _amo_alu_T_30 = 5'h14 == amo_r ? _amo_alu_T_12 : _amo_alu_T_28; // @[src/main/scala/chisel3/util/Mux.scala 81:58]
  wire [63:0] _amo_alu_T_32 = 5'h1c == amo_r ? _amo_alu_T_14 : _amo_alu_T_30; // @[src/main/scala/chisel3/util/Mux.scala 81:58]
  wire [63:0] amo_alu = 5'h1c == amo_r ? _amo_alu_T_16 : _amo_alu_T_32; // @[src/main/scala/chisel3/util/Mux.scala 81:58]
  wire [63:0] _amo_wdata_ans_T_2 = {32'h0,amo_alu[31:0]}; // @[playground/src/noop/common.scala 310:23]
  wire [63:0] _amo_wdata_ans_T_4 = {48'h0,amo_alu[15:0]}; // @[playground/src/noop/common.scala 311:23]
  wire [63:0] _amo_wdata_ans_T_6 = {56'h0,amo_alu[7:0]}; // @[playground/src/noop/common.scala 312:23]
  wire [63:0] _amo_wdata_ans_T_8 = 2'h2 == mode_r[1:0] ? _amo_wdata_ans_T_2 : amo_alu; // @[src/main/scala/chisel3/util/Mux.scala 81:58]
  wire [63:0] _amo_wdata_ans_T_10 = 2'h1 == mode_r[1:0] ? _amo_wdata_ans_T_4 : _amo_wdata_ans_T_8; // @[src/main/scala/chisel3/util/Mux.scala 81:58]
  wire [63:0] amo_wdata_ans = 2'h0 == mode_r[1:0] ? _amo_wdata_ans_T_6 : _amo_wdata_ans_T_10; // @[src/main/scala/chisel3/util/Mux.scala 81:58]
  wire [6:0] _amo_wdata_T_2 = {cur_addr[3:0],3'h0}; // @[playground/src/noop/dcache.scala 174:67]
  wire [190:0] _GEN_3560 = {{127'd0}, amo_wdata_ans}; // @[playground/src/noop/dcache.scala 174:60]
  wire [190:0] amo_wdata = _GEN_3560 << _amo_wdata_T_2; // @[playground/src/noop/dcache.scala 174:60]
  wire [190:0] _GEN_3561 = {{127'd0}, _GEN_131}; // @[playground/src/noop/dcache.scala 176:32]
  wire [190:0] inp_wdata = _GEN_3561 << _amo_wdata_T_2; // @[playground/src/noop/dcache.scala 176:32]
  wire [127:0] _inp_mask_T_2 = 2'h1 == _GEN_130[1:0] ? 128'hffff : 128'hff; // @[src/main/scala/chisel3/util/Mux.scala 81:58]
  wire [127:0] _inp_mask_T_4 = 2'h2 == _GEN_130[1:0] ? 128'hffffffff : _inp_mask_T_2; // @[src/main/scala/chisel3/util/Mux.scala 81:58]
  wire [127:0] _inp_mask_T_6 = 2'h3 == _GEN_130[1:0] ? 128'hffffffffffffffff : _inp_mask_T_4; // @[src/main/scala/chisel3/util/Mux.scala 81:58]
  wire [254:0] _GEN_3562 = {{127'd0}, _inp_mask_T_6}; // @[playground/src/noop/dcache.scala 182:24]
  wire [254:0] inp_mask = _GEN_3562 << _amo_wdata_T_2; // @[playground/src/noop/dcache.scala 182:24]
  wire  _data_addr_T = state == 3'h0; // @[playground/src/noop/dcache.scala 183:38]
  wire  _data_addr_T_1 = state == 3'h5; // @[playground/src/noop/dcache.scala 183:57]
  wire  _data_addr_T_2 = state == 3'h0 | state == 3'h5; // @[playground/src/noop/dcache.scala 183:48]
  wire [5:0] _data_addr_T_3 = state == 3'h0 | state == 3'h5 ? cur_ram_addr : cur_axi_addr; // @[playground/src/noop/dcache.scala 183:31]
  wire  _GEN_2524 = 2'h0 == _GEN_129; // @[playground/src/noop/dcache.scala 184:{25,25} playground/src/ram/ram.scala 41:17]
  wire  _GEN_2525 = 2'h1 == _GEN_129; // @[playground/src/noop/dcache.scala 184:{25,25} playground/src/ram/ram.scala 41:17]
  wire  _GEN_2526 = 2'h2 == _GEN_129; // @[playground/src/noop/dcache.scala 184:{25,25} playground/src/ram/ram.scala 41:17]
  wire  _GEN_2527 = 2'h3 == _GEN_129; // @[playground/src/noop/dcache.scala 184:{25,25} playground/src/ram/ram.scala 41:17]
  wire  _T_73 = cur_mode_sl == 2'h3; // @[playground/src/noop/dcache.scala 212:34]
  wire  _GEN_545 = cur_mode_sl == 2'h3 ? 1'h0 : _GEN_130[3]; // @[playground/src/noop/dcache.scala 189:13 212:42 217:25]
  wire  _GEN_617 = cacheHit & _GEN_545; // @[playground/src/noop/dcache.scala 189:13 211:33]
  wire  _GEN_624 = ~hs_in & _io_dcRW_ready_T ? 1'h0 : _GEN_617; // @[playground/src/noop/dcache.scala 189:13 209:42]
  wire  _GEN_631 = flush_r | io_flush ? 1'h0 : _GEN_624; // @[playground/src/noop/dcache.scala 189:13 207:38]
  reg  axiRdataEn; // @[playground/src/noop/dcache.scala 198:34]
  wire  _GEN_899 = axiRdataEn & io_dataAxi_rd_valid & offset[0]; // @[playground/src/noop/dcache.scala 189:13 243:52]
  wire  _GEN_1764 = 3'h4 == state ? 1'h0 : 3'h5 == state; // @[playground/src/noop/dcache.scala 189:13 205:18]
  wire  _GEN_1903 = 3'h3 == state ? 1'h0 : _GEN_1764; // @[playground/src/noop/dcache.scala 189:13 205:18]
  wire  _GEN_1910 = 3'h2 == state ? _GEN_899 : _GEN_1903; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_2117 = 3'h1 == state ? 1'h0 : _GEN_1910; // @[playground/src/noop/dcache.scala 189:13 205:18]
  wire  wen = 3'h0 == state ? _GEN_631 : _GEN_2117; // @[playground/src/noop/dcache.scala 205:18]
  wire [127:0] _data_wdata_T_2 = {io_dataAxi_rd_bits_data,rdatabuf}; // @[playground/src/noop/dcache.scala 187:64]
  wire [190:0] _data_wdata_T_3 = _data_addr_T ? inp_wdata : {{63'd0}, _data_wdata_T_2}; // @[playground/src/noop/dcache.scala 187:32]
  wire [190:0] _data_wdata_T_4 = _data_addr_T_1 ? amo_wdata : _data_wdata_T_3; // @[playground/src/noop/dcache.scala 186:31]
  wire [254:0] _GEN_546 = cur_mode_sl == 2'h3 ? 255'hffffffffffffffffffffffffffffffff : inp_mask; // @[playground/src/noop/dcache.scala 190:13 212:42 218:26]
  wire [254:0] _GEN_618 = cacheHit ? _GEN_546 : 255'hffffffffffffffffffffffffffffffff; // @[playground/src/noop/dcache.scala 190:13 211:33]
  wire [254:0] _GEN_625 = ~hs_in & _io_dcRW_ready_T ? 255'hffffffffffffffffffffffffffffffff : _GEN_618; // @[playground/src/noop/dcache.scala 190:13 209:42]
  wire [254:0] _GEN_632 = flush_r | io_flush ? 255'hffffffffffffffffffffffffffffffff : _GEN_625; // @[playground/src/noop/dcache.scala 190:13 207:38]
  wire [254:0] _GEN_1562 = 3'h5 == state ? inp_mask : 255'hffffffffffffffffffffffffffffffff; // @[playground/src/noop/dcache.scala 190:13 205:18 281:21]
  wire [254:0] _GEN_1765 = 3'h4 == state ? 255'hffffffffffffffffffffffffffffffff : _GEN_1562; // @[playground/src/noop/dcache.scala 190:13 205:18]
  wire [254:0] _GEN_1904 = 3'h3 == state ? 255'hffffffffffffffffffffffffffffffff : _GEN_1765; // @[playground/src/noop/dcache.scala 190:13 205:18]
  wire [254:0] _GEN_2108 = 3'h2 == state ? 255'hffffffffffffffffffffffffffffffff : _GEN_1904; // @[playground/src/noop/dcache.scala 190:13 205:18]
  wire [254:0] _GEN_2313 = 3'h1 == state ? 255'hffffffffffffffffffffffffffffffff : _GEN_2108; // @[playground/src/noop/dcache.scala 190:13 205:18]
  wire [254:0] _GEN_2322 = 3'h0 == state ? _GEN_632 : _GEN_2313; // @[playground/src/noop/dcache.scala 205:18]
  wire [127:0] mask = _GEN_2322[127:0]; // @[playground/src/noop/dcache.scala 159:23]
  wire  _GEN_2533 = 4'h0 == blockIdx; // @[playground/src/noop/dcache.scala 192:{34,34} 90:26]
  wire  _GEN_350 = _GEN_2524 & 4'h0 == blockIdx | dirty_0_0; // @[playground/src/noop/dcache.scala 192:{34,34} 90:26]
  wire  _GEN_2536 = 4'h1 == blockIdx; // @[playground/src/noop/dcache.scala 192:{34,34} 90:26]
  wire  _GEN_351 = _GEN_2524 & 4'h1 == blockIdx | dirty_0_1; // @[playground/src/noop/dcache.scala 192:{34,34} 90:26]
  wire  _GEN_2539 = 4'h2 == blockIdx; // @[playground/src/noop/dcache.scala 192:{34,34} 90:26]
  wire  _GEN_352 = _GEN_2524 & 4'h2 == blockIdx | dirty_0_2; // @[playground/src/noop/dcache.scala 192:{34,34} 90:26]
  wire  _GEN_2542 = 4'h3 == blockIdx; // @[playground/src/noop/dcache.scala 192:{34,34} 90:26]
  wire  _GEN_353 = _GEN_2524 & 4'h3 == blockIdx | dirty_0_3; // @[playground/src/noop/dcache.scala 192:{34,34} 90:26]
  wire  _GEN_2545 = 4'h4 == blockIdx; // @[playground/src/noop/dcache.scala 192:{34,34} 90:26]
  wire  _GEN_354 = _GEN_2524 & 4'h4 == blockIdx | dirty_0_4; // @[playground/src/noop/dcache.scala 192:{34,34} 90:26]
  wire  _GEN_2548 = 4'h5 == blockIdx; // @[playground/src/noop/dcache.scala 192:{34,34} 90:26]
  wire  _GEN_355 = _GEN_2524 & 4'h5 == blockIdx | dirty_0_5; // @[playground/src/noop/dcache.scala 192:{34,34} 90:26]
  wire  _GEN_2551 = 4'h6 == blockIdx; // @[playground/src/noop/dcache.scala 192:{34,34} 90:26]
  wire  _GEN_356 = _GEN_2524 & 4'h6 == blockIdx | dirty_0_6; // @[playground/src/noop/dcache.scala 192:{34,34} 90:26]
  wire  _GEN_2554 = 4'h7 == blockIdx; // @[playground/src/noop/dcache.scala 192:{34,34} 90:26]
  wire  _GEN_357 = _GEN_2524 & 4'h7 == blockIdx | dirty_0_7; // @[playground/src/noop/dcache.scala 192:{34,34} 90:26]
  wire  _GEN_2557 = 4'h8 == blockIdx; // @[playground/src/noop/dcache.scala 192:{34,34} 90:26]
  wire  _GEN_358 = _GEN_2524 & 4'h8 == blockIdx | dirty_0_8; // @[playground/src/noop/dcache.scala 192:{34,34} 90:26]
  wire  _GEN_2560 = 4'h9 == blockIdx; // @[playground/src/noop/dcache.scala 192:{34,34} 90:26]
  wire  _GEN_359 = _GEN_2524 & 4'h9 == blockIdx | dirty_0_9; // @[playground/src/noop/dcache.scala 192:{34,34} 90:26]
  wire  _GEN_2563 = 4'ha == blockIdx; // @[playground/src/noop/dcache.scala 192:{34,34} 90:26]
  wire  _GEN_360 = _GEN_2524 & 4'ha == blockIdx | dirty_0_10; // @[playground/src/noop/dcache.scala 192:{34,34} 90:26]
  wire  _GEN_2566 = 4'hb == blockIdx; // @[playground/src/noop/dcache.scala 192:{34,34} 90:26]
  wire  _GEN_361 = _GEN_2524 & 4'hb == blockIdx | dirty_0_11; // @[playground/src/noop/dcache.scala 192:{34,34} 90:26]
  wire  _GEN_2569 = 4'hc == blockIdx; // @[playground/src/noop/dcache.scala 192:{34,34} 90:26]
  wire  _GEN_362 = _GEN_2524 & 4'hc == blockIdx | dirty_0_12; // @[playground/src/noop/dcache.scala 192:{34,34} 90:26]
  wire  _GEN_2572 = 4'hd == blockIdx; // @[playground/src/noop/dcache.scala 192:{34,34} 90:26]
  wire  _GEN_363 = _GEN_2524 & 4'hd == blockIdx | dirty_0_13; // @[playground/src/noop/dcache.scala 192:{34,34} 90:26]
  wire  _GEN_2575 = 4'he == blockIdx; // @[playground/src/noop/dcache.scala 192:{34,34} 90:26]
  wire  _GEN_364 = _GEN_2524 & 4'he == blockIdx | dirty_0_14; // @[playground/src/noop/dcache.scala 192:{34,34} 90:26]
  wire  _GEN_2578 = 4'hf == blockIdx; // @[playground/src/noop/dcache.scala 192:{34,34} 90:26]
  wire  _GEN_365 = _GEN_2524 & 4'hf == blockIdx | dirty_0_15; // @[playground/src/noop/dcache.scala 192:{34,34} 90:26]
  wire  _GEN_366 = _GEN_2525 & 4'h0 == blockIdx | dirty_1_0; // @[playground/src/noop/dcache.scala 192:{34,34} 90:26]
  wire  _GEN_367 = _GEN_2525 & 4'h1 == blockIdx | dirty_1_1; // @[playground/src/noop/dcache.scala 192:{34,34} 90:26]
  wire  _GEN_368 = _GEN_2525 & 4'h2 == blockIdx | dirty_1_2; // @[playground/src/noop/dcache.scala 192:{34,34} 90:26]
  wire  _GEN_369 = _GEN_2525 & 4'h3 == blockIdx | dirty_1_3; // @[playground/src/noop/dcache.scala 192:{34,34} 90:26]
  wire  _GEN_370 = _GEN_2525 & 4'h4 == blockIdx | dirty_1_4; // @[playground/src/noop/dcache.scala 192:{34,34} 90:26]
  wire  _GEN_371 = _GEN_2525 & 4'h5 == blockIdx | dirty_1_5; // @[playground/src/noop/dcache.scala 192:{34,34} 90:26]
  wire  _GEN_372 = _GEN_2525 & 4'h6 == blockIdx | dirty_1_6; // @[playground/src/noop/dcache.scala 192:{34,34} 90:26]
  wire  _GEN_373 = _GEN_2525 & 4'h7 == blockIdx | dirty_1_7; // @[playground/src/noop/dcache.scala 192:{34,34} 90:26]
  wire  _GEN_374 = _GEN_2525 & 4'h8 == blockIdx | dirty_1_8; // @[playground/src/noop/dcache.scala 192:{34,34} 90:26]
  wire  _GEN_375 = _GEN_2525 & 4'h9 == blockIdx | dirty_1_9; // @[playground/src/noop/dcache.scala 192:{34,34} 90:26]
  wire  _GEN_376 = _GEN_2525 & 4'ha == blockIdx | dirty_1_10; // @[playground/src/noop/dcache.scala 192:{34,34} 90:26]
  wire  _GEN_377 = _GEN_2525 & 4'hb == blockIdx | dirty_1_11; // @[playground/src/noop/dcache.scala 192:{34,34} 90:26]
  wire  _GEN_378 = _GEN_2525 & 4'hc == blockIdx | dirty_1_12; // @[playground/src/noop/dcache.scala 192:{34,34} 90:26]
  wire  _GEN_379 = _GEN_2525 & 4'hd == blockIdx | dirty_1_13; // @[playground/src/noop/dcache.scala 192:{34,34} 90:26]
  wire  _GEN_380 = _GEN_2525 & 4'he == blockIdx | dirty_1_14; // @[playground/src/noop/dcache.scala 192:{34,34} 90:26]
  wire  _GEN_381 = _GEN_2525 & 4'hf == blockIdx | dirty_1_15; // @[playground/src/noop/dcache.scala 192:{34,34} 90:26]
  wire  _GEN_382 = _GEN_2526 & 4'h0 == blockIdx | dirty_2_0; // @[playground/src/noop/dcache.scala 192:{34,34} 90:26]
  wire  _GEN_383 = _GEN_2526 & 4'h1 == blockIdx | dirty_2_1; // @[playground/src/noop/dcache.scala 192:{34,34} 90:26]
  wire  _GEN_384 = _GEN_2526 & 4'h2 == blockIdx | dirty_2_2; // @[playground/src/noop/dcache.scala 192:{34,34} 90:26]
  wire  _GEN_385 = _GEN_2526 & 4'h3 == blockIdx | dirty_2_3; // @[playground/src/noop/dcache.scala 192:{34,34} 90:26]
  wire  _GEN_386 = _GEN_2526 & 4'h4 == blockIdx | dirty_2_4; // @[playground/src/noop/dcache.scala 192:{34,34} 90:26]
  wire  _GEN_387 = _GEN_2526 & 4'h5 == blockIdx | dirty_2_5; // @[playground/src/noop/dcache.scala 192:{34,34} 90:26]
  wire  _GEN_388 = _GEN_2526 & 4'h6 == blockIdx | dirty_2_6; // @[playground/src/noop/dcache.scala 192:{34,34} 90:26]
  wire  _GEN_389 = _GEN_2526 & 4'h7 == blockIdx | dirty_2_7; // @[playground/src/noop/dcache.scala 192:{34,34} 90:26]
  wire  _GEN_390 = _GEN_2526 & 4'h8 == blockIdx | dirty_2_8; // @[playground/src/noop/dcache.scala 192:{34,34} 90:26]
  wire  _GEN_391 = _GEN_2526 & 4'h9 == blockIdx | dirty_2_9; // @[playground/src/noop/dcache.scala 192:{34,34} 90:26]
  wire  _GEN_392 = _GEN_2526 & 4'ha == blockIdx | dirty_2_10; // @[playground/src/noop/dcache.scala 192:{34,34} 90:26]
  wire  _GEN_393 = _GEN_2526 & 4'hb == blockIdx | dirty_2_11; // @[playground/src/noop/dcache.scala 192:{34,34} 90:26]
  wire  _GEN_394 = _GEN_2526 & 4'hc == blockIdx | dirty_2_12; // @[playground/src/noop/dcache.scala 192:{34,34} 90:26]
  wire  _GEN_395 = _GEN_2526 & 4'hd == blockIdx | dirty_2_13; // @[playground/src/noop/dcache.scala 192:{34,34} 90:26]
  wire  _GEN_396 = _GEN_2526 & 4'he == blockIdx | dirty_2_14; // @[playground/src/noop/dcache.scala 192:{34,34} 90:26]
  wire  _GEN_397 = _GEN_2526 & 4'hf == blockIdx | dirty_2_15; // @[playground/src/noop/dcache.scala 192:{34,34} 90:26]
  wire  _GEN_398 = _GEN_2527 & 4'h0 == blockIdx | dirty_3_0; // @[playground/src/noop/dcache.scala 192:{34,34} 90:26]
  wire  _GEN_399 = _GEN_2527 & 4'h1 == blockIdx | dirty_3_1; // @[playground/src/noop/dcache.scala 192:{34,34} 90:26]
  wire  _GEN_400 = _GEN_2527 & 4'h2 == blockIdx | dirty_3_2; // @[playground/src/noop/dcache.scala 192:{34,34} 90:26]
  wire  _GEN_401 = _GEN_2527 & 4'h3 == blockIdx | dirty_3_3; // @[playground/src/noop/dcache.scala 192:{34,34} 90:26]
  wire  _GEN_402 = _GEN_2527 & 4'h4 == blockIdx | dirty_3_4; // @[playground/src/noop/dcache.scala 192:{34,34} 90:26]
  wire  _GEN_403 = _GEN_2527 & 4'h5 == blockIdx | dirty_3_5; // @[playground/src/noop/dcache.scala 192:{34,34} 90:26]
  wire  _GEN_404 = _GEN_2527 & 4'h6 == blockIdx | dirty_3_6; // @[playground/src/noop/dcache.scala 192:{34,34} 90:26]
  wire  _GEN_405 = _GEN_2527 & 4'h7 == blockIdx | dirty_3_7; // @[playground/src/noop/dcache.scala 192:{34,34} 90:26]
  wire  _GEN_406 = _GEN_2527 & 4'h8 == blockIdx | dirty_3_8; // @[playground/src/noop/dcache.scala 192:{34,34} 90:26]
  wire  _GEN_407 = _GEN_2527 & 4'h9 == blockIdx | dirty_3_9; // @[playground/src/noop/dcache.scala 192:{34,34} 90:26]
  wire  _GEN_408 = _GEN_2527 & 4'ha == blockIdx | dirty_3_10; // @[playground/src/noop/dcache.scala 192:{34,34} 90:26]
  wire  _GEN_409 = _GEN_2527 & 4'hb == blockIdx | dirty_3_11; // @[playground/src/noop/dcache.scala 192:{34,34} 90:26]
  wire  _GEN_410 = _GEN_2527 & 4'hc == blockIdx | dirty_3_12; // @[playground/src/noop/dcache.scala 192:{34,34} 90:26]
  wire  _GEN_411 = _GEN_2527 & 4'hd == blockIdx | dirty_3_13; // @[playground/src/noop/dcache.scala 192:{34,34} 90:26]
  wire  _GEN_412 = _GEN_2527 & 4'he == blockIdx | dirty_3_14; // @[playground/src/noop/dcache.scala 192:{34,34} 90:26]
  wire  _GEN_413 = _GEN_2527 & 4'hf == blockIdx | dirty_3_15; // @[playground/src/noop/dcache.scala 192:{34,34} 90:26]
  wire  _GEN_414 = wen & _data_addr_T_2 ? _GEN_350 : dirty_0_0; // @[playground/src/noop/dcache.scala 191:56 90:26]
  wire  _GEN_415 = wen & _data_addr_T_2 ? _GEN_351 : dirty_0_1; // @[playground/src/noop/dcache.scala 191:56 90:26]
  wire  _GEN_416 = wen & _data_addr_T_2 ? _GEN_352 : dirty_0_2; // @[playground/src/noop/dcache.scala 191:56 90:26]
  wire  _GEN_417 = wen & _data_addr_T_2 ? _GEN_353 : dirty_0_3; // @[playground/src/noop/dcache.scala 191:56 90:26]
  wire  _GEN_418 = wen & _data_addr_T_2 ? _GEN_354 : dirty_0_4; // @[playground/src/noop/dcache.scala 191:56 90:26]
  wire  _GEN_419 = wen & _data_addr_T_2 ? _GEN_355 : dirty_0_5; // @[playground/src/noop/dcache.scala 191:56 90:26]
  wire  _GEN_420 = wen & _data_addr_T_2 ? _GEN_356 : dirty_0_6; // @[playground/src/noop/dcache.scala 191:56 90:26]
  wire  _GEN_421 = wen & _data_addr_T_2 ? _GEN_357 : dirty_0_7; // @[playground/src/noop/dcache.scala 191:56 90:26]
  wire  _GEN_422 = wen & _data_addr_T_2 ? _GEN_358 : dirty_0_8; // @[playground/src/noop/dcache.scala 191:56 90:26]
  wire  _GEN_423 = wen & _data_addr_T_2 ? _GEN_359 : dirty_0_9; // @[playground/src/noop/dcache.scala 191:56 90:26]
  wire  _GEN_424 = wen & _data_addr_T_2 ? _GEN_360 : dirty_0_10; // @[playground/src/noop/dcache.scala 191:56 90:26]
  wire  _GEN_425 = wen & _data_addr_T_2 ? _GEN_361 : dirty_0_11; // @[playground/src/noop/dcache.scala 191:56 90:26]
  wire  _GEN_426 = wen & _data_addr_T_2 ? _GEN_362 : dirty_0_12; // @[playground/src/noop/dcache.scala 191:56 90:26]
  wire  _GEN_427 = wen & _data_addr_T_2 ? _GEN_363 : dirty_0_13; // @[playground/src/noop/dcache.scala 191:56 90:26]
  wire  _GEN_428 = wen & _data_addr_T_2 ? _GEN_364 : dirty_0_14; // @[playground/src/noop/dcache.scala 191:56 90:26]
  wire  _GEN_429 = wen & _data_addr_T_2 ? _GEN_365 : dirty_0_15; // @[playground/src/noop/dcache.scala 191:56 90:26]
  wire  _GEN_430 = wen & _data_addr_T_2 ? _GEN_366 : dirty_1_0; // @[playground/src/noop/dcache.scala 191:56 90:26]
  wire  _GEN_431 = wen & _data_addr_T_2 ? _GEN_367 : dirty_1_1; // @[playground/src/noop/dcache.scala 191:56 90:26]
  wire  _GEN_432 = wen & _data_addr_T_2 ? _GEN_368 : dirty_1_2; // @[playground/src/noop/dcache.scala 191:56 90:26]
  wire  _GEN_433 = wen & _data_addr_T_2 ? _GEN_369 : dirty_1_3; // @[playground/src/noop/dcache.scala 191:56 90:26]
  wire  _GEN_434 = wen & _data_addr_T_2 ? _GEN_370 : dirty_1_4; // @[playground/src/noop/dcache.scala 191:56 90:26]
  wire  _GEN_435 = wen & _data_addr_T_2 ? _GEN_371 : dirty_1_5; // @[playground/src/noop/dcache.scala 191:56 90:26]
  wire  _GEN_436 = wen & _data_addr_T_2 ? _GEN_372 : dirty_1_6; // @[playground/src/noop/dcache.scala 191:56 90:26]
  wire  _GEN_437 = wen & _data_addr_T_2 ? _GEN_373 : dirty_1_7; // @[playground/src/noop/dcache.scala 191:56 90:26]
  wire  _GEN_438 = wen & _data_addr_T_2 ? _GEN_374 : dirty_1_8; // @[playground/src/noop/dcache.scala 191:56 90:26]
  wire  _GEN_439 = wen & _data_addr_T_2 ? _GEN_375 : dirty_1_9; // @[playground/src/noop/dcache.scala 191:56 90:26]
  wire  _GEN_440 = wen & _data_addr_T_2 ? _GEN_376 : dirty_1_10; // @[playground/src/noop/dcache.scala 191:56 90:26]
  wire  _GEN_441 = wen & _data_addr_T_2 ? _GEN_377 : dirty_1_11; // @[playground/src/noop/dcache.scala 191:56 90:26]
  wire  _GEN_442 = wen & _data_addr_T_2 ? _GEN_378 : dirty_1_12; // @[playground/src/noop/dcache.scala 191:56 90:26]
  wire  _GEN_443 = wen & _data_addr_T_2 ? _GEN_379 : dirty_1_13; // @[playground/src/noop/dcache.scala 191:56 90:26]
  wire  _GEN_444 = wen & _data_addr_T_2 ? _GEN_380 : dirty_1_14; // @[playground/src/noop/dcache.scala 191:56 90:26]
  wire  _GEN_445 = wen & _data_addr_T_2 ? _GEN_381 : dirty_1_15; // @[playground/src/noop/dcache.scala 191:56 90:26]
  wire  _GEN_446 = wen & _data_addr_T_2 ? _GEN_382 : dirty_2_0; // @[playground/src/noop/dcache.scala 191:56 90:26]
  wire  _GEN_447 = wen & _data_addr_T_2 ? _GEN_383 : dirty_2_1; // @[playground/src/noop/dcache.scala 191:56 90:26]
  wire  _GEN_448 = wen & _data_addr_T_2 ? _GEN_384 : dirty_2_2; // @[playground/src/noop/dcache.scala 191:56 90:26]
  wire  _GEN_449 = wen & _data_addr_T_2 ? _GEN_385 : dirty_2_3; // @[playground/src/noop/dcache.scala 191:56 90:26]
  wire  _GEN_450 = wen & _data_addr_T_2 ? _GEN_386 : dirty_2_4; // @[playground/src/noop/dcache.scala 191:56 90:26]
  wire  _GEN_451 = wen & _data_addr_T_2 ? _GEN_387 : dirty_2_5; // @[playground/src/noop/dcache.scala 191:56 90:26]
  wire  _GEN_452 = wen & _data_addr_T_2 ? _GEN_388 : dirty_2_6; // @[playground/src/noop/dcache.scala 191:56 90:26]
  wire  _GEN_453 = wen & _data_addr_T_2 ? _GEN_389 : dirty_2_7; // @[playground/src/noop/dcache.scala 191:56 90:26]
  wire  _GEN_454 = wen & _data_addr_T_2 ? _GEN_390 : dirty_2_8; // @[playground/src/noop/dcache.scala 191:56 90:26]
  wire  _GEN_455 = wen & _data_addr_T_2 ? _GEN_391 : dirty_2_9; // @[playground/src/noop/dcache.scala 191:56 90:26]
  wire  _GEN_456 = wen & _data_addr_T_2 ? _GEN_392 : dirty_2_10; // @[playground/src/noop/dcache.scala 191:56 90:26]
  wire  _GEN_457 = wen & _data_addr_T_2 ? _GEN_393 : dirty_2_11; // @[playground/src/noop/dcache.scala 191:56 90:26]
  wire  _GEN_458 = wen & _data_addr_T_2 ? _GEN_394 : dirty_2_12; // @[playground/src/noop/dcache.scala 191:56 90:26]
  wire  _GEN_459 = wen & _data_addr_T_2 ? _GEN_395 : dirty_2_13; // @[playground/src/noop/dcache.scala 191:56 90:26]
  wire  _GEN_460 = wen & _data_addr_T_2 ? _GEN_396 : dirty_2_14; // @[playground/src/noop/dcache.scala 191:56 90:26]
  wire  _GEN_461 = wen & _data_addr_T_2 ? _GEN_397 : dirty_2_15; // @[playground/src/noop/dcache.scala 191:56 90:26]
  wire  _GEN_462 = wen & _data_addr_T_2 ? _GEN_398 : dirty_3_0; // @[playground/src/noop/dcache.scala 191:56 90:26]
  wire  _GEN_463 = wen & _data_addr_T_2 ? _GEN_399 : dirty_3_1; // @[playground/src/noop/dcache.scala 191:56 90:26]
  wire  _GEN_464 = wen & _data_addr_T_2 ? _GEN_400 : dirty_3_2; // @[playground/src/noop/dcache.scala 191:56 90:26]
  wire  _GEN_465 = wen & _data_addr_T_2 ? _GEN_401 : dirty_3_3; // @[playground/src/noop/dcache.scala 191:56 90:26]
  wire  _GEN_466 = wen & _data_addr_T_2 ? _GEN_402 : dirty_3_4; // @[playground/src/noop/dcache.scala 191:56 90:26]
  wire  _GEN_467 = wen & _data_addr_T_2 ? _GEN_403 : dirty_3_5; // @[playground/src/noop/dcache.scala 191:56 90:26]
  wire  _GEN_468 = wen & _data_addr_T_2 ? _GEN_404 : dirty_3_6; // @[playground/src/noop/dcache.scala 191:56 90:26]
  wire  _GEN_469 = wen & _data_addr_T_2 ? _GEN_405 : dirty_3_7; // @[playground/src/noop/dcache.scala 191:56 90:26]
  wire  _GEN_470 = wen & _data_addr_T_2 ? _GEN_406 : dirty_3_8; // @[playground/src/noop/dcache.scala 191:56 90:26]
  wire  _GEN_471 = wen & _data_addr_T_2 ? _GEN_407 : dirty_3_9; // @[playground/src/noop/dcache.scala 191:56 90:26]
  wire  _GEN_472 = wen & _data_addr_T_2 ? _GEN_408 : dirty_3_10; // @[playground/src/noop/dcache.scala 191:56 90:26]
  wire  _GEN_473 = wen & _data_addr_T_2 ? _GEN_409 : dirty_3_11; // @[playground/src/noop/dcache.scala 191:56 90:26]
  wire  _GEN_474 = wen & _data_addr_T_2 ? _GEN_410 : dirty_3_12; // @[playground/src/noop/dcache.scala 191:56 90:26]
  wire  _GEN_475 = wen & _data_addr_T_2 ? _GEN_411 : dirty_3_13; // @[playground/src/noop/dcache.scala 191:56 90:26]
  wire  _GEN_476 = wen & _data_addr_T_2 ? _GEN_412 : dirty_3_14; // @[playground/src/noop/dcache.scala 191:56 90:26]
  wire  _GEN_477 = wen & _data_addr_T_2 ? _GEN_413 : dirty_3_15; // @[playground/src/noop/dcache.scala 191:56 90:26]
  reg  axiRaddrEn; // @[playground/src/noop/dcache.scala 196:34]
  reg  axiWaddrEn; // @[playground/src/noop/dcache.scala 199:34]
  wire  _GEN_2724 = 2'h0 == matchWay_r; // @[playground/src/noop/dcache.scala 200:{30,30}]
  wire  _GEN_2725 = 4'h1 == blockIdx_r; // @[playground/src/noop/dcache.scala 200:{30,30}]
  wire [21:0] _GEN_479 = 2'h0 == matchWay_r & 4'h1 == blockIdx_r ? tag_0_1 : tag_0_0; // @[playground/src/noop/dcache.scala 200:{30,30}]
  wire  _GEN_2727 = 4'h2 == blockIdx_r; // @[playground/src/noop/dcache.scala 200:{30,30}]
  wire [21:0] _GEN_480 = 2'h0 == matchWay_r & 4'h2 == blockIdx_r ? tag_0_2 : _GEN_479; // @[playground/src/noop/dcache.scala 200:{30,30}]
  wire  _GEN_2729 = 4'h3 == blockIdx_r; // @[playground/src/noop/dcache.scala 200:{30,30}]
  wire [21:0] _GEN_481 = 2'h0 == matchWay_r & 4'h3 == blockIdx_r ? tag_0_3 : _GEN_480; // @[playground/src/noop/dcache.scala 200:{30,30}]
  wire  _GEN_2731 = 4'h4 == blockIdx_r; // @[playground/src/noop/dcache.scala 200:{30,30}]
  wire [21:0] _GEN_482 = 2'h0 == matchWay_r & 4'h4 == blockIdx_r ? tag_0_4 : _GEN_481; // @[playground/src/noop/dcache.scala 200:{30,30}]
  wire  _GEN_2733 = 4'h5 == blockIdx_r; // @[playground/src/noop/dcache.scala 200:{30,30}]
  wire [21:0] _GEN_483 = 2'h0 == matchWay_r & 4'h5 == blockIdx_r ? tag_0_5 : _GEN_482; // @[playground/src/noop/dcache.scala 200:{30,30}]
  wire  _GEN_2735 = 4'h6 == blockIdx_r; // @[playground/src/noop/dcache.scala 200:{30,30}]
  wire [21:0] _GEN_484 = 2'h0 == matchWay_r & 4'h6 == blockIdx_r ? tag_0_6 : _GEN_483; // @[playground/src/noop/dcache.scala 200:{30,30}]
  wire  _GEN_2737 = 4'h7 == blockIdx_r; // @[playground/src/noop/dcache.scala 200:{30,30}]
  wire [21:0] _GEN_485 = 2'h0 == matchWay_r & 4'h7 == blockIdx_r ? tag_0_7 : _GEN_484; // @[playground/src/noop/dcache.scala 200:{30,30}]
  wire  _GEN_2739 = 4'h8 == blockIdx_r; // @[playground/src/noop/dcache.scala 200:{30,30}]
  wire [21:0] _GEN_486 = 2'h0 == matchWay_r & 4'h8 == blockIdx_r ? tag_0_8 : _GEN_485; // @[playground/src/noop/dcache.scala 200:{30,30}]
  wire  _GEN_2741 = 4'h9 == blockIdx_r; // @[playground/src/noop/dcache.scala 200:{30,30}]
  wire [21:0] _GEN_487 = 2'h0 == matchWay_r & 4'h9 == blockIdx_r ? tag_0_9 : _GEN_486; // @[playground/src/noop/dcache.scala 200:{30,30}]
  wire  _GEN_2743 = 4'ha == blockIdx_r; // @[playground/src/noop/dcache.scala 200:{30,30}]
  wire [21:0] _GEN_488 = 2'h0 == matchWay_r & 4'ha == blockIdx_r ? tag_0_10 : _GEN_487; // @[playground/src/noop/dcache.scala 200:{30,30}]
  wire  _GEN_2745 = 4'hb == blockIdx_r; // @[playground/src/noop/dcache.scala 200:{30,30}]
  wire [21:0] _GEN_489 = 2'h0 == matchWay_r & 4'hb == blockIdx_r ? tag_0_11 : _GEN_488; // @[playground/src/noop/dcache.scala 200:{30,30}]
  wire  _GEN_2747 = 4'hc == blockIdx_r; // @[playground/src/noop/dcache.scala 200:{30,30}]
  wire [21:0] _GEN_490 = 2'h0 == matchWay_r & 4'hc == blockIdx_r ? tag_0_12 : _GEN_489; // @[playground/src/noop/dcache.scala 200:{30,30}]
  wire  _GEN_2749 = 4'hd == blockIdx_r; // @[playground/src/noop/dcache.scala 200:{30,30}]
  wire [21:0] _GEN_491 = 2'h0 == matchWay_r & 4'hd == blockIdx_r ? tag_0_13 : _GEN_490; // @[playground/src/noop/dcache.scala 200:{30,30}]
  wire  _GEN_2751 = 4'he == blockIdx_r; // @[playground/src/noop/dcache.scala 200:{30,30}]
  wire [21:0] _GEN_492 = 2'h0 == matchWay_r & 4'he == blockIdx_r ? tag_0_14 : _GEN_491; // @[playground/src/noop/dcache.scala 200:{30,30}]
  wire  _GEN_2753 = 4'hf == blockIdx_r; // @[playground/src/noop/dcache.scala 200:{30,30}]
  wire [21:0] _GEN_493 = 2'h0 == matchWay_r & 4'hf == blockIdx_r ? tag_0_15 : _GEN_492; // @[playground/src/noop/dcache.scala 200:{30,30}]
  wire  _GEN_2754 = 2'h1 == matchWay_r; // @[playground/src/noop/dcache.scala 200:{30,30}]
  wire  _GEN_2755 = 4'h0 == blockIdx_r; // @[playground/src/noop/dcache.scala 200:{30,30}]
  wire [21:0] _GEN_494 = 2'h1 == matchWay_r & 4'h0 == blockIdx_r ? tag_1_0 : _GEN_493; // @[playground/src/noop/dcache.scala 200:{30,30}]
  wire [21:0] _GEN_495 = 2'h1 == matchWay_r & 4'h1 == blockIdx_r ? tag_1_1 : _GEN_494; // @[playground/src/noop/dcache.scala 200:{30,30}]
  wire [21:0] _GEN_496 = 2'h1 == matchWay_r & 4'h2 == blockIdx_r ? tag_1_2 : _GEN_495; // @[playground/src/noop/dcache.scala 200:{30,30}]
  wire [21:0] _GEN_497 = 2'h1 == matchWay_r & 4'h3 == blockIdx_r ? tag_1_3 : _GEN_496; // @[playground/src/noop/dcache.scala 200:{30,30}]
  wire [21:0] _GEN_498 = 2'h1 == matchWay_r & 4'h4 == blockIdx_r ? tag_1_4 : _GEN_497; // @[playground/src/noop/dcache.scala 200:{30,30}]
  wire [21:0] _GEN_499 = 2'h1 == matchWay_r & 4'h5 == blockIdx_r ? tag_1_5 : _GEN_498; // @[playground/src/noop/dcache.scala 200:{30,30}]
  wire [21:0] _GEN_500 = 2'h1 == matchWay_r & 4'h6 == blockIdx_r ? tag_1_6 : _GEN_499; // @[playground/src/noop/dcache.scala 200:{30,30}]
  wire [21:0] _GEN_501 = 2'h1 == matchWay_r & 4'h7 == blockIdx_r ? tag_1_7 : _GEN_500; // @[playground/src/noop/dcache.scala 200:{30,30}]
  wire [21:0] _GEN_502 = 2'h1 == matchWay_r & 4'h8 == blockIdx_r ? tag_1_8 : _GEN_501; // @[playground/src/noop/dcache.scala 200:{30,30}]
  wire [21:0] _GEN_503 = 2'h1 == matchWay_r & 4'h9 == blockIdx_r ? tag_1_9 : _GEN_502; // @[playground/src/noop/dcache.scala 200:{30,30}]
  wire [21:0] _GEN_504 = 2'h1 == matchWay_r & 4'ha == blockIdx_r ? tag_1_10 : _GEN_503; // @[playground/src/noop/dcache.scala 200:{30,30}]
  wire [21:0] _GEN_505 = 2'h1 == matchWay_r & 4'hb == blockIdx_r ? tag_1_11 : _GEN_504; // @[playground/src/noop/dcache.scala 200:{30,30}]
  wire [21:0] _GEN_506 = 2'h1 == matchWay_r & 4'hc == blockIdx_r ? tag_1_12 : _GEN_505; // @[playground/src/noop/dcache.scala 200:{30,30}]
  wire [21:0] _GEN_507 = 2'h1 == matchWay_r & 4'hd == blockIdx_r ? tag_1_13 : _GEN_506; // @[playground/src/noop/dcache.scala 200:{30,30}]
  wire [21:0] _GEN_508 = 2'h1 == matchWay_r & 4'he == blockIdx_r ? tag_1_14 : _GEN_507; // @[playground/src/noop/dcache.scala 200:{30,30}]
  wire [21:0] _GEN_509 = 2'h1 == matchWay_r & 4'hf == blockIdx_r ? tag_1_15 : _GEN_508; // @[playground/src/noop/dcache.scala 200:{30,30}]
  wire  _GEN_2786 = 2'h2 == matchWay_r; // @[playground/src/noop/dcache.scala 200:{30,30}]
  wire [21:0] _GEN_510 = 2'h2 == matchWay_r & 4'h0 == blockIdx_r ? tag_2_0 : _GEN_509; // @[playground/src/noop/dcache.scala 200:{30,30}]
  wire [21:0] _GEN_511 = 2'h2 == matchWay_r & 4'h1 == blockIdx_r ? tag_2_1 : _GEN_510; // @[playground/src/noop/dcache.scala 200:{30,30}]
  wire [21:0] _GEN_512 = 2'h2 == matchWay_r & 4'h2 == blockIdx_r ? tag_2_2 : _GEN_511; // @[playground/src/noop/dcache.scala 200:{30,30}]
  wire [21:0] _GEN_513 = 2'h2 == matchWay_r & 4'h3 == blockIdx_r ? tag_2_3 : _GEN_512; // @[playground/src/noop/dcache.scala 200:{30,30}]
  wire [21:0] _GEN_514 = 2'h2 == matchWay_r & 4'h4 == blockIdx_r ? tag_2_4 : _GEN_513; // @[playground/src/noop/dcache.scala 200:{30,30}]
  wire [21:0] _GEN_515 = 2'h2 == matchWay_r & 4'h5 == blockIdx_r ? tag_2_5 : _GEN_514; // @[playground/src/noop/dcache.scala 200:{30,30}]
  wire [21:0] _GEN_516 = 2'h2 == matchWay_r & 4'h6 == blockIdx_r ? tag_2_6 : _GEN_515; // @[playground/src/noop/dcache.scala 200:{30,30}]
  wire [21:0] _GEN_517 = 2'h2 == matchWay_r & 4'h7 == blockIdx_r ? tag_2_7 : _GEN_516; // @[playground/src/noop/dcache.scala 200:{30,30}]
  wire [21:0] _GEN_518 = 2'h2 == matchWay_r & 4'h8 == blockIdx_r ? tag_2_8 : _GEN_517; // @[playground/src/noop/dcache.scala 200:{30,30}]
  wire [21:0] _GEN_519 = 2'h2 == matchWay_r & 4'h9 == blockIdx_r ? tag_2_9 : _GEN_518; // @[playground/src/noop/dcache.scala 200:{30,30}]
  wire [21:0] _GEN_520 = 2'h2 == matchWay_r & 4'ha == blockIdx_r ? tag_2_10 : _GEN_519; // @[playground/src/noop/dcache.scala 200:{30,30}]
  wire [21:0] _GEN_521 = 2'h2 == matchWay_r & 4'hb == blockIdx_r ? tag_2_11 : _GEN_520; // @[playground/src/noop/dcache.scala 200:{30,30}]
  wire [21:0] _GEN_522 = 2'h2 == matchWay_r & 4'hc == blockIdx_r ? tag_2_12 : _GEN_521; // @[playground/src/noop/dcache.scala 200:{30,30}]
  wire [21:0] _GEN_523 = 2'h2 == matchWay_r & 4'hd == blockIdx_r ? tag_2_13 : _GEN_522; // @[playground/src/noop/dcache.scala 200:{30,30}]
  wire [21:0] _GEN_524 = 2'h2 == matchWay_r & 4'he == blockIdx_r ? tag_2_14 : _GEN_523; // @[playground/src/noop/dcache.scala 200:{30,30}]
  wire [21:0] _GEN_525 = 2'h2 == matchWay_r & 4'hf == blockIdx_r ? tag_2_15 : _GEN_524; // @[playground/src/noop/dcache.scala 200:{30,30}]
  wire  _GEN_2818 = 2'h3 == matchWay_r; // @[playground/src/noop/dcache.scala 200:{30,30}]
  wire [21:0] _GEN_526 = 2'h3 == matchWay_r & 4'h0 == blockIdx_r ? tag_3_0 : _GEN_525; // @[playground/src/noop/dcache.scala 200:{30,30}]
  wire [21:0] _GEN_527 = 2'h3 == matchWay_r & 4'h1 == blockIdx_r ? tag_3_1 : _GEN_526; // @[playground/src/noop/dcache.scala 200:{30,30}]
  wire [21:0] _GEN_528 = 2'h3 == matchWay_r & 4'h2 == blockIdx_r ? tag_3_2 : _GEN_527; // @[playground/src/noop/dcache.scala 200:{30,30}]
  wire [21:0] _GEN_529 = 2'h3 == matchWay_r & 4'h3 == blockIdx_r ? tag_3_3 : _GEN_528; // @[playground/src/noop/dcache.scala 200:{30,30}]
  wire [21:0] _GEN_530 = 2'h3 == matchWay_r & 4'h4 == blockIdx_r ? tag_3_4 : _GEN_529; // @[playground/src/noop/dcache.scala 200:{30,30}]
  wire [21:0] _GEN_531 = 2'h3 == matchWay_r & 4'h5 == blockIdx_r ? tag_3_5 : _GEN_530; // @[playground/src/noop/dcache.scala 200:{30,30}]
  wire [21:0] _GEN_532 = 2'h3 == matchWay_r & 4'h6 == blockIdx_r ? tag_3_6 : _GEN_531; // @[playground/src/noop/dcache.scala 200:{30,30}]
  wire [21:0] _GEN_533 = 2'h3 == matchWay_r & 4'h7 == blockIdx_r ? tag_3_7 : _GEN_532; // @[playground/src/noop/dcache.scala 200:{30,30}]
  wire [21:0] _GEN_534 = 2'h3 == matchWay_r & 4'h8 == blockIdx_r ? tag_3_8 : _GEN_533; // @[playground/src/noop/dcache.scala 200:{30,30}]
  wire [21:0] _GEN_535 = 2'h3 == matchWay_r & 4'h9 == blockIdx_r ? tag_3_9 : _GEN_534; // @[playground/src/noop/dcache.scala 200:{30,30}]
  wire [21:0] _GEN_536 = 2'h3 == matchWay_r & 4'ha == blockIdx_r ? tag_3_10 : _GEN_535; // @[playground/src/noop/dcache.scala 200:{30,30}]
  wire [21:0] _GEN_537 = 2'h3 == matchWay_r & 4'hb == blockIdx_r ? tag_3_11 : _GEN_536; // @[playground/src/noop/dcache.scala 200:{30,30}]
  wire [21:0] _GEN_538 = 2'h3 == matchWay_r & 4'hc == blockIdx_r ? tag_3_12 : _GEN_537; // @[playground/src/noop/dcache.scala 200:{30,30}]
  wire [21:0] _GEN_539 = 2'h3 == matchWay_r & 4'hd == blockIdx_r ? tag_3_13 : _GEN_538; // @[playground/src/noop/dcache.scala 200:{30,30}]
  wire [21:0] _GEN_540 = 2'h3 == matchWay_r & 4'he == blockIdx_r ? tag_3_14 : _GEN_539; // @[playground/src/noop/dcache.scala 200:{30,30}]
  wire [21:0] _GEN_541 = 2'h3 == matchWay_r & 4'hf == blockIdx_r ? tag_3_15 : _GEN_540; // @[playground/src/noop/dcache.scala 200:{30,30}]
  wire [25:0] axiWaddr_hi = {_GEN_541,blockIdx_r}; // @[playground/src/noop/dcache.scala 200:30]
  reg  axiWdataEn; // @[playground/src/noop/dcache.scala 202:34]
  wire [2:0] _GEN_542 = cur_mode_sl == 2'h3 ? 3'h5 : state; // @[playground/src/noop/dcache.scala 152:24 212:42 213:27]
  wire  _GEN_548 = 2'h0 == matchWay & _GEN_2536 ? dirty_0_1 : dirty_0_0; // @[playground/src/noop/dcache.scala 223:{31,31}]
  wire  _GEN_549 = 2'h0 == matchWay & _GEN_2539 ? dirty_0_2 : _GEN_548; // @[playground/src/noop/dcache.scala 223:{31,31}]
  wire  _GEN_550 = 2'h0 == matchWay & _GEN_2542 ? dirty_0_3 : _GEN_549; // @[playground/src/noop/dcache.scala 223:{31,31}]
  wire  _GEN_551 = 2'h0 == matchWay & _GEN_2545 ? dirty_0_4 : _GEN_550; // @[playground/src/noop/dcache.scala 223:{31,31}]
  wire  _GEN_552 = 2'h0 == matchWay & _GEN_2548 ? dirty_0_5 : _GEN_551; // @[playground/src/noop/dcache.scala 223:{31,31}]
  wire  _GEN_553 = 2'h0 == matchWay & _GEN_2551 ? dirty_0_6 : _GEN_552; // @[playground/src/noop/dcache.scala 223:{31,31}]
  wire  _GEN_554 = 2'h0 == matchWay & _GEN_2554 ? dirty_0_7 : _GEN_553; // @[playground/src/noop/dcache.scala 223:{31,31}]
  wire  _GEN_555 = 2'h0 == matchWay & _GEN_2557 ? dirty_0_8 : _GEN_554; // @[playground/src/noop/dcache.scala 223:{31,31}]
  wire  _GEN_556 = 2'h0 == matchWay & _GEN_2560 ? dirty_0_9 : _GEN_555; // @[playground/src/noop/dcache.scala 223:{31,31}]
  wire  _GEN_557 = 2'h0 == matchWay & _GEN_2563 ? dirty_0_10 : _GEN_556; // @[playground/src/noop/dcache.scala 223:{31,31}]
  wire  _GEN_558 = 2'h0 == matchWay & _GEN_2566 ? dirty_0_11 : _GEN_557; // @[playground/src/noop/dcache.scala 223:{31,31}]
  wire  _GEN_559 = 2'h0 == matchWay & _GEN_2569 ? dirty_0_12 : _GEN_558; // @[playground/src/noop/dcache.scala 223:{31,31}]
  wire  _GEN_560 = 2'h0 == matchWay & _GEN_2572 ? dirty_0_13 : _GEN_559; // @[playground/src/noop/dcache.scala 223:{31,31}]
  wire  _GEN_561 = 2'h0 == matchWay & _GEN_2575 ? dirty_0_14 : _GEN_560; // @[playground/src/noop/dcache.scala 223:{31,31}]
  wire  _GEN_562 = 2'h0 == matchWay & _GEN_2578 ? dirty_0_15 : _GEN_561; // @[playground/src/noop/dcache.scala 223:{31,31}]
  wire  _GEN_563 = 2'h1 == matchWay & _GEN_2533 ? dirty_1_0 : _GEN_562; // @[playground/src/noop/dcache.scala 223:{31,31}]
  wire  _GEN_564 = 2'h1 == matchWay & _GEN_2536 ? dirty_1_1 : _GEN_563; // @[playground/src/noop/dcache.scala 223:{31,31}]
  wire  _GEN_565 = 2'h1 == matchWay & _GEN_2539 ? dirty_1_2 : _GEN_564; // @[playground/src/noop/dcache.scala 223:{31,31}]
  wire  _GEN_566 = 2'h1 == matchWay & _GEN_2542 ? dirty_1_3 : _GEN_565; // @[playground/src/noop/dcache.scala 223:{31,31}]
  wire  _GEN_567 = 2'h1 == matchWay & _GEN_2545 ? dirty_1_4 : _GEN_566; // @[playground/src/noop/dcache.scala 223:{31,31}]
  wire  _GEN_568 = 2'h1 == matchWay & _GEN_2548 ? dirty_1_5 : _GEN_567; // @[playground/src/noop/dcache.scala 223:{31,31}]
  wire  _GEN_569 = 2'h1 == matchWay & _GEN_2551 ? dirty_1_6 : _GEN_568; // @[playground/src/noop/dcache.scala 223:{31,31}]
  wire  _GEN_570 = 2'h1 == matchWay & _GEN_2554 ? dirty_1_7 : _GEN_569; // @[playground/src/noop/dcache.scala 223:{31,31}]
  wire  _GEN_571 = 2'h1 == matchWay & _GEN_2557 ? dirty_1_8 : _GEN_570; // @[playground/src/noop/dcache.scala 223:{31,31}]
  wire  _GEN_572 = 2'h1 == matchWay & _GEN_2560 ? dirty_1_9 : _GEN_571; // @[playground/src/noop/dcache.scala 223:{31,31}]
  wire  _GEN_573 = 2'h1 == matchWay & _GEN_2563 ? dirty_1_10 : _GEN_572; // @[playground/src/noop/dcache.scala 223:{31,31}]
  wire  _GEN_574 = 2'h1 == matchWay & _GEN_2566 ? dirty_1_11 : _GEN_573; // @[playground/src/noop/dcache.scala 223:{31,31}]
  wire  _GEN_575 = 2'h1 == matchWay & _GEN_2569 ? dirty_1_12 : _GEN_574; // @[playground/src/noop/dcache.scala 223:{31,31}]
  wire  _GEN_576 = 2'h1 == matchWay & _GEN_2572 ? dirty_1_13 : _GEN_575; // @[playground/src/noop/dcache.scala 223:{31,31}]
  wire  _GEN_577 = 2'h1 == matchWay & _GEN_2575 ? dirty_1_14 : _GEN_576; // @[playground/src/noop/dcache.scala 223:{31,31}]
  wire  _GEN_578 = 2'h1 == matchWay & _GEN_2578 ? dirty_1_15 : _GEN_577; // @[playground/src/noop/dcache.scala 223:{31,31}]
  wire  _GEN_579 = 2'h2 == matchWay & _GEN_2533 ? dirty_2_0 : _GEN_578; // @[playground/src/noop/dcache.scala 223:{31,31}]
  wire  _GEN_580 = 2'h2 == matchWay & _GEN_2536 ? dirty_2_1 : _GEN_579; // @[playground/src/noop/dcache.scala 223:{31,31}]
  wire  _GEN_581 = 2'h2 == matchWay & _GEN_2539 ? dirty_2_2 : _GEN_580; // @[playground/src/noop/dcache.scala 223:{31,31}]
  wire  _GEN_582 = 2'h2 == matchWay & _GEN_2542 ? dirty_2_3 : _GEN_581; // @[playground/src/noop/dcache.scala 223:{31,31}]
  wire  _GEN_583 = 2'h2 == matchWay & _GEN_2545 ? dirty_2_4 : _GEN_582; // @[playground/src/noop/dcache.scala 223:{31,31}]
  wire  _GEN_584 = 2'h2 == matchWay & _GEN_2548 ? dirty_2_5 : _GEN_583; // @[playground/src/noop/dcache.scala 223:{31,31}]
  wire  _GEN_585 = 2'h2 == matchWay & _GEN_2551 ? dirty_2_6 : _GEN_584; // @[playground/src/noop/dcache.scala 223:{31,31}]
  wire  _GEN_586 = 2'h2 == matchWay & _GEN_2554 ? dirty_2_7 : _GEN_585; // @[playground/src/noop/dcache.scala 223:{31,31}]
  wire  _GEN_587 = 2'h2 == matchWay & _GEN_2557 ? dirty_2_8 : _GEN_586; // @[playground/src/noop/dcache.scala 223:{31,31}]
  wire  _GEN_588 = 2'h2 == matchWay & _GEN_2560 ? dirty_2_9 : _GEN_587; // @[playground/src/noop/dcache.scala 223:{31,31}]
  wire  _GEN_589 = 2'h2 == matchWay & _GEN_2563 ? dirty_2_10 : _GEN_588; // @[playground/src/noop/dcache.scala 223:{31,31}]
  wire  _GEN_590 = 2'h2 == matchWay & _GEN_2566 ? dirty_2_11 : _GEN_589; // @[playground/src/noop/dcache.scala 223:{31,31}]
  wire  _GEN_591 = 2'h2 == matchWay & _GEN_2569 ? dirty_2_12 : _GEN_590; // @[playground/src/noop/dcache.scala 223:{31,31}]
  wire  _GEN_592 = 2'h2 == matchWay & _GEN_2572 ? dirty_2_13 : _GEN_591; // @[playground/src/noop/dcache.scala 223:{31,31}]
  wire  _GEN_593 = 2'h2 == matchWay & _GEN_2575 ? dirty_2_14 : _GEN_592; // @[playground/src/noop/dcache.scala 223:{31,31}]
  wire  _GEN_594 = 2'h2 == matchWay & _GEN_2578 ? dirty_2_15 : _GEN_593; // @[playground/src/noop/dcache.scala 223:{31,31}]
  wire  _GEN_595 = 2'h3 == matchWay & _GEN_2533 ? dirty_3_0 : _GEN_594; // @[playground/src/noop/dcache.scala 223:{31,31}]
  wire  _GEN_596 = 2'h3 == matchWay & _GEN_2536 ? dirty_3_1 : _GEN_595; // @[playground/src/noop/dcache.scala 223:{31,31}]
  wire  _GEN_597 = 2'h3 == matchWay & _GEN_2539 ? dirty_3_2 : _GEN_596; // @[playground/src/noop/dcache.scala 223:{31,31}]
  wire  _GEN_598 = 2'h3 == matchWay & _GEN_2542 ? dirty_3_3 : _GEN_597; // @[playground/src/noop/dcache.scala 223:{31,31}]
  wire  _GEN_599 = 2'h3 == matchWay & _GEN_2545 ? dirty_3_4 : _GEN_598; // @[playground/src/noop/dcache.scala 223:{31,31}]
  wire  _GEN_600 = 2'h3 == matchWay & _GEN_2548 ? dirty_3_5 : _GEN_599; // @[playground/src/noop/dcache.scala 223:{31,31}]
  wire  _GEN_601 = 2'h3 == matchWay & _GEN_2551 ? dirty_3_6 : _GEN_600; // @[playground/src/noop/dcache.scala 223:{31,31}]
  wire  _GEN_602 = 2'h3 == matchWay & _GEN_2554 ? dirty_3_7 : _GEN_601; // @[playground/src/noop/dcache.scala 223:{31,31}]
  wire  _GEN_603 = 2'h3 == matchWay & _GEN_2557 ? dirty_3_8 : _GEN_602; // @[playground/src/noop/dcache.scala 223:{31,31}]
  wire  _GEN_604 = 2'h3 == matchWay & _GEN_2560 ? dirty_3_9 : _GEN_603; // @[playground/src/noop/dcache.scala 223:{31,31}]
  wire  _GEN_605 = 2'h3 == matchWay & _GEN_2563 ? dirty_3_10 : _GEN_604; // @[playground/src/noop/dcache.scala 223:{31,31}]
  wire  _GEN_606 = 2'h3 == matchWay & _GEN_2566 ? dirty_3_11 : _GEN_605; // @[playground/src/noop/dcache.scala 223:{31,31}]
  wire  _GEN_607 = 2'h3 == matchWay & _GEN_2569 ? dirty_3_12 : _GEN_606; // @[playground/src/noop/dcache.scala 223:{31,31}]
  wire  _GEN_608 = 2'h3 == matchWay & _GEN_2572 ? dirty_3_13 : _GEN_607; // @[playground/src/noop/dcache.scala 223:{31,31}]
  wire  _GEN_609 = 2'h3 == matchWay & _GEN_2575 ? dirty_3_14 : _GEN_608; // @[playground/src/noop/dcache.scala 223:{31,31}]
  wire  _GEN_610 = 2'h3 == matchWay & _GEN_2578 ? dirty_3_15 : _GEN_609; // @[playground/src/noop/dcache.scala 223:{31,31}]
  wire [2:0] _GEN_611 = _GEN_610 ? 3'h3 : 3'h1; // @[playground/src/noop/dcache.scala 223:31 224:27 227:27]
  wire  _GEN_612 = _GEN_610 | axiWaddrEn; // @[playground/src/noop/dcache.scala 223:31 225:32 199:34]
  wire  _GEN_613 = _GEN_610 ? axiRaddrEn : 1'h1; // @[playground/src/noop/dcache.scala 223:31 196:34 228:32]
  wire [2:0] _GEN_614 = cacheHit ? _GEN_542 : _GEN_611; // @[playground/src/noop/dcache.scala 211:33]
  wire  _GEN_616 = cacheHit ? _T_73 : 1'h1; // @[playground/src/noop/dcache.scala 211:33 231:25]
  wire  _GEN_619 = cacheHit ? axiWaddrEn : _GEN_612; // @[playground/src/noop/dcache.scala 211:33 199:34]
  wire  _GEN_620 = cacheHit ? axiRaddrEn : _GEN_613; // @[playground/src/noop/dcache.scala 211:33 196:34]
  wire  _GEN_622 = ~hs_in & _io_dcRW_ready_T ? 1'h0 : cacheHit; // @[playground/src/noop/dcache.scala 101:13 209:42]
  wire  _GEN_629 = flush_r | io_flush ? 1'h0 : _GEN_622; // @[playground/src/noop/dcache.scala 101:13 207:38]
  wire  _GEN_637 = axiRaddrEn & io_dataAxi_ra_ready | axiRdataEn; // @[playground/src/noop/dcache.scala 236:52 239:28 198:34]
  wire [2:0] _offset_T_1 = offset + 3'h1; // @[playground/src/noop/dcache.scala 244:34]
  wire [63:0] _GEN_639 = offset[0] ? rdatabuf : io_dataAxi_rd_bits_data; // @[playground/src/noop/dcache.scala 245:32 111:34 248:30]
  wire  _GEN_2977 = 4'h0 == pre_blockIdx; // @[playground/src/noop/dcache.scala 252:{51,51} 88:26]
  wire [21:0] _GEN_640 = _GEN_2724 & 4'h0 == pre_blockIdx ? pre_tag : tag_0_0; // @[playground/src/noop/dcache.scala 252:{51,51} 88:26]
  wire  _GEN_2979 = 4'h1 == pre_blockIdx; // @[playground/src/noop/dcache.scala 252:{51,51} 88:26]
  wire [21:0] _GEN_641 = _GEN_2724 & 4'h1 == pre_blockIdx ? pre_tag : tag_0_1; // @[playground/src/noop/dcache.scala 252:{51,51} 88:26]
  wire  _GEN_2981 = 4'h2 == pre_blockIdx; // @[playground/src/noop/dcache.scala 252:{51,51} 88:26]
  wire [21:0] _GEN_642 = _GEN_2724 & 4'h2 == pre_blockIdx ? pre_tag : tag_0_2; // @[playground/src/noop/dcache.scala 252:{51,51} 88:26]
  wire  _GEN_2983 = 4'h3 == pre_blockIdx; // @[playground/src/noop/dcache.scala 252:{51,51} 88:26]
  wire [21:0] _GEN_643 = _GEN_2724 & 4'h3 == pre_blockIdx ? pre_tag : tag_0_3; // @[playground/src/noop/dcache.scala 252:{51,51} 88:26]
  wire  _GEN_2985 = 4'h4 == pre_blockIdx; // @[playground/src/noop/dcache.scala 252:{51,51} 88:26]
  wire [21:0] _GEN_644 = _GEN_2724 & 4'h4 == pre_blockIdx ? pre_tag : tag_0_4; // @[playground/src/noop/dcache.scala 252:{51,51} 88:26]
  wire  _GEN_2987 = 4'h5 == pre_blockIdx; // @[playground/src/noop/dcache.scala 252:{51,51} 88:26]
  wire [21:0] _GEN_645 = _GEN_2724 & 4'h5 == pre_blockIdx ? pre_tag : tag_0_5; // @[playground/src/noop/dcache.scala 252:{51,51} 88:26]
  wire  _GEN_2989 = 4'h6 == pre_blockIdx; // @[playground/src/noop/dcache.scala 252:{51,51} 88:26]
  wire [21:0] _GEN_646 = _GEN_2724 & 4'h6 == pre_blockIdx ? pre_tag : tag_0_6; // @[playground/src/noop/dcache.scala 252:{51,51} 88:26]
  wire  _GEN_2991 = 4'h7 == pre_blockIdx; // @[playground/src/noop/dcache.scala 252:{51,51} 88:26]
  wire [21:0] _GEN_647 = _GEN_2724 & 4'h7 == pre_blockIdx ? pre_tag : tag_0_7; // @[playground/src/noop/dcache.scala 252:{51,51} 88:26]
  wire  _GEN_2993 = 4'h8 == pre_blockIdx; // @[playground/src/noop/dcache.scala 252:{51,51} 88:26]
  wire [21:0] _GEN_648 = _GEN_2724 & 4'h8 == pre_blockIdx ? pre_tag : tag_0_8; // @[playground/src/noop/dcache.scala 252:{51,51} 88:26]
  wire  _GEN_2995 = 4'h9 == pre_blockIdx; // @[playground/src/noop/dcache.scala 252:{51,51} 88:26]
  wire [21:0] _GEN_649 = _GEN_2724 & 4'h9 == pre_blockIdx ? pre_tag : tag_0_9; // @[playground/src/noop/dcache.scala 252:{51,51} 88:26]
  wire  _GEN_2997 = 4'ha == pre_blockIdx; // @[playground/src/noop/dcache.scala 252:{51,51} 88:26]
  wire [21:0] _GEN_650 = _GEN_2724 & 4'ha == pre_blockIdx ? pre_tag : tag_0_10; // @[playground/src/noop/dcache.scala 252:{51,51} 88:26]
  wire  _GEN_2999 = 4'hb == pre_blockIdx; // @[playground/src/noop/dcache.scala 252:{51,51} 88:26]
  wire [21:0] _GEN_651 = _GEN_2724 & 4'hb == pre_blockIdx ? pre_tag : tag_0_11; // @[playground/src/noop/dcache.scala 252:{51,51} 88:26]
  wire  _GEN_3001 = 4'hc == pre_blockIdx; // @[playground/src/noop/dcache.scala 252:{51,51} 88:26]
  wire [21:0] _GEN_652 = _GEN_2724 & 4'hc == pre_blockIdx ? pre_tag : tag_0_12; // @[playground/src/noop/dcache.scala 252:{51,51} 88:26]
  wire  _GEN_3003 = 4'hd == pre_blockIdx; // @[playground/src/noop/dcache.scala 252:{51,51} 88:26]
  wire [21:0] _GEN_653 = _GEN_2724 & 4'hd == pre_blockIdx ? pre_tag : tag_0_13; // @[playground/src/noop/dcache.scala 252:{51,51} 88:26]
  wire  _GEN_3005 = 4'he == pre_blockIdx; // @[playground/src/noop/dcache.scala 252:{51,51} 88:26]
  wire [21:0] _GEN_654 = _GEN_2724 & 4'he == pre_blockIdx ? pre_tag : tag_0_14; // @[playground/src/noop/dcache.scala 252:{51,51} 88:26]
  wire  _GEN_3007 = 4'hf == pre_blockIdx; // @[playground/src/noop/dcache.scala 252:{51,51} 88:26]
  wire [21:0] _GEN_655 = _GEN_2724 & 4'hf == pre_blockIdx ? pre_tag : tag_0_15; // @[playground/src/noop/dcache.scala 252:{51,51} 88:26]
  wire [21:0] _GEN_656 = _GEN_2754 & 4'h0 == pre_blockIdx ? pre_tag : tag_1_0; // @[playground/src/noop/dcache.scala 252:{51,51} 88:26]
  wire [21:0] _GEN_657 = _GEN_2754 & 4'h1 == pre_blockIdx ? pre_tag : tag_1_1; // @[playground/src/noop/dcache.scala 252:{51,51} 88:26]
  wire [21:0] _GEN_658 = _GEN_2754 & 4'h2 == pre_blockIdx ? pre_tag : tag_1_2; // @[playground/src/noop/dcache.scala 252:{51,51} 88:26]
  wire [21:0] _GEN_659 = _GEN_2754 & 4'h3 == pre_blockIdx ? pre_tag : tag_1_3; // @[playground/src/noop/dcache.scala 252:{51,51} 88:26]
  wire [21:0] _GEN_660 = _GEN_2754 & 4'h4 == pre_blockIdx ? pre_tag : tag_1_4; // @[playground/src/noop/dcache.scala 252:{51,51} 88:26]
  wire [21:0] _GEN_661 = _GEN_2754 & 4'h5 == pre_blockIdx ? pre_tag : tag_1_5; // @[playground/src/noop/dcache.scala 252:{51,51} 88:26]
  wire [21:0] _GEN_662 = _GEN_2754 & 4'h6 == pre_blockIdx ? pre_tag : tag_1_6; // @[playground/src/noop/dcache.scala 252:{51,51} 88:26]
  wire [21:0] _GEN_663 = _GEN_2754 & 4'h7 == pre_blockIdx ? pre_tag : tag_1_7; // @[playground/src/noop/dcache.scala 252:{51,51} 88:26]
  wire [21:0] _GEN_664 = _GEN_2754 & 4'h8 == pre_blockIdx ? pre_tag : tag_1_8; // @[playground/src/noop/dcache.scala 252:{51,51} 88:26]
  wire [21:0] _GEN_665 = _GEN_2754 & 4'h9 == pre_blockIdx ? pre_tag : tag_1_9; // @[playground/src/noop/dcache.scala 252:{51,51} 88:26]
  wire [21:0] _GEN_666 = _GEN_2754 & 4'ha == pre_blockIdx ? pre_tag : tag_1_10; // @[playground/src/noop/dcache.scala 252:{51,51} 88:26]
  wire [21:0] _GEN_667 = _GEN_2754 & 4'hb == pre_blockIdx ? pre_tag : tag_1_11; // @[playground/src/noop/dcache.scala 252:{51,51} 88:26]
  wire [21:0] _GEN_668 = _GEN_2754 & 4'hc == pre_blockIdx ? pre_tag : tag_1_12; // @[playground/src/noop/dcache.scala 252:{51,51} 88:26]
  wire [21:0] _GEN_669 = _GEN_2754 & 4'hd == pre_blockIdx ? pre_tag : tag_1_13; // @[playground/src/noop/dcache.scala 252:{51,51} 88:26]
  wire [21:0] _GEN_670 = _GEN_2754 & 4'he == pre_blockIdx ? pre_tag : tag_1_14; // @[playground/src/noop/dcache.scala 252:{51,51} 88:26]
  wire [21:0] _GEN_671 = _GEN_2754 & 4'hf == pre_blockIdx ? pre_tag : tag_1_15; // @[playground/src/noop/dcache.scala 252:{51,51} 88:26]
  wire [21:0] _GEN_672 = _GEN_2786 & 4'h0 == pre_blockIdx ? pre_tag : tag_2_0; // @[playground/src/noop/dcache.scala 252:{51,51} 88:26]
  wire [21:0] _GEN_673 = _GEN_2786 & 4'h1 == pre_blockIdx ? pre_tag : tag_2_1; // @[playground/src/noop/dcache.scala 252:{51,51} 88:26]
  wire [21:0] _GEN_674 = _GEN_2786 & 4'h2 == pre_blockIdx ? pre_tag : tag_2_2; // @[playground/src/noop/dcache.scala 252:{51,51} 88:26]
  wire [21:0] _GEN_675 = _GEN_2786 & 4'h3 == pre_blockIdx ? pre_tag : tag_2_3; // @[playground/src/noop/dcache.scala 252:{51,51} 88:26]
  wire [21:0] _GEN_676 = _GEN_2786 & 4'h4 == pre_blockIdx ? pre_tag : tag_2_4; // @[playground/src/noop/dcache.scala 252:{51,51} 88:26]
  wire [21:0] _GEN_677 = _GEN_2786 & 4'h5 == pre_blockIdx ? pre_tag : tag_2_5; // @[playground/src/noop/dcache.scala 252:{51,51} 88:26]
  wire [21:0] _GEN_678 = _GEN_2786 & 4'h6 == pre_blockIdx ? pre_tag : tag_2_6; // @[playground/src/noop/dcache.scala 252:{51,51} 88:26]
  wire [21:0] _GEN_679 = _GEN_2786 & 4'h7 == pre_blockIdx ? pre_tag : tag_2_7; // @[playground/src/noop/dcache.scala 252:{51,51} 88:26]
  wire [21:0] _GEN_680 = _GEN_2786 & 4'h8 == pre_blockIdx ? pre_tag : tag_2_8; // @[playground/src/noop/dcache.scala 252:{51,51} 88:26]
  wire [21:0] _GEN_681 = _GEN_2786 & 4'h9 == pre_blockIdx ? pre_tag : tag_2_9; // @[playground/src/noop/dcache.scala 252:{51,51} 88:26]
  wire [21:0] _GEN_682 = _GEN_2786 & 4'ha == pre_blockIdx ? pre_tag : tag_2_10; // @[playground/src/noop/dcache.scala 252:{51,51} 88:26]
  wire [21:0] _GEN_683 = _GEN_2786 & 4'hb == pre_blockIdx ? pre_tag : tag_2_11; // @[playground/src/noop/dcache.scala 252:{51,51} 88:26]
  wire [21:0] _GEN_684 = _GEN_2786 & 4'hc == pre_blockIdx ? pre_tag : tag_2_12; // @[playground/src/noop/dcache.scala 252:{51,51} 88:26]
  wire [21:0] _GEN_685 = _GEN_2786 & 4'hd == pre_blockIdx ? pre_tag : tag_2_13; // @[playground/src/noop/dcache.scala 252:{51,51} 88:26]
  wire [21:0] _GEN_686 = _GEN_2786 & 4'he == pre_blockIdx ? pre_tag : tag_2_14; // @[playground/src/noop/dcache.scala 252:{51,51} 88:26]
  wire [21:0] _GEN_687 = _GEN_2786 & 4'hf == pre_blockIdx ? pre_tag : tag_2_15; // @[playground/src/noop/dcache.scala 252:{51,51} 88:26]
  wire [21:0] _GEN_688 = _GEN_2818 & 4'h0 == pre_blockIdx ? pre_tag : tag_3_0; // @[playground/src/noop/dcache.scala 252:{51,51} 88:26]
  wire [21:0] _GEN_689 = _GEN_2818 & 4'h1 == pre_blockIdx ? pre_tag : tag_3_1; // @[playground/src/noop/dcache.scala 252:{51,51} 88:26]
  wire [21:0] _GEN_690 = _GEN_2818 & 4'h2 == pre_blockIdx ? pre_tag : tag_3_2; // @[playground/src/noop/dcache.scala 252:{51,51} 88:26]
  wire [21:0] _GEN_691 = _GEN_2818 & 4'h3 == pre_blockIdx ? pre_tag : tag_3_3; // @[playground/src/noop/dcache.scala 252:{51,51} 88:26]
  wire [21:0] _GEN_692 = _GEN_2818 & 4'h4 == pre_blockIdx ? pre_tag : tag_3_4; // @[playground/src/noop/dcache.scala 252:{51,51} 88:26]
  wire [21:0] _GEN_693 = _GEN_2818 & 4'h5 == pre_blockIdx ? pre_tag : tag_3_5; // @[playground/src/noop/dcache.scala 252:{51,51} 88:26]
  wire [21:0] _GEN_694 = _GEN_2818 & 4'h6 == pre_blockIdx ? pre_tag : tag_3_6; // @[playground/src/noop/dcache.scala 252:{51,51} 88:26]
  wire [21:0] _GEN_695 = _GEN_2818 & 4'h7 == pre_blockIdx ? pre_tag : tag_3_7; // @[playground/src/noop/dcache.scala 252:{51,51} 88:26]
  wire [21:0] _GEN_696 = _GEN_2818 & 4'h8 == pre_blockIdx ? pre_tag : tag_3_8; // @[playground/src/noop/dcache.scala 252:{51,51} 88:26]
  wire [21:0] _GEN_697 = _GEN_2818 & 4'h9 == pre_blockIdx ? pre_tag : tag_3_9; // @[playground/src/noop/dcache.scala 252:{51,51} 88:26]
  wire [21:0] _GEN_698 = _GEN_2818 & 4'ha == pre_blockIdx ? pre_tag : tag_3_10; // @[playground/src/noop/dcache.scala 252:{51,51} 88:26]
  wire [21:0] _GEN_699 = _GEN_2818 & 4'hb == pre_blockIdx ? pre_tag : tag_3_11; // @[playground/src/noop/dcache.scala 252:{51,51} 88:26]
  wire [21:0] _GEN_700 = _GEN_2818 & 4'hc == pre_blockIdx ? pre_tag : tag_3_12; // @[playground/src/noop/dcache.scala 252:{51,51} 88:26]
  wire [21:0] _GEN_701 = _GEN_2818 & 4'hd == pre_blockIdx ? pre_tag : tag_3_13; // @[playground/src/noop/dcache.scala 252:{51,51} 88:26]
  wire [21:0] _GEN_702 = _GEN_2818 & 4'he == pre_blockIdx ? pre_tag : tag_3_14; // @[playground/src/noop/dcache.scala 252:{51,51} 88:26]
  wire [21:0] _GEN_703 = _GEN_2818 & 4'hf == pre_blockIdx ? pre_tag : tag_3_15; // @[playground/src/noop/dcache.scala 252:{51,51} 88:26]
  wire  _GEN_704 = _GEN_2724 & _GEN_2977 | valid_0_0; // @[playground/src/noop/dcache.scala 253:{53,53} 89:26]
  wire  _GEN_705 = _GEN_2724 & _GEN_2979 | valid_0_1; // @[playground/src/noop/dcache.scala 253:{53,53} 89:26]
  wire  _GEN_706 = _GEN_2724 & _GEN_2981 | valid_0_2; // @[playground/src/noop/dcache.scala 253:{53,53} 89:26]
  wire  _GEN_707 = _GEN_2724 & _GEN_2983 | valid_0_3; // @[playground/src/noop/dcache.scala 253:{53,53} 89:26]
  wire  _GEN_708 = _GEN_2724 & _GEN_2985 | valid_0_4; // @[playground/src/noop/dcache.scala 253:{53,53} 89:26]
  wire  _GEN_709 = _GEN_2724 & _GEN_2987 | valid_0_5; // @[playground/src/noop/dcache.scala 253:{53,53} 89:26]
  wire  _GEN_710 = _GEN_2724 & _GEN_2989 | valid_0_6; // @[playground/src/noop/dcache.scala 253:{53,53} 89:26]
  wire  _GEN_711 = _GEN_2724 & _GEN_2991 | valid_0_7; // @[playground/src/noop/dcache.scala 253:{53,53} 89:26]
  wire  _GEN_712 = _GEN_2724 & _GEN_2993 | valid_0_8; // @[playground/src/noop/dcache.scala 253:{53,53} 89:26]
  wire  _GEN_713 = _GEN_2724 & _GEN_2995 | valid_0_9; // @[playground/src/noop/dcache.scala 253:{53,53} 89:26]
  wire  _GEN_714 = _GEN_2724 & _GEN_2997 | valid_0_10; // @[playground/src/noop/dcache.scala 253:{53,53} 89:26]
  wire  _GEN_715 = _GEN_2724 & _GEN_2999 | valid_0_11; // @[playground/src/noop/dcache.scala 253:{53,53} 89:26]
  wire  _GEN_716 = _GEN_2724 & _GEN_3001 | valid_0_12; // @[playground/src/noop/dcache.scala 253:{53,53} 89:26]
  wire  _GEN_717 = _GEN_2724 & _GEN_3003 | valid_0_13; // @[playground/src/noop/dcache.scala 253:{53,53} 89:26]
  wire  _GEN_718 = _GEN_2724 & _GEN_3005 | valid_0_14; // @[playground/src/noop/dcache.scala 253:{53,53} 89:26]
  wire  _GEN_719 = _GEN_2724 & _GEN_3007 | valid_0_15; // @[playground/src/noop/dcache.scala 253:{53,53} 89:26]
  wire  _GEN_720 = _GEN_2754 & _GEN_2977 | valid_1_0; // @[playground/src/noop/dcache.scala 253:{53,53} 89:26]
  wire  _GEN_721 = _GEN_2754 & _GEN_2979 | valid_1_1; // @[playground/src/noop/dcache.scala 253:{53,53} 89:26]
  wire  _GEN_722 = _GEN_2754 & _GEN_2981 | valid_1_2; // @[playground/src/noop/dcache.scala 253:{53,53} 89:26]
  wire  _GEN_723 = _GEN_2754 & _GEN_2983 | valid_1_3; // @[playground/src/noop/dcache.scala 253:{53,53} 89:26]
  wire  _GEN_724 = _GEN_2754 & _GEN_2985 | valid_1_4; // @[playground/src/noop/dcache.scala 253:{53,53} 89:26]
  wire  _GEN_725 = _GEN_2754 & _GEN_2987 | valid_1_5; // @[playground/src/noop/dcache.scala 253:{53,53} 89:26]
  wire  _GEN_726 = _GEN_2754 & _GEN_2989 | valid_1_6; // @[playground/src/noop/dcache.scala 253:{53,53} 89:26]
  wire  _GEN_727 = _GEN_2754 & _GEN_2991 | valid_1_7; // @[playground/src/noop/dcache.scala 253:{53,53} 89:26]
  wire  _GEN_728 = _GEN_2754 & _GEN_2993 | valid_1_8; // @[playground/src/noop/dcache.scala 253:{53,53} 89:26]
  wire  _GEN_729 = _GEN_2754 & _GEN_2995 | valid_1_9; // @[playground/src/noop/dcache.scala 253:{53,53} 89:26]
  wire  _GEN_730 = _GEN_2754 & _GEN_2997 | valid_1_10; // @[playground/src/noop/dcache.scala 253:{53,53} 89:26]
  wire  _GEN_731 = _GEN_2754 & _GEN_2999 | valid_1_11; // @[playground/src/noop/dcache.scala 253:{53,53} 89:26]
  wire  _GEN_732 = _GEN_2754 & _GEN_3001 | valid_1_12; // @[playground/src/noop/dcache.scala 253:{53,53} 89:26]
  wire  _GEN_733 = _GEN_2754 & _GEN_3003 | valid_1_13; // @[playground/src/noop/dcache.scala 253:{53,53} 89:26]
  wire  _GEN_734 = _GEN_2754 & _GEN_3005 | valid_1_14; // @[playground/src/noop/dcache.scala 253:{53,53} 89:26]
  wire  _GEN_735 = _GEN_2754 & _GEN_3007 | valid_1_15; // @[playground/src/noop/dcache.scala 253:{53,53} 89:26]
  wire  _GEN_736 = _GEN_2786 & _GEN_2977 | valid_2_0; // @[playground/src/noop/dcache.scala 253:{53,53} 89:26]
  wire  _GEN_737 = _GEN_2786 & _GEN_2979 | valid_2_1; // @[playground/src/noop/dcache.scala 253:{53,53} 89:26]
  wire  _GEN_738 = _GEN_2786 & _GEN_2981 | valid_2_2; // @[playground/src/noop/dcache.scala 253:{53,53} 89:26]
  wire  _GEN_739 = _GEN_2786 & _GEN_2983 | valid_2_3; // @[playground/src/noop/dcache.scala 253:{53,53} 89:26]
  wire  _GEN_740 = _GEN_2786 & _GEN_2985 | valid_2_4; // @[playground/src/noop/dcache.scala 253:{53,53} 89:26]
  wire  _GEN_741 = _GEN_2786 & _GEN_2987 | valid_2_5; // @[playground/src/noop/dcache.scala 253:{53,53} 89:26]
  wire  _GEN_742 = _GEN_2786 & _GEN_2989 | valid_2_6; // @[playground/src/noop/dcache.scala 253:{53,53} 89:26]
  wire  _GEN_743 = _GEN_2786 & _GEN_2991 | valid_2_7; // @[playground/src/noop/dcache.scala 253:{53,53} 89:26]
  wire  _GEN_744 = _GEN_2786 & _GEN_2993 | valid_2_8; // @[playground/src/noop/dcache.scala 253:{53,53} 89:26]
  wire  _GEN_745 = _GEN_2786 & _GEN_2995 | valid_2_9; // @[playground/src/noop/dcache.scala 253:{53,53} 89:26]
  wire  _GEN_746 = _GEN_2786 & _GEN_2997 | valid_2_10; // @[playground/src/noop/dcache.scala 253:{53,53} 89:26]
  wire  _GEN_747 = _GEN_2786 & _GEN_2999 | valid_2_11; // @[playground/src/noop/dcache.scala 253:{53,53} 89:26]
  wire  _GEN_748 = _GEN_2786 & _GEN_3001 | valid_2_12; // @[playground/src/noop/dcache.scala 253:{53,53} 89:26]
  wire  _GEN_749 = _GEN_2786 & _GEN_3003 | valid_2_13; // @[playground/src/noop/dcache.scala 253:{53,53} 89:26]
  wire  _GEN_750 = _GEN_2786 & _GEN_3005 | valid_2_14; // @[playground/src/noop/dcache.scala 253:{53,53} 89:26]
  wire  _GEN_751 = _GEN_2786 & _GEN_3007 | valid_2_15; // @[playground/src/noop/dcache.scala 253:{53,53} 89:26]
  wire  _GEN_752 = _GEN_2818 & _GEN_2977 | valid_3_0; // @[playground/src/noop/dcache.scala 253:{53,53} 89:26]
  wire  _GEN_753 = _GEN_2818 & _GEN_2979 | valid_3_1; // @[playground/src/noop/dcache.scala 253:{53,53} 89:26]
  wire  _GEN_754 = _GEN_2818 & _GEN_2981 | valid_3_2; // @[playground/src/noop/dcache.scala 253:{53,53} 89:26]
  wire  _GEN_755 = _GEN_2818 & _GEN_2983 | valid_3_3; // @[playground/src/noop/dcache.scala 253:{53,53} 89:26]
  wire  _GEN_756 = _GEN_2818 & _GEN_2985 | valid_3_4; // @[playground/src/noop/dcache.scala 253:{53,53} 89:26]
  wire  _GEN_757 = _GEN_2818 & _GEN_2987 | valid_3_5; // @[playground/src/noop/dcache.scala 253:{53,53} 89:26]
  wire  _GEN_758 = _GEN_2818 & _GEN_2989 | valid_3_6; // @[playground/src/noop/dcache.scala 253:{53,53} 89:26]
  wire  _GEN_759 = _GEN_2818 & _GEN_2991 | valid_3_7; // @[playground/src/noop/dcache.scala 253:{53,53} 89:26]
  wire  _GEN_760 = _GEN_2818 & _GEN_2993 | valid_3_8; // @[playground/src/noop/dcache.scala 253:{53,53} 89:26]
  wire  _GEN_761 = _GEN_2818 & _GEN_2995 | valid_3_9; // @[playground/src/noop/dcache.scala 253:{53,53} 89:26]
  wire  _GEN_762 = _GEN_2818 & _GEN_2997 | valid_3_10; // @[playground/src/noop/dcache.scala 253:{53,53} 89:26]
  wire  _GEN_763 = _GEN_2818 & _GEN_2999 | valid_3_11; // @[playground/src/noop/dcache.scala 253:{53,53} 89:26]
  wire  _GEN_764 = _GEN_2818 & _GEN_3001 | valid_3_12; // @[playground/src/noop/dcache.scala 253:{53,53} 89:26]
  wire  _GEN_765 = _GEN_2818 & _GEN_3003 | valid_3_13; // @[playground/src/noop/dcache.scala 253:{53,53} 89:26]
  wire  _GEN_766 = _GEN_2818 & _GEN_3005 | valid_3_14; // @[playground/src/noop/dcache.scala 253:{53,53} 89:26]
  wire  _GEN_767 = _GEN_2818 & _GEN_3007 | valid_3_15; // @[playground/src/noop/dcache.scala 253:{53,53} 89:26]
  wire  _GEN_768 = io_dataAxi_rd_bits_last ? 1'h0 : axiRdataEn; // @[playground/src/noop/dcache.scala 250:46 251:32 198:34]
  wire [21:0] _GEN_769 = io_dataAxi_rd_bits_last ? _GEN_640 : tag_0_0; // @[playground/src/noop/dcache.scala 250:46 88:26]
  wire [21:0] _GEN_770 = io_dataAxi_rd_bits_last ? _GEN_641 : tag_0_1; // @[playground/src/noop/dcache.scala 250:46 88:26]
  wire [21:0] _GEN_771 = io_dataAxi_rd_bits_last ? _GEN_642 : tag_0_2; // @[playground/src/noop/dcache.scala 250:46 88:26]
  wire [21:0] _GEN_772 = io_dataAxi_rd_bits_last ? _GEN_643 : tag_0_3; // @[playground/src/noop/dcache.scala 250:46 88:26]
  wire [21:0] _GEN_773 = io_dataAxi_rd_bits_last ? _GEN_644 : tag_0_4; // @[playground/src/noop/dcache.scala 250:46 88:26]
  wire [21:0] _GEN_774 = io_dataAxi_rd_bits_last ? _GEN_645 : tag_0_5; // @[playground/src/noop/dcache.scala 250:46 88:26]
  wire [21:0] _GEN_775 = io_dataAxi_rd_bits_last ? _GEN_646 : tag_0_6; // @[playground/src/noop/dcache.scala 250:46 88:26]
  wire [21:0] _GEN_776 = io_dataAxi_rd_bits_last ? _GEN_647 : tag_0_7; // @[playground/src/noop/dcache.scala 250:46 88:26]
  wire [21:0] _GEN_777 = io_dataAxi_rd_bits_last ? _GEN_648 : tag_0_8; // @[playground/src/noop/dcache.scala 250:46 88:26]
  wire [21:0] _GEN_778 = io_dataAxi_rd_bits_last ? _GEN_649 : tag_0_9; // @[playground/src/noop/dcache.scala 250:46 88:26]
  wire [21:0] _GEN_779 = io_dataAxi_rd_bits_last ? _GEN_650 : tag_0_10; // @[playground/src/noop/dcache.scala 250:46 88:26]
  wire [21:0] _GEN_780 = io_dataAxi_rd_bits_last ? _GEN_651 : tag_0_11; // @[playground/src/noop/dcache.scala 250:46 88:26]
  wire [21:0] _GEN_781 = io_dataAxi_rd_bits_last ? _GEN_652 : tag_0_12; // @[playground/src/noop/dcache.scala 250:46 88:26]
  wire [21:0] _GEN_782 = io_dataAxi_rd_bits_last ? _GEN_653 : tag_0_13; // @[playground/src/noop/dcache.scala 250:46 88:26]
  wire [21:0] _GEN_783 = io_dataAxi_rd_bits_last ? _GEN_654 : tag_0_14; // @[playground/src/noop/dcache.scala 250:46 88:26]
  wire [21:0] _GEN_784 = io_dataAxi_rd_bits_last ? _GEN_655 : tag_0_15; // @[playground/src/noop/dcache.scala 250:46 88:26]
  wire [21:0] _GEN_785 = io_dataAxi_rd_bits_last ? _GEN_656 : tag_1_0; // @[playground/src/noop/dcache.scala 250:46 88:26]
  wire [21:0] _GEN_786 = io_dataAxi_rd_bits_last ? _GEN_657 : tag_1_1; // @[playground/src/noop/dcache.scala 250:46 88:26]
  wire [21:0] _GEN_787 = io_dataAxi_rd_bits_last ? _GEN_658 : tag_1_2; // @[playground/src/noop/dcache.scala 250:46 88:26]
  wire [21:0] _GEN_788 = io_dataAxi_rd_bits_last ? _GEN_659 : tag_1_3; // @[playground/src/noop/dcache.scala 250:46 88:26]
  wire [21:0] _GEN_789 = io_dataAxi_rd_bits_last ? _GEN_660 : tag_1_4; // @[playground/src/noop/dcache.scala 250:46 88:26]
  wire [21:0] _GEN_790 = io_dataAxi_rd_bits_last ? _GEN_661 : tag_1_5; // @[playground/src/noop/dcache.scala 250:46 88:26]
  wire [21:0] _GEN_791 = io_dataAxi_rd_bits_last ? _GEN_662 : tag_1_6; // @[playground/src/noop/dcache.scala 250:46 88:26]
  wire [21:0] _GEN_792 = io_dataAxi_rd_bits_last ? _GEN_663 : tag_1_7; // @[playground/src/noop/dcache.scala 250:46 88:26]
  wire [21:0] _GEN_793 = io_dataAxi_rd_bits_last ? _GEN_664 : tag_1_8; // @[playground/src/noop/dcache.scala 250:46 88:26]
  wire [21:0] _GEN_794 = io_dataAxi_rd_bits_last ? _GEN_665 : tag_1_9; // @[playground/src/noop/dcache.scala 250:46 88:26]
  wire [21:0] _GEN_795 = io_dataAxi_rd_bits_last ? _GEN_666 : tag_1_10; // @[playground/src/noop/dcache.scala 250:46 88:26]
  wire [21:0] _GEN_796 = io_dataAxi_rd_bits_last ? _GEN_667 : tag_1_11; // @[playground/src/noop/dcache.scala 250:46 88:26]
  wire [21:0] _GEN_797 = io_dataAxi_rd_bits_last ? _GEN_668 : tag_1_12; // @[playground/src/noop/dcache.scala 250:46 88:26]
  wire [21:0] _GEN_798 = io_dataAxi_rd_bits_last ? _GEN_669 : tag_1_13; // @[playground/src/noop/dcache.scala 250:46 88:26]
  wire [21:0] _GEN_799 = io_dataAxi_rd_bits_last ? _GEN_670 : tag_1_14; // @[playground/src/noop/dcache.scala 250:46 88:26]
  wire [21:0] _GEN_800 = io_dataAxi_rd_bits_last ? _GEN_671 : tag_1_15; // @[playground/src/noop/dcache.scala 250:46 88:26]
  wire [21:0] _GEN_801 = io_dataAxi_rd_bits_last ? _GEN_672 : tag_2_0; // @[playground/src/noop/dcache.scala 250:46 88:26]
  wire [21:0] _GEN_802 = io_dataAxi_rd_bits_last ? _GEN_673 : tag_2_1; // @[playground/src/noop/dcache.scala 250:46 88:26]
  wire [21:0] _GEN_803 = io_dataAxi_rd_bits_last ? _GEN_674 : tag_2_2; // @[playground/src/noop/dcache.scala 250:46 88:26]
  wire [21:0] _GEN_804 = io_dataAxi_rd_bits_last ? _GEN_675 : tag_2_3; // @[playground/src/noop/dcache.scala 250:46 88:26]
  wire [21:0] _GEN_805 = io_dataAxi_rd_bits_last ? _GEN_676 : tag_2_4; // @[playground/src/noop/dcache.scala 250:46 88:26]
  wire [21:0] _GEN_806 = io_dataAxi_rd_bits_last ? _GEN_677 : tag_2_5; // @[playground/src/noop/dcache.scala 250:46 88:26]
  wire [21:0] _GEN_807 = io_dataAxi_rd_bits_last ? _GEN_678 : tag_2_6; // @[playground/src/noop/dcache.scala 250:46 88:26]
  wire [21:0] _GEN_808 = io_dataAxi_rd_bits_last ? _GEN_679 : tag_2_7; // @[playground/src/noop/dcache.scala 250:46 88:26]
  wire [21:0] _GEN_809 = io_dataAxi_rd_bits_last ? _GEN_680 : tag_2_8; // @[playground/src/noop/dcache.scala 250:46 88:26]
  wire [21:0] _GEN_810 = io_dataAxi_rd_bits_last ? _GEN_681 : tag_2_9; // @[playground/src/noop/dcache.scala 250:46 88:26]
  wire [21:0] _GEN_811 = io_dataAxi_rd_bits_last ? _GEN_682 : tag_2_10; // @[playground/src/noop/dcache.scala 250:46 88:26]
  wire [21:0] _GEN_812 = io_dataAxi_rd_bits_last ? _GEN_683 : tag_2_11; // @[playground/src/noop/dcache.scala 250:46 88:26]
  wire [21:0] _GEN_813 = io_dataAxi_rd_bits_last ? _GEN_684 : tag_2_12; // @[playground/src/noop/dcache.scala 250:46 88:26]
  wire [21:0] _GEN_814 = io_dataAxi_rd_bits_last ? _GEN_685 : tag_2_13; // @[playground/src/noop/dcache.scala 250:46 88:26]
  wire [21:0] _GEN_815 = io_dataAxi_rd_bits_last ? _GEN_686 : tag_2_14; // @[playground/src/noop/dcache.scala 250:46 88:26]
  wire [21:0] _GEN_816 = io_dataAxi_rd_bits_last ? _GEN_687 : tag_2_15; // @[playground/src/noop/dcache.scala 250:46 88:26]
  wire [21:0] _GEN_817 = io_dataAxi_rd_bits_last ? _GEN_688 : tag_3_0; // @[playground/src/noop/dcache.scala 250:46 88:26]
  wire [21:0] _GEN_818 = io_dataAxi_rd_bits_last ? _GEN_689 : tag_3_1; // @[playground/src/noop/dcache.scala 250:46 88:26]
  wire [21:0] _GEN_819 = io_dataAxi_rd_bits_last ? _GEN_690 : tag_3_2; // @[playground/src/noop/dcache.scala 250:46 88:26]
  wire [21:0] _GEN_820 = io_dataAxi_rd_bits_last ? _GEN_691 : tag_3_3; // @[playground/src/noop/dcache.scala 250:46 88:26]
  wire [21:0] _GEN_821 = io_dataAxi_rd_bits_last ? _GEN_692 : tag_3_4; // @[playground/src/noop/dcache.scala 250:46 88:26]
  wire [21:0] _GEN_822 = io_dataAxi_rd_bits_last ? _GEN_693 : tag_3_5; // @[playground/src/noop/dcache.scala 250:46 88:26]
  wire [21:0] _GEN_823 = io_dataAxi_rd_bits_last ? _GEN_694 : tag_3_6; // @[playground/src/noop/dcache.scala 250:46 88:26]
  wire [21:0] _GEN_824 = io_dataAxi_rd_bits_last ? _GEN_695 : tag_3_7; // @[playground/src/noop/dcache.scala 250:46 88:26]
  wire [21:0] _GEN_825 = io_dataAxi_rd_bits_last ? _GEN_696 : tag_3_8; // @[playground/src/noop/dcache.scala 250:46 88:26]
  wire [21:0] _GEN_826 = io_dataAxi_rd_bits_last ? _GEN_697 : tag_3_9; // @[playground/src/noop/dcache.scala 250:46 88:26]
  wire [21:0] _GEN_827 = io_dataAxi_rd_bits_last ? _GEN_698 : tag_3_10; // @[playground/src/noop/dcache.scala 250:46 88:26]
  wire [21:0] _GEN_828 = io_dataAxi_rd_bits_last ? _GEN_699 : tag_3_11; // @[playground/src/noop/dcache.scala 250:46 88:26]
  wire [21:0] _GEN_829 = io_dataAxi_rd_bits_last ? _GEN_700 : tag_3_12; // @[playground/src/noop/dcache.scala 250:46 88:26]
  wire [21:0] _GEN_830 = io_dataAxi_rd_bits_last ? _GEN_701 : tag_3_13; // @[playground/src/noop/dcache.scala 250:46 88:26]
  wire [21:0] _GEN_831 = io_dataAxi_rd_bits_last ? _GEN_702 : tag_3_14; // @[playground/src/noop/dcache.scala 250:46 88:26]
  wire [21:0] _GEN_832 = io_dataAxi_rd_bits_last ? _GEN_703 : tag_3_15; // @[playground/src/noop/dcache.scala 250:46 88:26]
  wire  _GEN_833 = io_dataAxi_rd_bits_last ? _GEN_704 : valid_0_0; // @[playground/src/noop/dcache.scala 250:46 89:26]
  wire  _GEN_834 = io_dataAxi_rd_bits_last ? _GEN_705 : valid_0_1; // @[playground/src/noop/dcache.scala 250:46 89:26]
  wire  _GEN_835 = io_dataAxi_rd_bits_last ? _GEN_706 : valid_0_2; // @[playground/src/noop/dcache.scala 250:46 89:26]
  wire  _GEN_836 = io_dataAxi_rd_bits_last ? _GEN_707 : valid_0_3; // @[playground/src/noop/dcache.scala 250:46 89:26]
  wire  _GEN_837 = io_dataAxi_rd_bits_last ? _GEN_708 : valid_0_4; // @[playground/src/noop/dcache.scala 250:46 89:26]
  wire  _GEN_838 = io_dataAxi_rd_bits_last ? _GEN_709 : valid_0_5; // @[playground/src/noop/dcache.scala 250:46 89:26]
  wire  _GEN_839 = io_dataAxi_rd_bits_last ? _GEN_710 : valid_0_6; // @[playground/src/noop/dcache.scala 250:46 89:26]
  wire  _GEN_840 = io_dataAxi_rd_bits_last ? _GEN_711 : valid_0_7; // @[playground/src/noop/dcache.scala 250:46 89:26]
  wire  _GEN_841 = io_dataAxi_rd_bits_last ? _GEN_712 : valid_0_8; // @[playground/src/noop/dcache.scala 250:46 89:26]
  wire  _GEN_842 = io_dataAxi_rd_bits_last ? _GEN_713 : valid_0_9; // @[playground/src/noop/dcache.scala 250:46 89:26]
  wire  _GEN_843 = io_dataAxi_rd_bits_last ? _GEN_714 : valid_0_10; // @[playground/src/noop/dcache.scala 250:46 89:26]
  wire  _GEN_844 = io_dataAxi_rd_bits_last ? _GEN_715 : valid_0_11; // @[playground/src/noop/dcache.scala 250:46 89:26]
  wire  _GEN_845 = io_dataAxi_rd_bits_last ? _GEN_716 : valid_0_12; // @[playground/src/noop/dcache.scala 250:46 89:26]
  wire  _GEN_846 = io_dataAxi_rd_bits_last ? _GEN_717 : valid_0_13; // @[playground/src/noop/dcache.scala 250:46 89:26]
  wire  _GEN_847 = io_dataAxi_rd_bits_last ? _GEN_718 : valid_0_14; // @[playground/src/noop/dcache.scala 250:46 89:26]
  wire  _GEN_848 = io_dataAxi_rd_bits_last ? _GEN_719 : valid_0_15; // @[playground/src/noop/dcache.scala 250:46 89:26]
  wire  _GEN_849 = io_dataAxi_rd_bits_last ? _GEN_720 : valid_1_0; // @[playground/src/noop/dcache.scala 250:46 89:26]
  wire  _GEN_850 = io_dataAxi_rd_bits_last ? _GEN_721 : valid_1_1; // @[playground/src/noop/dcache.scala 250:46 89:26]
  wire  _GEN_851 = io_dataAxi_rd_bits_last ? _GEN_722 : valid_1_2; // @[playground/src/noop/dcache.scala 250:46 89:26]
  wire  _GEN_852 = io_dataAxi_rd_bits_last ? _GEN_723 : valid_1_3; // @[playground/src/noop/dcache.scala 250:46 89:26]
  wire  _GEN_853 = io_dataAxi_rd_bits_last ? _GEN_724 : valid_1_4; // @[playground/src/noop/dcache.scala 250:46 89:26]
  wire  _GEN_854 = io_dataAxi_rd_bits_last ? _GEN_725 : valid_1_5; // @[playground/src/noop/dcache.scala 250:46 89:26]
  wire  _GEN_855 = io_dataAxi_rd_bits_last ? _GEN_726 : valid_1_6; // @[playground/src/noop/dcache.scala 250:46 89:26]
  wire  _GEN_856 = io_dataAxi_rd_bits_last ? _GEN_727 : valid_1_7; // @[playground/src/noop/dcache.scala 250:46 89:26]
  wire  _GEN_857 = io_dataAxi_rd_bits_last ? _GEN_728 : valid_1_8; // @[playground/src/noop/dcache.scala 250:46 89:26]
  wire  _GEN_858 = io_dataAxi_rd_bits_last ? _GEN_729 : valid_1_9; // @[playground/src/noop/dcache.scala 250:46 89:26]
  wire  _GEN_859 = io_dataAxi_rd_bits_last ? _GEN_730 : valid_1_10; // @[playground/src/noop/dcache.scala 250:46 89:26]
  wire  _GEN_860 = io_dataAxi_rd_bits_last ? _GEN_731 : valid_1_11; // @[playground/src/noop/dcache.scala 250:46 89:26]
  wire  _GEN_861 = io_dataAxi_rd_bits_last ? _GEN_732 : valid_1_12; // @[playground/src/noop/dcache.scala 250:46 89:26]
  wire  _GEN_862 = io_dataAxi_rd_bits_last ? _GEN_733 : valid_1_13; // @[playground/src/noop/dcache.scala 250:46 89:26]
  wire  _GEN_863 = io_dataAxi_rd_bits_last ? _GEN_734 : valid_1_14; // @[playground/src/noop/dcache.scala 250:46 89:26]
  wire  _GEN_864 = io_dataAxi_rd_bits_last ? _GEN_735 : valid_1_15; // @[playground/src/noop/dcache.scala 250:46 89:26]
  wire  _GEN_865 = io_dataAxi_rd_bits_last ? _GEN_736 : valid_2_0; // @[playground/src/noop/dcache.scala 250:46 89:26]
  wire  _GEN_866 = io_dataAxi_rd_bits_last ? _GEN_737 : valid_2_1; // @[playground/src/noop/dcache.scala 250:46 89:26]
  wire  _GEN_867 = io_dataAxi_rd_bits_last ? _GEN_738 : valid_2_2; // @[playground/src/noop/dcache.scala 250:46 89:26]
  wire  _GEN_868 = io_dataAxi_rd_bits_last ? _GEN_739 : valid_2_3; // @[playground/src/noop/dcache.scala 250:46 89:26]
  wire  _GEN_869 = io_dataAxi_rd_bits_last ? _GEN_740 : valid_2_4; // @[playground/src/noop/dcache.scala 250:46 89:26]
  wire  _GEN_870 = io_dataAxi_rd_bits_last ? _GEN_741 : valid_2_5; // @[playground/src/noop/dcache.scala 250:46 89:26]
  wire  _GEN_871 = io_dataAxi_rd_bits_last ? _GEN_742 : valid_2_6; // @[playground/src/noop/dcache.scala 250:46 89:26]
  wire  _GEN_872 = io_dataAxi_rd_bits_last ? _GEN_743 : valid_2_7; // @[playground/src/noop/dcache.scala 250:46 89:26]
  wire  _GEN_873 = io_dataAxi_rd_bits_last ? _GEN_744 : valid_2_8; // @[playground/src/noop/dcache.scala 250:46 89:26]
  wire  _GEN_874 = io_dataAxi_rd_bits_last ? _GEN_745 : valid_2_9; // @[playground/src/noop/dcache.scala 250:46 89:26]
  wire  _GEN_875 = io_dataAxi_rd_bits_last ? _GEN_746 : valid_2_10; // @[playground/src/noop/dcache.scala 250:46 89:26]
  wire  _GEN_876 = io_dataAxi_rd_bits_last ? _GEN_747 : valid_2_11; // @[playground/src/noop/dcache.scala 250:46 89:26]
  wire  _GEN_877 = io_dataAxi_rd_bits_last ? _GEN_748 : valid_2_12; // @[playground/src/noop/dcache.scala 250:46 89:26]
  wire  _GEN_878 = io_dataAxi_rd_bits_last ? _GEN_749 : valid_2_13; // @[playground/src/noop/dcache.scala 250:46 89:26]
  wire  _GEN_879 = io_dataAxi_rd_bits_last ? _GEN_750 : valid_2_14; // @[playground/src/noop/dcache.scala 250:46 89:26]
  wire  _GEN_880 = io_dataAxi_rd_bits_last ? _GEN_751 : valid_2_15; // @[playground/src/noop/dcache.scala 250:46 89:26]
  wire  _GEN_881 = io_dataAxi_rd_bits_last ? _GEN_752 : valid_3_0; // @[playground/src/noop/dcache.scala 250:46 89:26]
  wire  _GEN_882 = io_dataAxi_rd_bits_last ? _GEN_753 : valid_3_1; // @[playground/src/noop/dcache.scala 250:46 89:26]
  wire  _GEN_883 = io_dataAxi_rd_bits_last ? _GEN_754 : valid_3_2; // @[playground/src/noop/dcache.scala 250:46 89:26]
  wire  _GEN_884 = io_dataAxi_rd_bits_last ? _GEN_755 : valid_3_3; // @[playground/src/noop/dcache.scala 250:46 89:26]
  wire  _GEN_885 = io_dataAxi_rd_bits_last ? _GEN_756 : valid_3_4; // @[playground/src/noop/dcache.scala 250:46 89:26]
  wire  _GEN_886 = io_dataAxi_rd_bits_last ? _GEN_757 : valid_3_5; // @[playground/src/noop/dcache.scala 250:46 89:26]
  wire  _GEN_887 = io_dataAxi_rd_bits_last ? _GEN_758 : valid_3_6; // @[playground/src/noop/dcache.scala 250:46 89:26]
  wire  _GEN_888 = io_dataAxi_rd_bits_last ? _GEN_759 : valid_3_7; // @[playground/src/noop/dcache.scala 250:46 89:26]
  wire  _GEN_889 = io_dataAxi_rd_bits_last ? _GEN_760 : valid_3_8; // @[playground/src/noop/dcache.scala 250:46 89:26]
  wire  _GEN_890 = io_dataAxi_rd_bits_last ? _GEN_761 : valid_3_9; // @[playground/src/noop/dcache.scala 250:46 89:26]
  wire  _GEN_891 = io_dataAxi_rd_bits_last ? _GEN_762 : valid_3_10; // @[playground/src/noop/dcache.scala 250:46 89:26]
  wire  _GEN_892 = io_dataAxi_rd_bits_last ? _GEN_763 : valid_3_11; // @[playground/src/noop/dcache.scala 250:46 89:26]
  wire  _GEN_893 = io_dataAxi_rd_bits_last ? _GEN_764 : valid_3_12; // @[playground/src/noop/dcache.scala 250:46 89:26]
  wire  _GEN_894 = io_dataAxi_rd_bits_last ? _GEN_765 : valid_3_13; // @[playground/src/noop/dcache.scala 250:46 89:26]
  wire  _GEN_895 = io_dataAxi_rd_bits_last ? _GEN_766 : valid_3_14; // @[playground/src/noop/dcache.scala 250:46 89:26]
  wire  _GEN_896 = io_dataAxi_rd_bits_last ? _GEN_767 : valid_3_15; // @[playground/src/noop/dcache.scala 250:46 89:26]
  wire [2:0] _GEN_897 = io_dataAxi_rd_bits_last ? 3'h0 : state; // @[playground/src/noop/dcache.scala 152:24 250:46 254:27]
  wire [2:0] _GEN_898 = axiRdataEn & io_dataAxi_rd_valid ? _offset_T_1 : offset; // @[playground/src/noop/dcache.scala 243:52 244:24 110:34]
  wire [63:0] _GEN_900 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_639 : rdatabuf; // @[playground/src/noop/dcache.scala 111:34 243:52]
  wire  _GEN_901 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_768 : axiRdataEn; // @[playground/src/noop/dcache.scala 198:34 243:52]
  wire [21:0] _GEN_902 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_769 : tag_0_0; // @[playground/src/noop/dcache.scala 243:52 88:26]
  wire [21:0] _GEN_903 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_770 : tag_0_1; // @[playground/src/noop/dcache.scala 243:52 88:26]
  wire [21:0] _GEN_904 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_771 : tag_0_2; // @[playground/src/noop/dcache.scala 243:52 88:26]
  wire [21:0] _GEN_905 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_772 : tag_0_3; // @[playground/src/noop/dcache.scala 243:52 88:26]
  wire [21:0] _GEN_906 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_773 : tag_0_4; // @[playground/src/noop/dcache.scala 243:52 88:26]
  wire [21:0] _GEN_907 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_774 : tag_0_5; // @[playground/src/noop/dcache.scala 243:52 88:26]
  wire [21:0] _GEN_908 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_775 : tag_0_6; // @[playground/src/noop/dcache.scala 243:52 88:26]
  wire [21:0] _GEN_909 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_776 : tag_0_7; // @[playground/src/noop/dcache.scala 243:52 88:26]
  wire [21:0] _GEN_910 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_777 : tag_0_8; // @[playground/src/noop/dcache.scala 243:52 88:26]
  wire [21:0] _GEN_911 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_778 : tag_0_9; // @[playground/src/noop/dcache.scala 243:52 88:26]
  wire [21:0] _GEN_912 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_779 : tag_0_10; // @[playground/src/noop/dcache.scala 243:52 88:26]
  wire [21:0] _GEN_913 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_780 : tag_0_11; // @[playground/src/noop/dcache.scala 243:52 88:26]
  wire [21:0] _GEN_914 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_781 : tag_0_12; // @[playground/src/noop/dcache.scala 243:52 88:26]
  wire [21:0] _GEN_915 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_782 : tag_0_13; // @[playground/src/noop/dcache.scala 243:52 88:26]
  wire [21:0] _GEN_916 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_783 : tag_0_14; // @[playground/src/noop/dcache.scala 243:52 88:26]
  wire [21:0] _GEN_917 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_784 : tag_0_15; // @[playground/src/noop/dcache.scala 243:52 88:26]
  wire [21:0] _GEN_918 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_785 : tag_1_0; // @[playground/src/noop/dcache.scala 243:52 88:26]
  wire [21:0] _GEN_919 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_786 : tag_1_1; // @[playground/src/noop/dcache.scala 243:52 88:26]
  wire [21:0] _GEN_920 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_787 : tag_1_2; // @[playground/src/noop/dcache.scala 243:52 88:26]
  wire [21:0] _GEN_921 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_788 : tag_1_3; // @[playground/src/noop/dcache.scala 243:52 88:26]
  wire [21:0] _GEN_922 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_789 : tag_1_4; // @[playground/src/noop/dcache.scala 243:52 88:26]
  wire [21:0] _GEN_923 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_790 : tag_1_5; // @[playground/src/noop/dcache.scala 243:52 88:26]
  wire [21:0] _GEN_924 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_791 : tag_1_6; // @[playground/src/noop/dcache.scala 243:52 88:26]
  wire [21:0] _GEN_925 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_792 : tag_1_7; // @[playground/src/noop/dcache.scala 243:52 88:26]
  wire [21:0] _GEN_926 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_793 : tag_1_8; // @[playground/src/noop/dcache.scala 243:52 88:26]
  wire [21:0] _GEN_927 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_794 : tag_1_9; // @[playground/src/noop/dcache.scala 243:52 88:26]
  wire [21:0] _GEN_928 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_795 : tag_1_10; // @[playground/src/noop/dcache.scala 243:52 88:26]
  wire [21:0] _GEN_929 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_796 : tag_1_11; // @[playground/src/noop/dcache.scala 243:52 88:26]
  wire [21:0] _GEN_930 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_797 : tag_1_12; // @[playground/src/noop/dcache.scala 243:52 88:26]
  wire [21:0] _GEN_931 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_798 : tag_1_13; // @[playground/src/noop/dcache.scala 243:52 88:26]
  wire [21:0] _GEN_932 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_799 : tag_1_14; // @[playground/src/noop/dcache.scala 243:52 88:26]
  wire [21:0] _GEN_933 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_800 : tag_1_15; // @[playground/src/noop/dcache.scala 243:52 88:26]
  wire [21:0] _GEN_934 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_801 : tag_2_0; // @[playground/src/noop/dcache.scala 243:52 88:26]
  wire [21:0] _GEN_935 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_802 : tag_2_1; // @[playground/src/noop/dcache.scala 243:52 88:26]
  wire [21:0] _GEN_936 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_803 : tag_2_2; // @[playground/src/noop/dcache.scala 243:52 88:26]
  wire [21:0] _GEN_937 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_804 : tag_2_3; // @[playground/src/noop/dcache.scala 243:52 88:26]
  wire [21:0] _GEN_938 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_805 : tag_2_4; // @[playground/src/noop/dcache.scala 243:52 88:26]
  wire [21:0] _GEN_939 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_806 : tag_2_5; // @[playground/src/noop/dcache.scala 243:52 88:26]
  wire [21:0] _GEN_940 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_807 : tag_2_6; // @[playground/src/noop/dcache.scala 243:52 88:26]
  wire [21:0] _GEN_941 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_808 : tag_2_7; // @[playground/src/noop/dcache.scala 243:52 88:26]
  wire [21:0] _GEN_942 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_809 : tag_2_8; // @[playground/src/noop/dcache.scala 243:52 88:26]
  wire [21:0] _GEN_943 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_810 : tag_2_9; // @[playground/src/noop/dcache.scala 243:52 88:26]
  wire [21:0] _GEN_944 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_811 : tag_2_10; // @[playground/src/noop/dcache.scala 243:52 88:26]
  wire [21:0] _GEN_945 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_812 : tag_2_11; // @[playground/src/noop/dcache.scala 243:52 88:26]
  wire [21:0] _GEN_946 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_813 : tag_2_12; // @[playground/src/noop/dcache.scala 243:52 88:26]
  wire [21:0] _GEN_947 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_814 : tag_2_13; // @[playground/src/noop/dcache.scala 243:52 88:26]
  wire [21:0] _GEN_948 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_815 : tag_2_14; // @[playground/src/noop/dcache.scala 243:52 88:26]
  wire [21:0] _GEN_949 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_816 : tag_2_15; // @[playground/src/noop/dcache.scala 243:52 88:26]
  wire [21:0] _GEN_950 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_817 : tag_3_0; // @[playground/src/noop/dcache.scala 243:52 88:26]
  wire [21:0] _GEN_951 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_818 : tag_3_1; // @[playground/src/noop/dcache.scala 243:52 88:26]
  wire [21:0] _GEN_952 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_819 : tag_3_2; // @[playground/src/noop/dcache.scala 243:52 88:26]
  wire [21:0] _GEN_953 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_820 : tag_3_3; // @[playground/src/noop/dcache.scala 243:52 88:26]
  wire [21:0] _GEN_954 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_821 : tag_3_4; // @[playground/src/noop/dcache.scala 243:52 88:26]
  wire [21:0] _GEN_955 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_822 : tag_3_5; // @[playground/src/noop/dcache.scala 243:52 88:26]
  wire [21:0] _GEN_956 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_823 : tag_3_6; // @[playground/src/noop/dcache.scala 243:52 88:26]
  wire [21:0] _GEN_957 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_824 : tag_3_7; // @[playground/src/noop/dcache.scala 243:52 88:26]
  wire [21:0] _GEN_958 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_825 : tag_3_8; // @[playground/src/noop/dcache.scala 243:52 88:26]
  wire [21:0] _GEN_959 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_826 : tag_3_9; // @[playground/src/noop/dcache.scala 243:52 88:26]
  wire [21:0] _GEN_960 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_827 : tag_3_10; // @[playground/src/noop/dcache.scala 243:52 88:26]
  wire [21:0] _GEN_961 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_828 : tag_3_11; // @[playground/src/noop/dcache.scala 243:52 88:26]
  wire [21:0] _GEN_962 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_829 : tag_3_12; // @[playground/src/noop/dcache.scala 243:52 88:26]
  wire [21:0] _GEN_963 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_830 : tag_3_13; // @[playground/src/noop/dcache.scala 243:52 88:26]
  wire [21:0] _GEN_964 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_831 : tag_3_14; // @[playground/src/noop/dcache.scala 243:52 88:26]
  wire [21:0] _GEN_965 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_832 : tag_3_15; // @[playground/src/noop/dcache.scala 243:52 88:26]
  wire  _GEN_966 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_833 : valid_0_0; // @[playground/src/noop/dcache.scala 243:52 89:26]
  wire  _GEN_967 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_834 : valid_0_1; // @[playground/src/noop/dcache.scala 243:52 89:26]
  wire  _GEN_968 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_835 : valid_0_2; // @[playground/src/noop/dcache.scala 243:52 89:26]
  wire  _GEN_969 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_836 : valid_0_3; // @[playground/src/noop/dcache.scala 243:52 89:26]
  wire  _GEN_970 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_837 : valid_0_4; // @[playground/src/noop/dcache.scala 243:52 89:26]
  wire  _GEN_971 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_838 : valid_0_5; // @[playground/src/noop/dcache.scala 243:52 89:26]
  wire  _GEN_972 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_839 : valid_0_6; // @[playground/src/noop/dcache.scala 243:52 89:26]
  wire  _GEN_973 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_840 : valid_0_7; // @[playground/src/noop/dcache.scala 243:52 89:26]
  wire  _GEN_974 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_841 : valid_0_8; // @[playground/src/noop/dcache.scala 243:52 89:26]
  wire  _GEN_975 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_842 : valid_0_9; // @[playground/src/noop/dcache.scala 243:52 89:26]
  wire  _GEN_976 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_843 : valid_0_10; // @[playground/src/noop/dcache.scala 243:52 89:26]
  wire  _GEN_977 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_844 : valid_0_11; // @[playground/src/noop/dcache.scala 243:52 89:26]
  wire  _GEN_978 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_845 : valid_0_12; // @[playground/src/noop/dcache.scala 243:52 89:26]
  wire  _GEN_979 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_846 : valid_0_13; // @[playground/src/noop/dcache.scala 243:52 89:26]
  wire  _GEN_980 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_847 : valid_0_14; // @[playground/src/noop/dcache.scala 243:52 89:26]
  wire  _GEN_981 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_848 : valid_0_15; // @[playground/src/noop/dcache.scala 243:52 89:26]
  wire  _GEN_982 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_849 : valid_1_0; // @[playground/src/noop/dcache.scala 243:52 89:26]
  wire  _GEN_983 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_850 : valid_1_1; // @[playground/src/noop/dcache.scala 243:52 89:26]
  wire  _GEN_984 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_851 : valid_1_2; // @[playground/src/noop/dcache.scala 243:52 89:26]
  wire  _GEN_985 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_852 : valid_1_3; // @[playground/src/noop/dcache.scala 243:52 89:26]
  wire  _GEN_986 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_853 : valid_1_4; // @[playground/src/noop/dcache.scala 243:52 89:26]
  wire  _GEN_987 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_854 : valid_1_5; // @[playground/src/noop/dcache.scala 243:52 89:26]
  wire  _GEN_988 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_855 : valid_1_6; // @[playground/src/noop/dcache.scala 243:52 89:26]
  wire  _GEN_989 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_856 : valid_1_7; // @[playground/src/noop/dcache.scala 243:52 89:26]
  wire  _GEN_990 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_857 : valid_1_8; // @[playground/src/noop/dcache.scala 243:52 89:26]
  wire  _GEN_991 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_858 : valid_1_9; // @[playground/src/noop/dcache.scala 243:52 89:26]
  wire  _GEN_992 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_859 : valid_1_10; // @[playground/src/noop/dcache.scala 243:52 89:26]
  wire  _GEN_993 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_860 : valid_1_11; // @[playground/src/noop/dcache.scala 243:52 89:26]
  wire  _GEN_994 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_861 : valid_1_12; // @[playground/src/noop/dcache.scala 243:52 89:26]
  wire  _GEN_995 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_862 : valid_1_13; // @[playground/src/noop/dcache.scala 243:52 89:26]
  wire  _GEN_996 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_863 : valid_1_14; // @[playground/src/noop/dcache.scala 243:52 89:26]
  wire  _GEN_997 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_864 : valid_1_15; // @[playground/src/noop/dcache.scala 243:52 89:26]
  wire  _GEN_998 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_865 : valid_2_0; // @[playground/src/noop/dcache.scala 243:52 89:26]
  wire  _GEN_999 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_866 : valid_2_1; // @[playground/src/noop/dcache.scala 243:52 89:26]
  wire  _GEN_1000 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_867 : valid_2_2; // @[playground/src/noop/dcache.scala 243:52 89:26]
  wire  _GEN_1001 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_868 : valid_2_3; // @[playground/src/noop/dcache.scala 243:52 89:26]
  wire  _GEN_1002 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_869 : valid_2_4; // @[playground/src/noop/dcache.scala 243:52 89:26]
  wire  _GEN_1003 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_870 : valid_2_5; // @[playground/src/noop/dcache.scala 243:52 89:26]
  wire  _GEN_1004 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_871 : valid_2_6; // @[playground/src/noop/dcache.scala 243:52 89:26]
  wire  _GEN_1005 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_872 : valid_2_7; // @[playground/src/noop/dcache.scala 243:52 89:26]
  wire  _GEN_1006 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_873 : valid_2_8; // @[playground/src/noop/dcache.scala 243:52 89:26]
  wire  _GEN_1007 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_874 : valid_2_9; // @[playground/src/noop/dcache.scala 243:52 89:26]
  wire  _GEN_1008 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_875 : valid_2_10; // @[playground/src/noop/dcache.scala 243:52 89:26]
  wire  _GEN_1009 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_876 : valid_2_11; // @[playground/src/noop/dcache.scala 243:52 89:26]
  wire  _GEN_1010 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_877 : valid_2_12; // @[playground/src/noop/dcache.scala 243:52 89:26]
  wire  _GEN_1011 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_878 : valid_2_13; // @[playground/src/noop/dcache.scala 243:52 89:26]
  wire  _GEN_1012 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_879 : valid_2_14; // @[playground/src/noop/dcache.scala 243:52 89:26]
  wire  _GEN_1013 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_880 : valid_2_15; // @[playground/src/noop/dcache.scala 243:52 89:26]
  wire  _GEN_1014 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_881 : valid_3_0; // @[playground/src/noop/dcache.scala 243:52 89:26]
  wire  _GEN_1015 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_882 : valid_3_1; // @[playground/src/noop/dcache.scala 243:52 89:26]
  wire  _GEN_1016 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_883 : valid_3_2; // @[playground/src/noop/dcache.scala 243:52 89:26]
  wire  _GEN_1017 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_884 : valid_3_3; // @[playground/src/noop/dcache.scala 243:52 89:26]
  wire  _GEN_1018 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_885 : valid_3_4; // @[playground/src/noop/dcache.scala 243:52 89:26]
  wire  _GEN_1019 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_886 : valid_3_5; // @[playground/src/noop/dcache.scala 243:52 89:26]
  wire  _GEN_1020 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_887 : valid_3_6; // @[playground/src/noop/dcache.scala 243:52 89:26]
  wire  _GEN_1021 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_888 : valid_3_7; // @[playground/src/noop/dcache.scala 243:52 89:26]
  wire  _GEN_1022 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_889 : valid_3_8; // @[playground/src/noop/dcache.scala 243:52 89:26]
  wire  _GEN_1023 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_890 : valid_3_9; // @[playground/src/noop/dcache.scala 243:52 89:26]
  wire  _GEN_1024 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_891 : valid_3_10; // @[playground/src/noop/dcache.scala 243:52 89:26]
  wire  _GEN_1025 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_892 : valid_3_11; // @[playground/src/noop/dcache.scala 243:52 89:26]
  wire  _GEN_1026 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_893 : valid_3_12; // @[playground/src/noop/dcache.scala 243:52 89:26]
  wire  _GEN_1027 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_894 : valid_3_13; // @[playground/src/noop/dcache.scala 243:52 89:26]
  wire  _GEN_1028 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_895 : valid_3_14; // @[playground/src/noop/dcache.scala 243:52 89:26]
  wire  _GEN_1029 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_896 : valid_3_15; // @[playground/src/noop/dcache.scala 243:52 89:26]
  wire [2:0] _GEN_1030 = axiRdataEn & io_dataAxi_rd_valid ? _GEN_897 : state; // @[playground/src/noop/dcache.scala 152:24 243:52]
  wire [2:0] _GEN_1031 = axiWaddrEn & io_dataAxi_wa_ready ? 3'h4 : state; // @[playground/src/noop/dcache.scala 152:24 260:52 261:29]
  wire  _GEN_1032 = axiWaddrEn & io_dataAxi_wa_ready ? 1'h0 : axiWaddrEn; // @[playground/src/noop/dcache.scala 260:52 262:29 199:34]
  wire  _GEN_1033 = axiWaddrEn & io_dataAxi_wa_ready | axiWdataEn; // @[playground/src/noop/dcache.scala 260:52 263:29 202:34]
  wire  _GEN_1034 = _GEN_2724 & _GEN_2755 ? 1'h0 : valid_0_0; // @[playground/src/noop/dcache.scala 274:{51,51} 89:26]
  wire  _GEN_1035 = _GEN_2724 & _GEN_2725 ? 1'h0 : valid_0_1; // @[playground/src/noop/dcache.scala 274:{51,51} 89:26]
  wire  _GEN_1036 = _GEN_2724 & _GEN_2727 ? 1'h0 : valid_0_2; // @[playground/src/noop/dcache.scala 274:{51,51} 89:26]
  wire  _GEN_1037 = _GEN_2724 & _GEN_2729 ? 1'h0 : valid_0_3; // @[playground/src/noop/dcache.scala 274:{51,51} 89:26]
  wire  _GEN_1038 = _GEN_2724 & _GEN_2731 ? 1'h0 : valid_0_4; // @[playground/src/noop/dcache.scala 274:{51,51} 89:26]
  wire  _GEN_1039 = _GEN_2724 & _GEN_2733 ? 1'h0 : valid_0_5; // @[playground/src/noop/dcache.scala 274:{51,51} 89:26]
  wire  _GEN_1040 = _GEN_2724 & _GEN_2735 ? 1'h0 : valid_0_6; // @[playground/src/noop/dcache.scala 274:{51,51} 89:26]
  wire  _GEN_1041 = _GEN_2724 & _GEN_2737 ? 1'h0 : valid_0_7; // @[playground/src/noop/dcache.scala 274:{51,51} 89:26]
  wire  _GEN_1042 = _GEN_2724 & _GEN_2739 ? 1'h0 : valid_0_8; // @[playground/src/noop/dcache.scala 274:{51,51} 89:26]
  wire  _GEN_1043 = _GEN_2724 & _GEN_2741 ? 1'h0 : valid_0_9; // @[playground/src/noop/dcache.scala 274:{51,51} 89:26]
  wire  _GEN_1044 = _GEN_2724 & _GEN_2743 ? 1'h0 : valid_0_10; // @[playground/src/noop/dcache.scala 274:{51,51} 89:26]
  wire  _GEN_1045 = _GEN_2724 & _GEN_2745 ? 1'h0 : valid_0_11; // @[playground/src/noop/dcache.scala 274:{51,51} 89:26]
  wire  _GEN_1046 = _GEN_2724 & _GEN_2747 ? 1'h0 : valid_0_12; // @[playground/src/noop/dcache.scala 274:{51,51} 89:26]
  wire  _GEN_1047 = _GEN_2724 & _GEN_2749 ? 1'h0 : valid_0_13; // @[playground/src/noop/dcache.scala 274:{51,51} 89:26]
  wire  _GEN_1048 = _GEN_2724 & _GEN_2751 ? 1'h0 : valid_0_14; // @[playground/src/noop/dcache.scala 274:{51,51} 89:26]
  wire  _GEN_1049 = _GEN_2724 & _GEN_2753 ? 1'h0 : valid_0_15; // @[playground/src/noop/dcache.scala 274:{51,51} 89:26]
  wire  _GEN_1050 = _GEN_2754 & _GEN_2755 ? 1'h0 : valid_1_0; // @[playground/src/noop/dcache.scala 274:{51,51} 89:26]
  wire  _GEN_1051 = _GEN_2754 & _GEN_2725 ? 1'h0 : valid_1_1; // @[playground/src/noop/dcache.scala 274:{51,51} 89:26]
  wire  _GEN_1052 = _GEN_2754 & _GEN_2727 ? 1'h0 : valid_1_2; // @[playground/src/noop/dcache.scala 274:{51,51} 89:26]
  wire  _GEN_1053 = _GEN_2754 & _GEN_2729 ? 1'h0 : valid_1_3; // @[playground/src/noop/dcache.scala 274:{51,51} 89:26]
  wire  _GEN_1054 = _GEN_2754 & _GEN_2731 ? 1'h0 : valid_1_4; // @[playground/src/noop/dcache.scala 274:{51,51} 89:26]
  wire  _GEN_1055 = _GEN_2754 & _GEN_2733 ? 1'h0 : valid_1_5; // @[playground/src/noop/dcache.scala 274:{51,51} 89:26]
  wire  _GEN_1056 = _GEN_2754 & _GEN_2735 ? 1'h0 : valid_1_6; // @[playground/src/noop/dcache.scala 274:{51,51} 89:26]
  wire  _GEN_1057 = _GEN_2754 & _GEN_2737 ? 1'h0 : valid_1_7; // @[playground/src/noop/dcache.scala 274:{51,51} 89:26]
  wire  _GEN_1058 = _GEN_2754 & _GEN_2739 ? 1'h0 : valid_1_8; // @[playground/src/noop/dcache.scala 274:{51,51} 89:26]
  wire  _GEN_1059 = _GEN_2754 & _GEN_2741 ? 1'h0 : valid_1_9; // @[playground/src/noop/dcache.scala 274:{51,51} 89:26]
  wire  _GEN_1060 = _GEN_2754 & _GEN_2743 ? 1'h0 : valid_1_10; // @[playground/src/noop/dcache.scala 274:{51,51} 89:26]
  wire  _GEN_1061 = _GEN_2754 & _GEN_2745 ? 1'h0 : valid_1_11; // @[playground/src/noop/dcache.scala 274:{51,51} 89:26]
  wire  _GEN_1062 = _GEN_2754 & _GEN_2747 ? 1'h0 : valid_1_12; // @[playground/src/noop/dcache.scala 274:{51,51} 89:26]
  wire  _GEN_1063 = _GEN_2754 & _GEN_2749 ? 1'h0 : valid_1_13; // @[playground/src/noop/dcache.scala 274:{51,51} 89:26]
  wire  _GEN_1064 = _GEN_2754 & _GEN_2751 ? 1'h0 : valid_1_14; // @[playground/src/noop/dcache.scala 274:{51,51} 89:26]
  wire  _GEN_1065 = _GEN_2754 & _GEN_2753 ? 1'h0 : valid_1_15; // @[playground/src/noop/dcache.scala 274:{51,51} 89:26]
  wire  _GEN_1066 = _GEN_2786 & _GEN_2755 ? 1'h0 : valid_2_0; // @[playground/src/noop/dcache.scala 274:{51,51} 89:26]
  wire  _GEN_1067 = _GEN_2786 & _GEN_2725 ? 1'h0 : valid_2_1; // @[playground/src/noop/dcache.scala 274:{51,51} 89:26]
  wire  _GEN_1068 = _GEN_2786 & _GEN_2727 ? 1'h0 : valid_2_2; // @[playground/src/noop/dcache.scala 274:{51,51} 89:26]
  wire  _GEN_1069 = _GEN_2786 & _GEN_2729 ? 1'h0 : valid_2_3; // @[playground/src/noop/dcache.scala 274:{51,51} 89:26]
  wire  _GEN_1070 = _GEN_2786 & _GEN_2731 ? 1'h0 : valid_2_4; // @[playground/src/noop/dcache.scala 274:{51,51} 89:26]
  wire  _GEN_1071 = _GEN_2786 & _GEN_2733 ? 1'h0 : valid_2_5; // @[playground/src/noop/dcache.scala 274:{51,51} 89:26]
  wire  _GEN_1072 = _GEN_2786 & _GEN_2735 ? 1'h0 : valid_2_6; // @[playground/src/noop/dcache.scala 274:{51,51} 89:26]
  wire  _GEN_1073 = _GEN_2786 & _GEN_2737 ? 1'h0 : valid_2_7; // @[playground/src/noop/dcache.scala 274:{51,51} 89:26]
  wire  _GEN_1074 = _GEN_2786 & _GEN_2739 ? 1'h0 : valid_2_8; // @[playground/src/noop/dcache.scala 274:{51,51} 89:26]
  wire  _GEN_1075 = _GEN_2786 & _GEN_2741 ? 1'h0 : valid_2_9; // @[playground/src/noop/dcache.scala 274:{51,51} 89:26]
  wire  _GEN_1076 = _GEN_2786 & _GEN_2743 ? 1'h0 : valid_2_10; // @[playground/src/noop/dcache.scala 274:{51,51} 89:26]
  wire  _GEN_1077 = _GEN_2786 & _GEN_2745 ? 1'h0 : valid_2_11; // @[playground/src/noop/dcache.scala 274:{51,51} 89:26]
  wire  _GEN_1078 = _GEN_2786 & _GEN_2747 ? 1'h0 : valid_2_12; // @[playground/src/noop/dcache.scala 274:{51,51} 89:26]
  wire  _GEN_1079 = _GEN_2786 & _GEN_2749 ? 1'h0 : valid_2_13; // @[playground/src/noop/dcache.scala 274:{51,51} 89:26]
  wire  _GEN_1080 = _GEN_2786 & _GEN_2751 ? 1'h0 : valid_2_14; // @[playground/src/noop/dcache.scala 274:{51,51} 89:26]
  wire  _GEN_1081 = _GEN_2786 & _GEN_2753 ? 1'h0 : valid_2_15; // @[playground/src/noop/dcache.scala 274:{51,51} 89:26]
  wire  _GEN_1082 = _GEN_2818 & _GEN_2755 ? 1'h0 : valid_3_0; // @[playground/src/noop/dcache.scala 274:{51,51} 89:26]
  wire  _GEN_1083 = _GEN_2818 & _GEN_2725 ? 1'h0 : valid_3_1; // @[playground/src/noop/dcache.scala 274:{51,51} 89:26]
  wire  _GEN_1084 = _GEN_2818 & _GEN_2727 ? 1'h0 : valid_3_2; // @[playground/src/noop/dcache.scala 274:{51,51} 89:26]
  wire  _GEN_1085 = _GEN_2818 & _GEN_2729 ? 1'h0 : valid_3_3; // @[playground/src/noop/dcache.scala 274:{51,51} 89:26]
  wire  _GEN_1086 = _GEN_2818 & _GEN_2731 ? 1'h0 : valid_3_4; // @[playground/src/noop/dcache.scala 274:{51,51} 89:26]
  wire  _GEN_1087 = _GEN_2818 & _GEN_2733 ? 1'h0 : valid_3_5; // @[playground/src/noop/dcache.scala 274:{51,51} 89:26]
  wire  _GEN_1088 = _GEN_2818 & _GEN_2735 ? 1'h0 : valid_3_6; // @[playground/src/noop/dcache.scala 274:{51,51} 89:26]
  wire  _GEN_1089 = _GEN_2818 & _GEN_2737 ? 1'h0 : valid_3_7; // @[playground/src/noop/dcache.scala 274:{51,51} 89:26]
  wire  _GEN_1090 = _GEN_2818 & _GEN_2739 ? 1'h0 : valid_3_8; // @[playground/src/noop/dcache.scala 274:{51,51} 89:26]
  wire  _GEN_1091 = _GEN_2818 & _GEN_2741 ? 1'h0 : valid_3_9; // @[playground/src/noop/dcache.scala 274:{51,51} 89:26]
  wire  _GEN_1092 = _GEN_2818 & _GEN_2743 ? 1'h0 : valid_3_10; // @[playground/src/noop/dcache.scala 274:{51,51} 89:26]
  wire  _GEN_1093 = _GEN_2818 & _GEN_2745 ? 1'h0 : valid_3_11; // @[playground/src/noop/dcache.scala 274:{51,51} 89:26]
  wire  _GEN_1094 = _GEN_2818 & _GEN_2747 ? 1'h0 : valid_3_12; // @[playground/src/noop/dcache.scala 274:{51,51} 89:26]
  wire  _GEN_1095 = _GEN_2818 & _GEN_2749 ? 1'h0 : valid_3_13; // @[playground/src/noop/dcache.scala 274:{51,51} 89:26]
  wire  _GEN_1096 = _GEN_2818 & _GEN_2751 ? 1'h0 : valid_3_14; // @[playground/src/noop/dcache.scala 274:{51,51} 89:26]
  wire  _GEN_1097 = _GEN_2818 & _GEN_2753 ? 1'h0 : valid_3_15; // @[playground/src/noop/dcache.scala 274:{51,51} 89:26]
  wire  _GEN_1098 = _GEN_2724 & _GEN_2755 ? 1'h0 : _GEN_414; // @[playground/src/noop/dcache.scala 275:{51,51}]
  wire  _GEN_1099 = _GEN_2724 & _GEN_2725 ? 1'h0 : _GEN_415; // @[playground/src/noop/dcache.scala 275:{51,51}]
  wire  _GEN_1100 = _GEN_2724 & _GEN_2727 ? 1'h0 : _GEN_416; // @[playground/src/noop/dcache.scala 275:{51,51}]
  wire  _GEN_1101 = _GEN_2724 & _GEN_2729 ? 1'h0 : _GEN_417; // @[playground/src/noop/dcache.scala 275:{51,51}]
  wire  _GEN_1102 = _GEN_2724 & _GEN_2731 ? 1'h0 : _GEN_418; // @[playground/src/noop/dcache.scala 275:{51,51}]
  wire  _GEN_1103 = _GEN_2724 & _GEN_2733 ? 1'h0 : _GEN_419; // @[playground/src/noop/dcache.scala 275:{51,51}]
  wire  _GEN_1104 = _GEN_2724 & _GEN_2735 ? 1'h0 : _GEN_420; // @[playground/src/noop/dcache.scala 275:{51,51}]
  wire  _GEN_1105 = _GEN_2724 & _GEN_2737 ? 1'h0 : _GEN_421; // @[playground/src/noop/dcache.scala 275:{51,51}]
  wire  _GEN_1106 = _GEN_2724 & _GEN_2739 ? 1'h0 : _GEN_422; // @[playground/src/noop/dcache.scala 275:{51,51}]
  wire  _GEN_1107 = _GEN_2724 & _GEN_2741 ? 1'h0 : _GEN_423; // @[playground/src/noop/dcache.scala 275:{51,51}]
  wire  _GEN_1108 = _GEN_2724 & _GEN_2743 ? 1'h0 : _GEN_424; // @[playground/src/noop/dcache.scala 275:{51,51}]
  wire  _GEN_1109 = _GEN_2724 & _GEN_2745 ? 1'h0 : _GEN_425; // @[playground/src/noop/dcache.scala 275:{51,51}]
  wire  _GEN_1110 = _GEN_2724 & _GEN_2747 ? 1'h0 : _GEN_426; // @[playground/src/noop/dcache.scala 275:{51,51}]
  wire  _GEN_1111 = _GEN_2724 & _GEN_2749 ? 1'h0 : _GEN_427; // @[playground/src/noop/dcache.scala 275:{51,51}]
  wire  _GEN_1112 = _GEN_2724 & _GEN_2751 ? 1'h0 : _GEN_428; // @[playground/src/noop/dcache.scala 275:{51,51}]
  wire  _GEN_1113 = _GEN_2724 & _GEN_2753 ? 1'h0 : _GEN_429; // @[playground/src/noop/dcache.scala 275:{51,51}]
  wire  _GEN_1114 = _GEN_2754 & _GEN_2755 ? 1'h0 : _GEN_430; // @[playground/src/noop/dcache.scala 275:{51,51}]
  wire  _GEN_1115 = _GEN_2754 & _GEN_2725 ? 1'h0 : _GEN_431; // @[playground/src/noop/dcache.scala 275:{51,51}]
  wire  _GEN_1116 = _GEN_2754 & _GEN_2727 ? 1'h0 : _GEN_432; // @[playground/src/noop/dcache.scala 275:{51,51}]
  wire  _GEN_1117 = _GEN_2754 & _GEN_2729 ? 1'h0 : _GEN_433; // @[playground/src/noop/dcache.scala 275:{51,51}]
  wire  _GEN_1118 = _GEN_2754 & _GEN_2731 ? 1'h0 : _GEN_434; // @[playground/src/noop/dcache.scala 275:{51,51}]
  wire  _GEN_1119 = _GEN_2754 & _GEN_2733 ? 1'h0 : _GEN_435; // @[playground/src/noop/dcache.scala 275:{51,51}]
  wire  _GEN_1120 = _GEN_2754 & _GEN_2735 ? 1'h0 : _GEN_436; // @[playground/src/noop/dcache.scala 275:{51,51}]
  wire  _GEN_1121 = _GEN_2754 & _GEN_2737 ? 1'h0 : _GEN_437; // @[playground/src/noop/dcache.scala 275:{51,51}]
  wire  _GEN_1122 = _GEN_2754 & _GEN_2739 ? 1'h0 : _GEN_438; // @[playground/src/noop/dcache.scala 275:{51,51}]
  wire  _GEN_1123 = _GEN_2754 & _GEN_2741 ? 1'h0 : _GEN_439; // @[playground/src/noop/dcache.scala 275:{51,51}]
  wire  _GEN_1124 = _GEN_2754 & _GEN_2743 ? 1'h0 : _GEN_440; // @[playground/src/noop/dcache.scala 275:{51,51}]
  wire  _GEN_1125 = _GEN_2754 & _GEN_2745 ? 1'h0 : _GEN_441; // @[playground/src/noop/dcache.scala 275:{51,51}]
  wire  _GEN_1126 = _GEN_2754 & _GEN_2747 ? 1'h0 : _GEN_442; // @[playground/src/noop/dcache.scala 275:{51,51}]
  wire  _GEN_1127 = _GEN_2754 & _GEN_2749 ? 1'h0 : _GEN_443; // @[playground/src/noop/dcache.scala 275:{51,51}]
  wire  _GEN_1128 = _GEN_2754 & _GEN_2751 ? 1'h0 : _GEN_444; // @[playground/src/noop/dcache.scala 275:{51,51}]
  wire  _GEN_1129 = _GEN_2754 & _GEN_2753 ? 1'h0 : _GEN_445; // @[playground/src/noop/dcache.scala 275:{51,51}]
  wire  _GEN_1130 = _GEN_2786 & _GEN_2755 ? 1'h0 : _GEN_446; // @[playground/src/noop/dcache.scala 275:{51,51}]
  wire  _GEN_1131 = _GEN_2786 & _GEN_2725 ? 1'h0 : _GEN_447; // @[playground/src/noop/dcache.scala 275:{51,51}]
  wire  _GEN_1132 = _GEN_2786 & _GEN_2727 ? 1'h0 : _GEN_448; // @[playground/src/noop/dcache.scala 275:{51,51}]
  wire  _GEN_1133 = _GEN_2786 & _GEN_2729 ? 1'h0 : _GEN_449; // @[playground/src/noop/dcache.scala 275:{51,51}]
  wire  _GEN_1134 = _GEN_2786 & _GEN_2731 ? 1'h0 : _GEN_450; // @[playground/src/noop/dcache.scala 275:{51,51}]
  wire  _GEN_1135 = _GEN_2786 & _GEN_2733 ? 1'h0 : _GEN_451; // @[playground/src/noop/dcache.scala 275:{51,51}]
  wire  _GEN_1136 = _GEN_2786 & _GEN_2735 ? 1'h0 : _GEN_452; // @[playground/src/noop/dcache.scala 275:{51,51}]
  wire  _GEN_1137 = _GEN_2786 & _GEN_2737 ? 1'h0 : _GEN_453; // @[playground/src/noop/dcache.scala 275:{51,51}]
  wire  _GEN_1138 = _GEN_2786 & _GEN_2739 ? 1'h0 : _GEN_454; // @[playground/src/noop/dcache.scala 275:{51,51}]
  wire  _GEN_1139 = _GEN_2786 & _GEN_2741 ? 1'h0 : _GEN_455; // @[playground/src/noop/dcache.scala 275:{51,51}]
  wire  _GEN_1140 = _GEN_2786 & _GEN_2743 ? 1'h0 : _GEN_456; // @[playground/src/noop/dcache.scala 275:{51,51}]
  wire  _GEN_1141 = _GEN_2786 & _GEN_2745 ? 1'h0 : _GEN_457; // @[playground/src/noop/dcache.scala 275:{51,51}]
  wire  _GEN_1142 = _GEN_2786 & _GEN_2747 ? 1'h0 : _GEN_458; // @[playground/src/noop/dcache.scala 275:{51,51}]
  wire  _GEN_1143 = _GEN_2786 & _GEN_2749 ? 1'h0 : _GEN_459; // @[playground/src/noop/dcache.scala 275:{51,51}]
  wire  _GEN_1144 = _GEN_2786 & _GEN_2751 ? 1'h0 : _GEN_460; // @[playground/src/noop/dcache.scala 275:{51,51}]
  wire  _GEN_1145 = _GEN_2786 & _GEN_2753 ? 1'h0 : _GEN_461; // @[playground/src/noop/dcache.scala 275:{51,51}]
  wire  _GEN_1146 = _GEN_2818 & _GEN_2755 ? 1'h0 : _GEN_462; // @[playground/src/noop/dcache.scala 275:{51,51}]
  wire  _GEN_1147 = _GEN_2818 & _GEN_2725 ? 1'h0 : _GEN_463; // @[playground/src/noop/dcache.scala 275:{51,51}]
  wire  _GEN_1148 = _GEN_2818 & _GEN_2727 ? 1'h0 : _GEN_464; // @[playground/src/noop/dcache.scala 275:{51,51}]
  wire  _GEN_1149 = _GEN_2818 & _GEN_2729 ? 1'h0 : _GEN_465; // @[playground/src/noop/dcache.scala 275:{51,51}]
  wire  _GEN_1150 = _GEN_2818 & _GEN_2731 ? 1'h0 : _GEN_466; // @[playground/src/noop/dcache.scala 275:{51,51}]
  wire  _GEN_1151 = _GEN_2818 & _GEN_2733 ? 1'h0 : _GEN_467; // @[playground/src/noop/dcache.scala 275:{51,51}]
  wire  _GEN_1152 = _GEN_2818 & _GEN_2735 ? 1'h0 : _GEN_468; // @[playground/src/noop/dcache.scala 275:{51,51}]
  wire  _GEN_1153 = _GEN_2818 & _GEN_2737 ? 1'h0 : _GEN_469; // @[playground/src/noop/dcache.scala 275:{51,51}]
  wire  _GEN_1154 = _GEN_2818 & _GEN_2739 ? 1'h0 : _GEN_470; // @[playground/src/noop/dcache.scala 275:{51,51}]
  wire  _GEN_1155 = _GEN_2818 & _GEN_2741 ? 1'h0 : _GEN_471; // @[playground/src/noop/dcache.scala 275:{51,51}]
  wire  _GEN_1156 = _GEN_2818 & _GEN_2743 ? 1'h0 : _GEN_472; // @[playground/src/noop/dcache.scala 275:{51,51}]
  wire  _GEN_1157 = _GEN_2818 & _GEN_2745 ? 1'h0 : _GEN_473; // @[playground/src/noop/dcache.scala 275:{51,51}]
  wire  _GEN_1158 = _GEN_2818 & _GEN_2747 ? 1'h0 : _GEN_474; // @[playground/src/noop/dcache.scala 275:{51,51}]
  wire  _GEN_1159 = _GEN_2818 & _GEN_2749 ? 1'h0 : _GEN_475; // @[playground/src/noop/dcache.scala 275:{51,51}]
  wire  _GEN_1160 = _GEN_2818 & _GEN_2751 ? 1'h0 : _GEN_476; // @[playground/src/noop/dcache.scala 275:{51,51}]
  wire  _GEN_1161 = _GEN_2818 & _GEN_2753 ? 1'h0 : _GEN_477; // @[playground/src/noop/dcache.scala 275:{51,51}]
  wire [2:0] _GEN_1162 = io_dataAxi_wd_bits_last ? 3'h0 : state; // @[playground/src/noop/dcache.scala 152:24 271:46 272:27]
  wire  _GEN_1164 = io_dataAxi_wd_bits_last ? _GEN_1034 : valid_0_0; // @[playground/src/noop/dcache.scala 271:46 89:26]
  wire  _GEN_1165 = io_dataAxi_wd_bits_last ? _GEN_1035 : valid_0_1; // @[playground/src/noop/dcache.scala 271:46 89:26]
  wire  _GEN_1166 = io_dataAxi_wd_bits_last ? _GEN_1036 : valid_0_2; // @[playground/src/noop/dcache.scala 271:46 89:26]
  wire  _GEN_1167 = io_dataAxi_wd_bits_last ? _GEN_1037 : valid_0_3; // @[playground/src/noop/dcache.scala 271:46 89:26]
  wire  _GEN_1168 = io_dataAxi_wd_bits_last ? _GEN_1038 : valid_0_4; // @[playground/src/noop/dcache.scala 271:46 89:26]
  wire  _GEN_1169 = io_dataAxi_wd_bits_last ? _GEN_1039 : valid_0_5; // @[playground/src/noop/dcache.scala 271:46 89:26]
  wire  _GEN_1170 = io_dataAxi_wd_bits_last ? _GEN_1040 : valid_0_6; // @[playground/src/noop/dcache.scala 271:46 89:26]
  wire  _GEN_1171 = io_dataAxi_wd_bits_last ? _GEN_1041 : valid_0_7; // @[playground/src/noop/dcache.scala 271:46 89:26]
  wire  _GEN_1172 = io_dataAxi_wd_bits_last ? _GEN_1042 : valid_0_8; // @[playground/src/noop/dcache.scala 271:46 89:26]
  wire  _GEN_1173 = io_dataAxi_wd_bits_last ? _GEN_1043 : valid_0_9; // @[playground/src/noop/dcache.scala 271:46 89:26]
  wire  _GEN_1174 = io_dataAxi_wd_bits_last ? _GEN_1044 : valid_0_10; // @[playground/src/noop/dcache.scala 271:46 89:26]
  wire  _GEN_1175 = io_dataAxi_wd_bits_last ? _GEN_1045 : valid_0_11; // @[playground/src/noop/dcache.scala 271:46 89:26]
  wire  _GEN_1176 = io_dataAxi_wd_bits_last ? _GEN_1046 : valid_0_12; // @[playground/src/noop/dcache.scala 271:46 89:26]
  wire  _GEN_1177 = io_dataAxi_wd_bits_last ? _GEN_1047 : valid_0_13; // @[playground/src/noop/dcache.scala 271:46 89:26]
  wire  _GEN_1178 = io_dataAxi_wd_bits_last ? _GEN_1048 : valid_0_14; // @[playground/src/noop/dcache.scala 271:46 89:26]
  wire  _GEN_1179 = io_dataAxi_wd_bits_last ? _GEN_1049 : valid_0_15; // @[playground/src/noop/dcache.scala 271:46 89:26]
  wire  _GEN_1180 = io_dataAxi_wd_bits_last ? _GEN_1050 : valid_1_0; // @[playground/src/noop/dcache.scala 271:46 89:26]
  wire  _GEN_1181 = io_dataAxi_wd_bits_last ? _GEN_1051 : valid_1_1; // @[playground/src/noop/dcache.scala 271:46 89:26]
  wire  _GEN_1182 = io_dataAxi_wd_bits_last ? _GEN_1052 : valid_1_2; // @[playground/src/noop/dcache.scala 271:46 89:26]
  wire  _GEN_1183 = io_dataAxi_wd_bits_last ? _GEN_1053 : valid_1_3; // @[playground/src/noop/dcache.scala 271:46 89:26]
  wire  _GEN_1184 = io_dataAxi_wd_bits_last ? _GEN_1054 : valid_1_4; // @[playground/src/noop/dcache.scala 271:46 89:26]
  wire  _GEN_1185 = io_dataAxi_wd_bits_last ? _GEN_1055 : valid_1_5; // @[playground/src/noop/dcache.scala 271:46 89:26]
  wire  _GEN_1186 = io_dataAxi_wd_bits_last ? _GEN_1056 : valid_1_6; // @[playground/src/noop/dcache.scala 271:46 89:26]
  wire  _GEN_1187 = io_dataAxi_wd_bits_last ? _GEN_1057 : valid_1_7; // @[playground/src/noop/dcache.scala 271:46 89:26]
  wire  _GEN_1188 = io_dataAxi_wd_bits_last ? _GEN_1058 : valid_1_8; // @[playground/src/noop/dcache.scala 271:46 89:26]
  wire  _GEN_1189 = io_dataAxi_wd_bits_last ? _GEN_1059 : valid_1_9; // @[playground/src/noop/dcache.scala 271:46 89:26]
  wire  _GEN_1190 = io_dataAxi_wd_bits_last ? _GEN_1060 : valid_1_10; // @[playground/src/noop/dcache.scala 271:46 89:26]
  wire  _GEN_1191 = io_dataAxi_wd_bits_last ? _GEN_1061 : valid_1_11; // @[playground/src/noop/dcache.scala 271:46 89:26]
  wire  _GEN_1192 = io_dataAxi_wd_bits_last ? _GEN_1062 : valid_1_12; // @[playground/src/noop/dcache.scala 271:46 89:26]
  wire  _GEN_1193 = io_dataAxi_wd_bits_last ? _GEN_1063 : valid_1_13; // @[playground/src/noop/dcache.scala 271:46 89:26]
  wire  _GEN_1194 = io_dataAxi_wd_bits_last ? _GEN_1064 : valid_1_14; // @[playground/src/noop/dcache.scala 271:46 89:26]
  wire  _GEN_1195 = io_dataAxi_wd_bits_last ? _GEN_1065 : valid_1_15; // @[playground/src/noop/dcache.scala 271:46 89:26]
  wire  _GEN_1196 = io_dataAxi_wd_bits_last ? _GEN_1066 : valid_2_0; // @[playground/src/noop/dcache.scala 271:46 89:26]
  wire  _GEN_1197 = io_dataAxi_wd_bits_last ? _GEN_1067 : valid_2_1; // @[playground/src/noop/dcache.scala 271:46 89:26]
  wire  _GEN_1198 = io_dataAxi_wd_bits_last ? _GEN_1068 : valid_2_2; // @[playground/src/noop/dcache.scala 271:46 89:26]
  wire  _GEN_1199 = io_dataAxi_wd_bits_last ? _GEN_1069 : valid_2_3; // @[playground/src/noop/dcache.scala 271:46 89:26]
  wire  _GEN_1200 = io_dataAxi_wd_bits_last ? _GEN_1070 : valid_2_4; // @[playground/src/noop/dcache.scala 271:46 89:26]
  wire  _GEN_1201 = io_dataAxi_wd_bits_last ? _GEN_1071 : valid_2_5; // @[playground/src/noop/dcache.scala 271:46 89:26]
  wire  _GEN_1202 = io_dataAxi_wd_bits_last ? _GEN_1072 : valid_2_6; // @[playground/src/noop/dcache.scala 271:46 89:26]
  wire  _GEN_1203 = io_dataAxi_wd_bits_last ? _GEN_1073 : valid_2_7; // @[playground/src/noop/dcache.scala 271:46 89:26]
  wire  _GEN_1204 = io_dataAxi_wd_bits_last ? _GEN_1074 : valid_2_8; // @[playground/src/noop/dcache.scala 271:46 89:26]
  wire  _GEN_1205 = io_dataAxi_wd_bits_last ? _GEN_1075 : valid_2_9; // @[playground/src/noop/dcache.scala 271:46 89:26]
  wire  _GEN_1206 = io_dataAxi_wd_bits_last ? _GEN_1076 : valid_2_10; // @[playground/src/noop/dcache.scala 271:46 89:26]
  wire  _GEN_1207 = io_dataAxi_wd_bits_last ? _GEN_1077 : valid_2_11; // @[playground/src/noop/dcache.scala 271:46 89:26]
  wire  _GEN_1208 = io_dataAxi_wd_bits_last ? _GEN_1078 : valid_2_12; // @[playground/src/noop/dcache.scala 271:46 89:26]
  wire  _GEN_1209 = io_dataAxi_wd_bits_last ? _GEN_1079 : valid_2_13; // @[playground/src/noop/dcache.scala 271:46 89:26]
  wire  _GEN_1210 = io_dataAxi_wd_bits_last ? _GEN_1080 : valid_2_14; // @[playground/src/noop/dcache.scala 271:46 89:26]
  wire  _GEN_1211 = io_dataAxi_wd_bits_last ? _GEN_1081 : valid_2_15; // @[playground/src/noop/dcache.scala 271:46 89:26]
  wire  _GEN_1212 = io_dataAxi_wd_bits_last ? _GEN_1082 : valid_3_0; // @[playground/src/noop/dcache.scala 271:46 89:26]
  wire  _GEN_1213 = io_dataAxi_wd_bits_last ? _GEN_1083 : valid_3_1; // @[playground/src/noop/dcache.scala 271:46 89:26]
  wire  _GEN_1214 = io_dataAxi_wd_bits_last ? _GEN_1084 : valid_3_2; // @[playground/src/noop/dcache.scala 271:46 89:26]
  wire  _GEN_1215 = io_dataAxi_wd_bits_last ? _GEN_1085 : valid_3_3; // @[playground/src/noop/dcache.scala 271:46 89:26]
  wire  _GEN_1216 = io_dataAxi_wd_bits_last ? _GEN_1086 : valid_3_4; // @[playground/src/noop/dcache.scala 271:46 89:26]
  wire  _GEN_1217 = io_dataAxi_wd_bits_last ? _GEN_1087 : valid_3_5; // @[playground/src/noop/dcache.scala 271:46 89:26]
  wire  _GEN_1218 = io_dataAxi_wd_bits_last ? _GEN_1088 : valid_3_6; // @[playground/src/noop/dcache.scala 271:46 89:26]
  wire  _GEN_1219 = io_dataAxi_wd_bits_last ? _GEN_1089 : valid_3_7; // @[playground/src/noop/dcache.scala 271:46 89:26]
  wire  _GEN_1220 = io_dataAxi_wd_bits_last ? _GEN_1090 : valid_3_8; // @[playground/src/noop/dcache.scala 271:46 89:26]
  wire  _GEN_1221 = io_dataAxi_wd_bits_last ? _GEN_1091 : valid_3_9; // @[playground/src/noop/dcache.scala 271:46 89:26]
  wire  _GEN_1222 = io_dataAxi_wd_bits_last ? _GEN_1092 : valid_3_10; // @[playground/src/noop/dcache.scala 271:46 89:26]
  wire  _GEN_1223 = io_dataAxi_wd_bits_last ? _GEN_1093 : valid_3_11; // @[playground/src/noop/dcache.scala 271:46 89:26]
  wire  _GEN_1224 = io_dataAxi_wd_bits_last ? _GEN_1094 : valid_3_12; // @[playground/src/noop/dcache.scala 271:46 89:26]
  wire  _GEN_1225 = io_dataAxi_wd_bits_last ? _GEN_1095 : valid_3_13; // @[playground/src/noop/dcache.scala 271:46 89:26]
  wire  _GEN_1226 = io_dataAxi_wd_bits_last ? _GEN_1096 : valid_3_14; // @[playground/src/noop/dcache.scala 271:46 89:26]
  wire  _GEN_1227 = io_dataAxi_wd_bits_last ? _GEN_1097 : valid_3_15; // @[playground/src/noop/dcache.scala 271:46 89:26]
  wire  _GEN_1228 = io_dataAxi_wd_bits_last ? _GEN_1098 : _GEN_414; // @[playground/src/noop/dcache.scala 271:46]
  wire  _GEN_1229 = io_dataAxi_wd_bits_last ? _GEN_1099 : _GEN_415; // @[playground/src/noop/dcache.scala 271:46]
  wire  _GEN_1230 = io_dataAxi_wd_bits_last ? _GEN_1100 : _GEN_416; // @[playground/src/noop/dcache.scala 271:46]
  wire  _GEN_1231 = io_dataAxi_wd_bits_last ? _GEN_1101 : _GEN_417; // @[playground/src/noop/dcache.scala 271:46]
  wire  _GEN_1232 = io_dataAxi_wd_bits_last ? _GEN_1102 : _GEN_418; // @[playground/src/noop/dcache.scala 271:46]
  wire  _GEN_1233 = io_dataAxi_wd_bits_last ? _GEN_1103 : _GEN_419; // @[playground/src/noop/dcache.scala 271:46]
  wire  _GEN_1234 = io_dataAxi_wd_bits_last ? _GEN_1104 : _GEN_420; // @[playground/src/noop/dcache.scala 271:46]
  wire  _GEN_1235 = io_dataAxi_wd_bits_last ? _GEN_1105 : _GEN_421; // @[playground/src/noop/dcache.scala 271:46]
  wire  _GEN_1236 = io_dataAxi_wd_bits_last ? _GEN_1106 : _GEN_422; // @[playground/src/noop/dcache.scala 271:46]
  wire  _GEN_1237 = io_dataAxi_wd_bits_last ? _GEN_1107 : _GEN_423; // @[playground/src/noop/dcache.scala 271:46]
  wire  _GEN_1238 = io_dataAxi_wd_bits_last ? _GEN_1108 : _GEN_424; // @[playground/src/noop/dcache.scala 271:46]
  wire  _GEN_1239 = io_dataAxi_wd_bits_last ? _GEN_1109 : _GEN_425; // @[playground/src/noop/dcache.scala 271:46]
  wire  _GEN_1240 = io_dataAxi_wd_bits_last ? _GEN_1110 : _GEN_426; // @[playground/src/noop/dcache.scala 271:46]
  wire  _GEN_1241 = io_dataAxi_wd_bits_last ? _GEN_1111 : _GEN_427; // @[playground/src/noop/dcache.scala 271:46]
  wire  _GEN_1242 = io_dataAxi_wd_bits_last ? _GEN_1112 : _GEN_428; // @[playground/src/noop/dcache.scala 271:46]
  wire  _GEN_1243 = io_dataAxi_wd_bits_last ? _GEN_1113 : _GEN_429; // @[playground/src/noop/dcache.scala 271:46]
  wire  _GEN_1244 = io_dataAxi_wd_bits_last ? _GEN_1114 : _GEN_430; // @[playground/src/noop/dcache.scala 271:46]
  wire  _GEN_1245 = io_dataAxi_wd_bits_last ? _GEN_1115 : _GEN_431; // @[playground/src/noop/dcache.scala 271:46]
  wire  _GEN_1246 = io_dataAxi_wd_bits_last ? _GEN_1116 : _GEN_432; // @[playground/src/noop/dcache.scala 271:46]
  wire  _GEN_1247 = io_dataAxi_wd_bits_last ? _GEN_1117 : _GEN_433; // @[playground/src/noop/dcache.scala 271:46]
  wire  _GEN_1248 = io_dataAxi_wd_bits_last ? _GEN_1118 : _GEN_434; // @[playground/src/noop/dcache.scala 271:46]
  wire  _GEN_1249 = io_dataAxi_wd_bits_last ? _GEN_1119 : _GEN_435; // @[playground/src/noop/dcache.scala 271:46]
  wire  _GEN_1250 = io_dataAxi_wd_bits_last ? _GEN_1120 : _GEN_436; // @[playground/src/noop/dcache.scala 271:46]
  wire  _GEN_1251 = io_dataAxi_wd_bits_last ? _GEN_1121 : _GEN_437; // @[playground/src/noop/dcache.scala 271:46]
  wire  _GEN_1252 = io_dataAxi_wd_bits_last ? _GEN_1122 : _GEN_438; // @[playground/src/noop/dcache.scala 271:46]
  wire  _GEN_1253 = io_dataAxi_wd_bits_last ? _GEN_1123 : _GEN_439; // @[playground/src/noop/dcache.scala 271:46]
  wire  _GEN_1254 = io_dataAxi_wd_bits_last ? _GEN_1124 : _GEN_440; // @[playground/src/noop/dcache.scala 271:46]
  wire  _GEN_1255 = io_dataAxi_wd_bits_last ? _GEN_1125 : _GEN_441; // @[playground/src/noop/dcache.scala 271:46]
  wire  _GEN_1256 = io_dataAxi_wd_bits_last ? _GEN_1126 : _GEN_442; // @[playground/src/noop/dcache.scala 271:46]
  wire  _GEN_1257 = io_dataAxi_wd_bits_last ? _GEN_1127 : _GEN_443; // @[playground/src/noop/dcache.scala 271:46]
  wire  _GEN_1258 = io_dataAxi_wd_bits_last ? _GEN_1128 : _GEN_444; // @[playground/src/noop/dcache.scala 271:46]
  wire  _GEN_1259 = io_dataAxi_wd_bits_last ? _GEN_1129 : _GEN_445; // @[playground/src/noop/dcache.scala 271:46]
  wire  _GEN_1260 = io_dataAxi_wd_bits_last ? _GEN_1130 : _GEN_446; // @[playground/src/noop/dcache.scala 271:46]
  wire  _GEN_1261 = io_dataAxi_wd_bits_last ? _GEN_1131 : _GEN_447; // @[playground/src/noop/dcache.scala 271:46]
  wire  _GEN_1262 = io_dataAxi_wd_bits_last ? _GEN_1132 : _GEN_448; // @[playground/src/noop/dcache.scala 271:46]
  wire  _GEN_1263 = io_dataAxi_wd_bits_last ? _GEN_1133 : _GEN_449; // @[playground/src/noop/dcache.scala 271:46]
  wire  _GEN_1264 = io_dataAxi_wd_bits_last ? _GEN_1134 : _GEN_450; // @[playground/src/noop/dcache.scala 271:46]
  wire  _GEN_1265 = io_dataAxi_wd_bits_last ? _GEN_1135 : _GEN_451; // @[playground/src/noop/dcache.scala 271:46]
  wire  _GEN_1266 = io_dataAxi_wd_bits_last ? _GEN_1136 : _GEN_452; // @[playground/src/noop/dcache.scala 271:46]
  wire  _GEN_1267 = io_dataAxi_wd_bits_last ? _GEN_1137 : _GEN_453; // @[playground/src/noop/dcache.scala 271:46]
  wire  _GEN_1268 = io_dataAxi_wd_bits_last ? _GEN_1138 : _GEN_454; // @[playground/src/noop/dcache.scala 271:46]
  wire  _GEN_1269 = io_dataAxi_wd_bits_last ? _GEN_1139 : _GEN_455; // @[playground/src/noop/dcache.scala 271:46]
  wire  _GEN_1270 = io_dataAxi_wd_bits_last ? _GEN_1140 : _GEN_456; // @[playground/src/noop/dcache.scala 271:46]
  wire  _GEN_1271 = io_dataAxi_wd_bits_last ? _GEN_1141 : _GEN_457; // @[playground/src/noop/dcache.scala 271:46]
  wire  _GEN_1272 = io_dataAxi_wd_bits_last ? _GEN_1142 : _GEN_458; // @[playground/src/noop/dcache.scala 271:46]
  wire  _GEN_1273 = io_dataAxi_wd_bits_last ? _GEN_1143 : _GEN_459; // @[playground/src/noop/dcache.scala 271:46]
  wire  _GEN_1274 = io_dataAxi_wd_bits_last ? _GEN_1144 : _GEN_460; // @[playground/src/noop/dcache.scala 271:46]
  wire  _GEN_1275 = io_dataAxi_wd_bits_last ? _GEN_1145 : _GEN_461; // @[playground/src/noop/dcache.scala 271:46]
  wire  _GEN_1276 = io_dataAxi_wd_bits_last ? _GEN_1146 : _GEN_462; // @[playground/src/noop/dcache.scala 271:46]
  wire  _GEN_1277 = io_dataAxi_wd_bits_last ? _GEN_1147 : _GEN_463; // @[playground/src/noop/dcache.scala 271:46]
  wire  _GEN_1278 = io_dataAxi_wd_bits_last ? _GEN_1148 : _GEN_464; // @[playground/src/noop/dcache.scala 271:46]
  wire  _GEN_1279 = io_dataAxi_wd_bits_last ? _GEN_1149 : _GEN_465; // @[playground/src/noop/dcache.scala 271:46]
  wire  _GEN_1280 = io_dataAxi_wd_bits_last ? _GEN_1150 : _GEN_466; // @[playground/src/noop/dcache.scala 271:46]
  wire  _GEN_1281 = io_dataAxi_wd_bits_last ? _GEN_1151 : _GEN_467; // @[playground/src/noop/dcache.scala 271:46]
  wire  _GEN_1282 = io_dataAxi_wd_bits_last ? _GEN_1152 : _GEN_468; // @[playground/src/noop/dcache.scala 271:46]
  wire  _GEN_1283 = io_dataAxi_wd_bits_last ? _GEN_1153 : _GEN_469; // @[playground/src/noop/dcache.scala 271:46]
  wire  _GEN_1284 = io_dataAxi_wd_bits_last ? _GEN_1154 : _GEN_470; // @[playground/src/noop/dcache.scala 271:46]
  wire  _GEN_1285 = io_dataAxi_wd_bits_last ? _GEN_1155 : _GEN_471; // @[playground/src/noop/dcache.scala 271:46]
  wire  _GEN_1286 = io_dataAxi_wd_bits_last ? _GEN_1156 : _GEN_472; // @[playground/src/noop/dcache.scala 271:46]
  wire  _GEN_1287 = io_dataAxi_wd_bits_last ? _GEN_1157 : _GEN_473; // @[playground/src/noop/dcache.scala 271:46]
  wire  _GEN_1288 = io_dataAxi_wd_bits_last ? _GEN_1158 : _GEN_474; // @[playground/src/noop/dcache.scala 271:46]
  wire  _GEN_1289 = io_dataAxi_wd_bits_last ? _GEN_1159 : _GEN_475; // @[playground/src/noop/dcache.scala 271:46]
  wire  _GEN_1290 = io_dataAxi_wd_bits_last ? _GEN_1160 : _GEN_476; // @[playground/src/noop/dcache.scala 271:46]
  wire  _GEN_1291 = io_dataAxi_wd_bits_last ? _GEN_1161 : _GEN_477; // @[playground/src/noop/dcache.scala 271:46]
  wire [2:0] _GEN_1292 = axiWdataEn & io_dataAxi_wd_ready ? _offset_T_1 : offset; // @[playground/src/noop/dcache.scala 268:52 269:24 110:34]
  wire  _GEN_1293 = axiWdataEn & io_dataAxi_wd_ready ? 1'h0 : 1'h1; // @[playground/src/noop/dcache.scala 267:24 268:52]
  wire [2:0] _GEN_1294 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1162 : state; // @[playground/src/noop/dcache.scala 152:24 268:52]
  wire  _GEN_1295 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1164 : valid_0_0; // @[playground/src/noop/dcache.scala 268:52 89:26]
  wire  _GEN_1296 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1165 : valid_0_1; // @[playground/src/noop/dcache.scala 268:52 89:26]
  wire  _GEN_1297 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1166 : valid_0_2; // @[playground/src/noop/dcache.scala 268:52 89:26]
  wire  _GEN_1298 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1167 : valid_0_3; // @[playground/src/noop/dcache.scala 268:52 89:26]
  wire  _GEN_1299 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1168 : valid_0_4; // @[playground/src/noop/dcache.scala 268:52 89:26]
  wire  _GEN_1300 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1169 : valid_0_5; // @[playground/src/noop/dcache.scala 268:52 89:26]
  wire  _GEN_1301 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1170 : valid_0_6; // @[playground/src/noop/dcache.scala 268:52 89:26]
  wire  _GEN_1302 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1171 : valid_0_7; // @[playground/src/noop/dcache.scala 268:52 89:26]
  wire  _GEN_1303 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1172 : valid_0_8; // @[playground/src/noop/dcache.scala 268:52 89:26]
  wire  _GEN_1304 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1173 : valid_0_9; // @[playground/src/noop/dcache.scala 268:52 89:26]
  wire  _GEN_1305 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1174 : valid_0_10; // @[playground/src/noop/dcache.scala 268:52 89:26]
  wire  _GEN_1306 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1175 : valid_0_11; // @[playground/src/noop/dcache.scala 268:52 89:26]
  wire  _GEN_1307 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1176 : valid_0_12; // @[playground/src/noop/dcache.scala 268:52 89:26]
  wire  _GEN_1308 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1177 : valid_0_13; // @[playground/src/noop/dcache.scala 268:52 89:26]
  wire  _GEN_1309 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1178 : valid_0_14; // @[playground/src/noop/dcache.scala 268:52 89:26]
  wire  _GEN_1310 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1179 : valid_0_15; // @[playground/src/noop/dcache.scala 268:52 89:26]
  wire  _GEN_1311 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1180 : valid_1_0; // @[playground/src/noop/dcache.scala 268:52 89:26]
  wire  _GEN_1312 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1181 : valid_1_1; // @[playground/src/noop/dcache.scala 268:52 89:26]
  wire  _GEN_1313 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1182 : valid_1_2; // @[playground/src/noop/dcache.scala 268:52 89:26]
  wire  _GEN_1314 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1183 : valid_1_3; // @[playground/src/noop/dcache.scala 268:52 89:26]
  wire  _GEN_1315 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1184 : valid_1_4; // @[playground/src/noop/dcache.scala 268:52 89:26]
  wire  _GEN_1316 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1185 : valid_1_5; // @[playground/src/noop/dcache.scala 268:52 89:26]
  wire  _GEN_1317 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1186 : valid_1_6; // @[playground/src/noop/dcache.scala 268:52 89:26]
  wire  _GEN_1318 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1187 : valid_1_7; // @[playground/src/noop/dcache.scala 268:52 89:26]
  wire  _GEN_1319 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1188 : valid_1_8; // @[playground/src/noop/dcache.scala 268:52 89:26]
  wire  _GEN_1320 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1189 : valid_1_9; // @[playground/src/noop/dcache.scala 268:52 89:26]
  wire  _GEN_1321 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1190 : valid_1_10; // @[playground/src/noop/dcache.scala 268:52 89:26]
  wire  _GEN_1322 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1191 : valid_1_11; // @[playground/src/noop/dcache.scala 268:52 89:26]
  wire  _GEN_1323 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1192 : valid_1_12; // @[playground/src/noop/dcache.scala 268:52 89:26]
  wire  _GEN_1324 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1193 : valid_1_13; // @[playground/src/noop/dcache.scala 268:52 89:26]
  wire  _GEN_1325 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1194 : valid_1_14; // @[playground/src/noop/dcache.scala 268:52 89:26]
  wire  _GEN_1326 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1195 : valid_1_15; // @[playground/src/noop/dcache.scala 268:52 89:26]
  wire  _GEN_1327 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1196 : valid_2_0; // @[playground/src/noop/dcache.scala 268:52 89:26]
  wire  _GEN_1328 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1197 : valid_2_1; // @[playground/src/noop/dcache.scala 268:52 89:26]
  wire  _GEN_1329 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1198 : valid_2_2; // @[playground/src/noop/dcache.scala 268:52 89:26]
  wire  _GEN_1330 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1199 : valid_2_3; // @[playground/src/noop/dcache.scala 268:52 89:26]
  wire  _GEN_1331 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1200 : valid_2_4; // @[playground/src/noop/dcache.scala 268:52 89:26]
  wire  _GEN_1332 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1201 : valid_2_5; // @[playground/src/noop/dcache.scala 268:52 89:26]
  wire  _GEN_1333 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1202 : valid_2_6; // @[playground/src/noop/dcache.scala 268:52 89:26]
  wire  _GEN_1334 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1203 : valid_2_7; // @[playground/src/noop/dcache.scala 268:52 89:26]
  wire  _GEN_1335 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1204 : valid_2_8; // @[playground/src/noop/dcache.scala 268:52 89:26]
  wire  _GEN_1336 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1205 : valid_2_9; // @[playground/src/noop/dcache.scala 268:52 89:26]
  wire  _GEN_1337 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1206 : valid_2_10; // @[playground/src/noop/dcache.scala 268:52 89:26]
  wire  _GEN_1338 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1207 : valid_2_11; // @[playground/src/noop/dcache.scala 268:52 89:26]
  wire  _GEN_1339 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1208 : valid_2_12; // @[playground/src/noop/dcache.scala 268:52 89:26]
  wire  _GEN_1340 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1209 : valid_2_13; // @[playground/src/noop/dcache.scala 268:52 89:26]
  wire  _GEN_1341 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1210 : valid_2_14; // @[playground/src/noop/dcache.scala 268:52 89:26]
  wire  _GEN_1342 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1211 : valid_2_15; // @[playground/src/noop/dcache.scala 268:52 89:26]
  wire  _GEN_1343 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1212 : valid_3_0; // @[playground/src/noop/dcache.scala 268:52 89:26]
  wire  _GEN_1344 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1213 : valid_3_1; // @[playground/src/noop/dcache.scala 268:52 89:26]
  wire  _GEN_1345 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1214 : valid_3_2; // @[playground/src/noop/dcache.scala 268:52 89:26]
  wire  _GEN_1346 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1215 : valid_3_3; // @[playground/src/noop/dcache.scala 268:52 89:26]
  wire  _GEN_1347 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1216 : valid_3_4; // @[playground/src/noop/dcache.scala 268:52 89:26]
  wire  _GEN_1348 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1217 : valid_3_5; // @[playground/src/noop/dcache.scala 268:52 89:26]
  wire  _GEN_1349 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1218 : valid_3_6; // @[playground/src/noop/dcache.scala 268:52 89:26]
  wire  _GEN_1350 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1219 : valid_3_7; // @[playground/src/noop/dcache.scala 268:52 89:26]
  wire  _GEN_1351 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1220 : valid_3_8; // @[playground/src/noop/dcache.scala 268:52 89:26]
  wire  _GEN_1352 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1221 : valid_3_9; // @[playground/src/noop/dcache.scala 268:52 89:26]
  wire  _GEN_1353 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1222 : valid_3_10; // @[playground/src/noop/dcache.scala 268:52 89:26]
  wire  _GEN_1354 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1223 : valid_3_11; // @[playground/src/noop/dcache.scala 268:52 89:26]
  wire  _GEN_1355 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1224 : valid_3_12; // @[playground/src/noop/dcache.scala 268:52 89:26]
  wire  _GEN_1356 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1225 : valid_3_13; // @[playground/src/noop/dcache.scala 268:52 89:26]
  wire  _GEN_1357 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1226 : valid_3_14; // @[playground/src/noop/dcache.scala 268:52 89:26]
  wire  _GEN_1358 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1227 : valid_3_15; // @[playground/src/noop/dcache.scala 268:52 89:26]
  wire  _GEN_1359 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1228 : _GEN_414; // @[playground/src/noop/dcache.scala 268:52]
  wire  _GEN_1360 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1229 : _GEN_415; // @[playground/src/noop/dcache.scala 268:52]
  wire  _GEN_1361 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1230 : _GEN_416; // @[playground/src/noop/dcache.scala 268:52]
  wire  _GEN_1362 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1231 : _GEN_417; // @[playground/src/noop/dcache.scala 268:52]
  wire  _GEN_1363 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1232 : _GEN_418; // @[playground/src/noop/dcache.scala 268:52]
  wire  _GEN_1364 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1233 : _GEN_419; // @[playground/src/noop/dcache.scala 268:52]
  wire  _GEN_1365 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1234 : _GEN_420; // @[playground/src/noop/dcache.scala 268:52]
  wire  _GEN_1366 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1235 : _GEN_421; // @[playground/src/noop/dcache.scala 268:52]
  wire  _GEN_1367 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1236 : _GEN_422; // @[playground/src/noop/dcache.scala 268:52]
  wire  _GEN_1368 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1237 : _GEN_423; // @[playground/src/noop/dcache.scala 268:52]
  wire  _GEN_1369 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1238 : _GEN_424; // @[playground/src/noop/dcache.scala 268:52]
  wire  _GEN_1370 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1239 : _GEN_425; // @[playground/src/noop/dcache.scala 268:52]
  wire  _GEN_1371 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1240 : _GEN_426; // @[playground/src/noop/dcache.scala 268:52]
  wire  _GEN_1372 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1241 : _GEN_427; // @[playground/src/noop/dcache.scala 268:52]
  wire  _GEN_1373 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1242 : _GEN_428; // @[playground/src/noop/dcache.scala 268:52]
  wire  _GEN_1374 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1243 : _GEN_429; // @[playground/src/noop/dcache.scala 268:52]
  wire  _GEN_1375 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1244 : _GEN_430; // @[playground/src/noop/dcache.scala 268:52]
  wire  _GEN_1376 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1245 : _GEN_431; // @[playground/src/noop/dcache.scala 268:52]
  wire  _GEN_1377 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1246 : _GEN_432; // @[playground/src/noop/dcache.scala 268:52]
  wire  _GEN_1378 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1247 : _GEN_433; // @[playground/src/noop/dcache.scala 268:52]
  wire  _GEN_1379 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1248 : _GEN_434; // @[playground/src/noop/dcache.scala 268:52]
  wire  _GEN_1380 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1249 : _GEN_435; // @[playground/src/noop/dcache.scala 268:52]
  wire  _GEN_1381 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1250 : _GEN_436; // @[playground/src/noop/dcache.scala 268:52]
  wire  _GEN_1382 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1251 : _GEN_437; // @[playground/src/noop/dcache.scala 268:52]
  wire  _GEN_1383 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1252 : _GEN_438; // @[playground/src/noop/dcache.scala 268:52]
  wire  _GEN_1384 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1253 : _GEN_439; // @[playground/src/noop/dcache.scala 268:52]
  wire  _GEN_1385 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1254 : _GEN_440; // @[playground/src/noop/dcache.scala 268:52]
  wire  _GEN_1386 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1255 : _GEN_441; // @[playground/src/noop/dcache.scala 268:52]
  wire  _GEN_1387 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1256 : _GEN_442; // @[playground/src/noop/dcache.scala 268:52]
  wire  _GEN_1388 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1257 : _GEN_443; // @[playground/src/noop/dcache.scala 268:52]
  wire  _GEN_1389 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1258 : _GEN_444; // @[playground/src/noop/dcache.scala 268:52]
  wire  _GEN_1390 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1259 : _GEN_445; // @[playground/src/noop/dcache.scala 268:52]
  wire  _GEN_1391 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1260 : _GEN_446; // @[playground/src/noop/dcache.scala 268:52]
  wire  _GEN_1392 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1261 : _GEN_447; // @[playground/src/noop/dcache.scala 268:52]
  wire  _GEN_1393 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1262 : _GEN_448; // @[playground/src/noop/dcache.scala 268:52]
  wire  _GEN_1394 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1263 : _GEN_449; // @[playground/src/noop/dcache.scala 268:52]
  wire  _GEN_1395 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1264 : _GEN_450; // @[playground/src/noop/dcache.scala 268:52]
  wire  _GEN_1396 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1265 : _GEN_451; // @[playground/src/noop/dcache.scala 268:52]
  wire  _GEN_1397 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1266 : _GEN_452; // @[playground/src/noop/dcache.scala 268:52]
  wire  _GEN_1398 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1267 : _GEN_453; // @[playground/src/noop/dcache.scala 268:52]
  wire  _GEN_1399 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1268 : _GEN_454; // @[playground/src/noop/dcache.scala 268:52]
  wire  _GEN_1400 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1269 : _GEN_455; // @[playground/src/noop/dcache.scala 268:52]
  wire  _GEN_1401 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1270 : _GEN_456; // @[playground/src/noop/dcache.scala 268:52]
  wire  _GEN_1402 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1271 : _GEN_457; // @[playground/src/noop/dcache.scala 268:52]
  wire  _GEN_1403 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1272 : _GEN_458; // @[playground/src/noop/dcache.scala 268:52]
  wire  _GEN_1404 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1273 : _GEN_459; // @[playground/src/noop/dcache.scala 268:52]
  wire  _GEN_1405 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1274 : _GEN_460; // @[playground/src/noop/dcache.scala 268:52]
  wire  _GEN_1406 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1275 : _GEN_461; // @[playground/src/noop/dcache.scala 268:52]
  wire  _GEN_1407 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1276 : _GEN_462; // @[playground/src/noop/dcache.scala 268:52]
  wire  _GEN_1408 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1277 : _GEN_463; // @[playground/src/noop/dcache.scala 268:52]
  wire  _GEN_1409 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1278 : _GEN_464; // @[playground/src/noop/dcache.scala 268:52]
  wire  _GEN_1410 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1279 : _GEN_465; // @[playground/src/noop/dcache.scala 268:52]
  wire  _GEN_1411 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1280 : _GEN_466; // @[playground/src/noop/dcache.scala 268:52]
  wire  _GEN_1412 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1281 : _GEN_467; // @[playground/src/noop/dcache.scala 268:52]
  wire  _GEN_1413 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1282 : _GEN_468; // @[playground/src/noop/dcache.scala 268:52]
  wire  _GEN_1414 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1283 : _GEN_469; // @[playground/src/noop/dcache.scala 268:52]
  wire  _GEN_1415 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1284 : _GEN_470; // @[playground/src/noop/dcache.scala 268:52]
  wire  _GEN_1416 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1285 : _GEN_471; // @[playground/src/noop/dcache.scala 268:52]
  wire  _GEN_1417 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1286 : _GEN_472; // @[playground/src/noop/dcache.scala 268:52]
  wire  _GEN_1418 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1287 : _GEN_473; // @[playground/src/noop/dcache.scala 268:52]
  wire  _GEN_1419 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1288 : _GEN_474; // @[playground/src/noop/dcache.scala 268:52]
  wire  _GEN_1420 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1289 : _GEN_475; // @[playground/src/noop/dcache.scala 268:52]
  wire  _GEN_1421 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1290 : _GEN_476; // @[playground/src/noop/dcache.scala 268:52]
  wire  _GEN_1422 = axiWdataEn & io_dataAxi_wd_ready ? _GEN_1291 : _GEN_477; // @[playground/src/noop/dcache.scala 268:52]
  wire  _GEN_1423 = flush_done ? 1'h0 : _GEN_134; // @[playground/src/noop/dcache.scala 286:29 287:25]
  wire [2:0] _GEN_1424 = flush_done ? 3'h0 : 3'h3; // @[playground/src/noop/dcache.scala 286:29 288:23 291:23]
  wire  _GEN_1425 = flush_done ? 1'h0 : valid_0_0; // @[playground/src/noop/dcache.scala 286:29 289:23 89:26]
  wire  _GEN_1426 = flush_done ? 1'h0 : valid_0_1; // @[playground/src/noop/dcache.scala 286:29 289:23 89:26]
  wire  _GEN_1427 = flush_done ? 1'h0 : valid_0_2; // @[playground/src/noop/dcache.scala 286:29 289:23 89:26]
  wire  _GEN_1428 = flush_done ? 1'h0 : valid_0_3; // @[playground/src/noop/dcache.scala 286:29 289:23 89:26]
  wire  _GEN_1429 = flush_done ? 1'h0 : valid_0_4; // @[playground/src/noop/dcache.scala 286:29 289:23 89:26]
  wire  _GEN_1430 = flush_done ? 1'h0 : valid_0_5; // @[playground/src/noop/dcache.scala 286:29 289:23 89:26]
  wire  _GEN_1431 = flush_done ? 1'h0 : valid_0_6; // @[playground/src/noop/dcache.scala 286:29 289:23 89:26]
  wire  _GEN_1432 = flush_done ? 1'h0 : valid_0_7; // @[playground/src/noop/dcache.scala 286:29 289:23 89:26]
  wire  _GEN_1433 = flush_done ? 1'h0 : valid_0_8; // @[playground/src/noop/dcache.scala 286:29 289:23 89:26]
  wire  _GEN_1434 = flush_done ? 1'h0 : valid_0_9; // @[playground/src/noop/dcache.scala 286:29 289:23 89:26]
  wire  _GEN_1435 = flush_done ? 1'h0 : valid_0_10; // @[playground/src/noop/dcache.scala 286:29 289:23 89:26]
  wire  _GEN_1436 = flush_done ? 1'h0 : valid_0_11; // @[playground/src/noop/dcache.scala 286:29 289:23 89:26]
  wire  _GEN_1437 = flush_done ? 1'h0 : valid_0_12; // @[playground/src/noop/dcache.scala 286:29 289:23 89:26]
  wire  _GEN_1438 = flush_done ? 1'h0 : valid_0_13; // @[playground/src/noop/dcache.scala 286:29 289:23 89:26]
  wire  _GEN_1439 = flush_done ? 1'h0 : valid_0_14; // @[playground/src/noop/dcache.scala 286:29 289:23 89:26]
  wire  _GEN_1440 = flush_done ? 1'h0 : valid_0_15; // @[playground/src/noop/dcache.scala 286:29 289:23 89:26]
  wire  _GEN_1441 = flush_done ? 1'h0 : valid_1_0; // @[playground/src/noop/dcache.scala 286:29 289:23 89:26]
  wire  _GEN_1442 = flush_done ? 1'h0 : valid_1_1; // @[playground/src/noop/dcache.scala 286:29 289:23 89:26]
  wire  _GEN_1443 = flush_done ? 1'h0 : valid_1_2; // @[playground/src/noop/dcache.scala 286:29 289:23 89:26]
  wire  _GEN_1444 = flush_done ? 1'h0 : valid_1_3; // @[playground/src/noop/dcache.scala 286:29 289:23 89:26]
  wire  _GEN_1445 = flush_done ? 1'h0 : valid_1_4; // @[playground/src/noop/dcache.scala 286:29 289:23 89:26]
  wire  _GEN_1446 = flush_done ? 1'h0 : valid_1_5; // @[playground/src/noop/dcache.scala 286:29 289:23 89:26]
  wire  _GEN_1447 = flush_done ? 1'h0 : valid_1_6; // @[playground/src/noop/dcache.scala 286:29 289:23 89:26]
  wire  _GEN_1448 = flush_done ? 1'h0 : valid_1_7; // @[playground/src/noop/dcache.scala 286:29 289:23 89:26]
  wire  _GEN_1449 = flush_done ? 1'h0 : valid_1_8; // @[playground/src/noop/dcache.scala 286:29 289:23 89:26]
  wire  _GEN_1450 = flush_done ? 1'h0 : valid_1_9; // @[playground/src/noop/dcache.scala 286:29 289:23 89:26]
  wire  _GEN_1451 = flush_done ? 1'h0 : valid_1_10; // @[playground/src/noop/dcache.scala 286:29 289:23 89:26]
  wire  _GEN_1452 = flush_done ? 1'h0 : valid_1_11; // @[playground/src/noop/dcache.scala 286:29 289:23 89:26]
  wire  _GEN_1453 = flush_done ? 1'h0 : valid_1_12; // @[playground/src/noop/dcache.scala 286:29 289:23 89:26]
  wire  _GEN_1454 = flush_done ? 1'h0 : valid_1_13; // @[playground/src/noop/dcache.scala 286:29 289:23 89:26]
  wire  _GEN_1455 = flush_done ? 1'h0 : valid_1_14; // @[playground/src/noop/dcache.scala 286:29 289:23 89:26]
  wire  _GEN_1456 = flush_done ? 1'h0 : valid_1_15; // @[playground/src/noop/dcache.scala 286:29 289:23 89:26]
  wire  _GEN_1457 = flush_done ? 1'h0 : valid_2_0; // @[playground/src/noop/dcache.scala 286:29 289:23 89:26]
  wire  _GEN_1458 = flush_done ? 1'h0 : valid_2_1; // @[playground/src/noop/dcache.scala 286:29 289:23 89:26]
  wire  _GEN_1459 = flush_done ? 1'h0 : valid_2_2; // @[playground/src/noop/dcache.scala 286:29 289:23 89:26]
  wire  _GEN_1460 = flush_done ? 1'h0 : valid_2_3; // @[playground/src/noop/dcache.scala 286:29 289:23 89:26]
  wire  _GEN_1461 = flush_done ? 1'h0 : valid_2_4; // @[playground/src/noop/dcache.scala 286:29 289:23 89:26]
  wire  _GEN_1462 = flush_done ? 1'h0 : valid_2_5; // @[playground/src/noop/dcache.scala 286:29 289:23 89:26]
  wire  _GEN_1463 = flush_done ? 1'h0 : valid_2_6; // @[playground/src/noop/dcache.scala 286:29 289:23 89:26]
  wire  _GEN_1464 = flush_done ? 1'h0 : valid_2_7; // @[playground/src/noop/dcache.scala 286:29 289:23 89:26]
  wire  _GEN_1465 = flush_done ? 1'h0 : valid_2_8; // @[playground/src/noop/dcache.scala 286:29 289:23 89:26]
  wire  _GEN_1466 = flush_done ? 1'h0 : valid_2_9; // @[playground/src/noop/dcache.scala 286:29 289:23 89:26]
  wire  _GEN_1467 = flush_done ? 1'h0 : valid_2_10; // @[playground/src/noop/dcache.scala 286:29 289:23 89:26]
  wire  _GEN_1468 = flush_done ? 1'h0 : valid_2_11; // @[playground/src/noop/dcache.scala 286:29 289:23 89:26]
  wire  _GEN_1469 = flush_done ? 1'h0 : valid_2_12; // @[playground/src/noop/dcache.scala 286:29 289:23 89:26]
  wire  _GEN_1470 = flush_done ? 1'h0 : valid_2_13; // @[playground/src/noop/dcache.scala 286:29 289:23 89:26]
  wire  _GEN_1471 = flush_done ? 1'h0 : valid_2_14; // @[playground/src/noop/dcache.scala 286:29 289:23 89:26]
  wire  _GEN_1472 = flush_done ? 1'h0 : valid_2_15; // @[playground/src/noop/dcache.scala 286:29 289:23 89:26]
  wire  _GEN_1473 = flush_done ? 1'h0 : valid_3_0; // @[playground/src/noop/dcache.scala 286:29 289:23 89:26]
  wire  _GEN_1474 = flush_done ? 1'h0 : valid_3_1; // @[playground/src/noop/dcache.scala 286:29 289:23 89:26]
  wire  _GEN_1475 = flush_done ? 1'h0 : valid_3_2; // @[playground/src/noop/dcache.scala 286:29 289:23 89:26]
  wire  _GEN_1476 = flush_done ? 1'h0 : valid_3_3; // @[playground/src/noop/dcache.scala 286:29 289:23 89:26]
  wire  _GEN_1477 = flush_done ? 1'h0 : valid_3_4; // @[playground/src/noop/dcache.scala 286:29 289:23 89:26]
  wire  _GEN_1478 = flush_done ? 1'h0 : valid_3_5; // @[playground/src/noop/dcache.scala 286:29 289:23 89:26]
  wire  _GEN_1479 = flush_done ? 1'h0 : valid_3_6; // @[playground/src/noop/dcache.scala 286:29 289:23 89:26]
  wire  _GEN_1480 = flush_done ? 1'h0 : valid_3_7; // @[playground/src/noop/dcache.scala 286:29 289:23 89:26]
  wire  _GEN_1481 = flush_done ? 1'h0 : valid_3_8; // @[playground/src/noop/dcache.scala 286:29 289:23 89:26]
  wire  _GEN_1482 = flush_done ? 1'h0 : valid_3_9; // @[playground/src/noop/dcache.scala 286:29 289:23 89:26]
  wire  _GEN_1483 = flush_done ? 1'h0 : valid_3_10; // @[playground/src/noop/dcache.scala 286:29 289:23 89:26]
  wire  _GEN_1484 = flush_done ? 1'h0 : valid_3_11; // @[playground/src/noop/dcache.scala 286:29 289:23 89:26]
  wire  _GEN_1485 = flush_done ? 1'h0 : valid_3_12; // @[playground/src/noop/dcache.scala 286:29 289:23 89:26]
  wire  _GEN_1486 = flush_done ? 1'h0 : valid_3_13; // @[playground/src/noop/dcache.scala 286:29 289:23 89:26]
  wire  _GEN_1487 = flush_done ? 1'h0 : valid_3_14; // @[playground/src/noop/dcache.scala 286:29 289:23 89:26]
  wire  _GEN_1488 = flush_done ? 1'h0 : valid_3_15; // @[playground/src/noop/dcache.scala 286:29 289:23 89:26]
  wire  _GEN_1489 = flush_done ? axiWaddrEn : 1'h1; // @[playground/src/noop/dcache.scala 286:29 199:34 292:28]
  wire [1:0] _GEN_1490 = flush_done ? _GEN_129 : flush_way; // @[playground/src/noop/dcache.scala 286:29 293:28]
  wire [3:0] _GEN_1491 = flush_done ? _GEN_133 : flush_idx; // @[playground/src/noop/dcache.scala 286:29 294:28]
  wire  _GEN_1492 = 3'h6 == state ? _GEN_1423 : _GEN_134; // @[playground/src/noop/dcache.scala 205:18]
  wire [2:0] _GEN_1493 = 3'h6 == state ? _GEN_1424 : state; // @[playground/src/noop/dcache.scala 205:18 152:24]
  wire  _GEN_1494 = 3'h6 == state ? _GEN_1425 : valid_0_0; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1495 = 3'h6 == state ? _GEN_1426 : valid_0_1; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1496 = 3'h6 == state ? _GEN_1427 : valid_0_2; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1497 = 3'h6 == state ? _GEN_1428 : valid_0_3; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1498 = 3'h6 == state ? _GEN_1429 : valid_0_4; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1499 = 3'h6 == state ? _GEN_1430 : valid_0_5; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1500 = 3'h6 == state ? _GEN_1431 : valid_0_6; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1501 = 3'h6 == state ? _GEN_1432 : valid_0_7; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1502 = 3'h6 == state ? _GEN_1433 : valid_0_8; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1503 = 3'h6 == state ? _GEN_1434 : valid_0_9; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1504 = 3'h6 == state ? _GEN_1435 : valid_0_10; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1505 = 3'h6 == state ? _GEN_1436 : valid_0_11; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1506 = 3'h6 == state ? _GEN_1437 : valid_0_12; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1507 = 3'h6 == state ? _GEN_1438 : valid_0_13; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1508 = 3'h6 == state ? _GEN_1439 : valid_0_14; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1509 = 3'h6 == state ? _GEN_1440 : valid_0_15; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1510 = 3'h6 == state ? _GEN_1441 : valid_1_0; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1511 = 3'h6 == state ? _GEN_1442 : valid_1_1; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1512 = 3'h6 == state ? _GEN_1443 : valid_1_2; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1513 = 3'h6 == state ? _GEN_1444 : valid_1_3; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1514 = 3'h6 == state ? _GEN_1445 : valid_1_4; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1515 = 3'h6 == state ? _GEN_1446 : valid_1_5; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1516 = 3'h6 == state ? _GEN_1447 : valid_1_6; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1517 = 3'h6 == state ? _GEN_1448 : valid_1_7; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1518 = 3'h6 == state ? _GEN_1449 : valid_1_8; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1519 = 3'h6 == state ? _GEN_1450 : valid_1_9; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1520 = 3'h6 == state ? _GEN_1451 : valid_1_10; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1521 = 3'h6 == state ? _GEN_1452 : valid_1_11; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1522 = 3'h6 == state ? _GEN_1453 : valid_1_12; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1523 = 3'h6 == state ? _GEN_1454 : valid_1_13; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1524 = 3'h6 == state ? _GEN_1455 : valid_1_14; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1525 = 3'h6 == state ? _GEN_1456 : valid_1_15; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1526 = 3'h6 == state ? _GEN_1457 : valid_2_0; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1527 = 3'h6 == state ? _GEN_1458 : valid_2_1; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1528 = 3'h6 == state ? _GEN_1459 : valid_2_2; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1529 = 3'h6 == state ? _GEN_1460 : valid_2_3; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1530 = 3'h6 == state ? _GEN_1461 : valid_2_4; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1531 = 3'h6 == state ? _GEN_1462 : valid_2_5; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1532 = 3'h6 == state ? _GEN_1463 : valid_2_6; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1533 = 3'h6 == state ? _GEN_1464 : valid_2_7; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1534 = 3'h6 == state ? _GEN_1465 : valid_2_8; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1535 = 3'h6 == state ? _GEN_1466 : valid_2_9; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1536 = 3'h6 == state ? _GEN_1467 : valid_2_10; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1537 = 3'h6 == state ? _GEN_1468 : valid_2_11; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1538 = 3'h6 == state ? _GEN_1469 : valid_2_12; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1539 = 3'h6 == state ? _GEN_1470 : valid_2_13; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1540 = 3'h6 == state ? _GEN_1471 : valid_2_14; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1541 = 3'h6 == state ? _GEN_1472 : valid_2_15; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1542 = 3'h6 == state ? _GEN_1473 : valid_3_0; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1543 = 3'h6 == state ? _GEN_1474 : valid_3_1; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1544 = 3'h6 == state ? _GEN_1475 : valid_3_2; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1545 = 3'h6 == state ? _GEN_1476 : valid_3_3; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1546 = 3'h6 == state ? _GEN_1477 : valid_3_4; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1547 = 3'h6 == state ? _GEN_1478 : valid_3_5; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1548 = 3'h6 == state ? _GEN_1479 : valid_3_6; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1549 = 3'h6 == state ? _GEN_1480 : valid_3_7; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1550 = 3'h6 == state ? _GEN_1481 : valid_3_8; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1551 = 3'h6 == state ? _GEN_1482 : valid_3_9; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1552 = 3'h6 == state ? _GEN_1483 : valid_3_10; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1553 = 3'h6 == state ? _GEN_1484 : valid_3_11; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1554 = 3'h6 == state ? _GEN_1485 : valid_3_12; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1555 = 3'h6 == state ? _GEN_1486 : valid_3_13; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1556 = 3'h6 == state ? _GEN_1487 : valid_3_14; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1557 = 3'h6 == state ? _GEN_1488 : valid_3_15; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1558 = 3'h6 == state ? _GEN_1489 : axiWaddrEn; // @[playground/src/noop/dcache.scala 205:18 199:34]
  wire [1:0] _GEN_1559 = 3'h6 == state ? _GEN_1490 : _GEN_129; // @[playground/src/noop/dcache.scala 205:18]
  wire [3:0] _GEN_1560 = 3'h6 == state ? _GEN_1491 : _GEN_133; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1563 = 3'h5 == state ? 1'h0 : wait_r; // @[playground/src/noop/dcache.scala 205:18 282:21 95:30]
  wire [2:0] _GEN_1564 = 3'h5 == state ? 3'h0 : _GEN_1493; // @[playground/src/noop/dcache.scala 205:18 283:21]
  wire  _GEN_1565 = 3'h5 == state ? _GEN_134 : _GEN_1492; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1566 = 3'h5 == state ? valid_0_0 : _GEN_1494; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1567 = 3'h5 == state ? valid_0_1 : _GEN_1495; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1568 = 3'h5 == state ? valid_0_2 : _GEN_1496; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1569 = 3'h5 == state ? valid_0_3 : _GEN_1497; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1570 = 3'h5 == state ? valid_0_4 : _GEN_1498; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1571 = 3'h5 == state ? valid_0_5 : _GEN_1499; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1572 = 3'h5 == state ? valid_0_6 : _GEN_1500; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1573 = 3'h5 == state ? valid_0_7 : _GEN_1501; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1574 = 3'h5 == state ? valid_0_8 : _GEN_1502; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1575 = 3'h5 == state ? valid_0_9 : _GEN_1503; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1576 = 3'h5 == state ? valid_0_10 : _GEN_1504; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1577 = 3'h5 == state ? valid_0_11 : _GEN_1505; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1578 = 3'h5 == state ? valid_0_12 : _GEN_1506; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1579 = 3'h5 == state ? valid_0_13 : _GEN_1507; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1580 = 3'h5 == state ? valid_0_14 : _GEN_1508; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1581 = 3'h5 == state ? valid_0_15 : _GEN_1509; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1582 = 3'h5 == state ? valid_1_0 : _GEN_1510; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1583 = 3'h5 == state ? valid_1_1 : _GEN_1511; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1584 = 3'h5 == state ? valid_1_2 : _GEN_1512; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1585 = 3'h5 == state ? valid_1_3 : _GEN_1513; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1586 = 3'h5 == state ? valid_1_4 : _GEN_1514; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1587 = 3'h5 == state ? valid_1_5 : _GEN_1515; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1588 = 3'h5 == state ? valid_1_6 : _GEN_1516; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1589 = 3'h5 == state ? valid_1_7 : _GEN_1517; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1590 = 3'h5 == state ? valid_1_8 : _GEN_1518; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1591 = 3'h5 == state ? valid_1_9 : _GEN_1519; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1592 = 3'h5 == state ? valid_1_10 : _GEN_1520; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1593 = 3'h5 == state ? valid_1_11 : _GEN_1521; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1594 = 3'h5 == state ? valid_1_12 : _GEN_1522; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1595 = 3'h5 == state ? valid_1_13 : _GEN_1523; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1596 = 3'h5 == state ? valid_1_14 : _GEN_1524; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1597 = 3'h5 == state ? valid_1_15 : _GEN_1525; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1598 = 3'h5 == state ? valid_2_0 : _GEN_1526; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1599 = 3'h5 == state ? valid_2_1 : _GEN_1527; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1600 = 3'h5 == state ? valid_2_2 : _GEN_1528; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1601 = 3'h5 == state ? valid_2_3 : _GEN_1529; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1602 = 3'h5 == state ? valid_2_4 : _GEN_1530; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1603 = 3'h5 == state ? valid_2_5 : _GEN_1531; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1604 = 3'h5 == state ? valid_2_6 : _GEN_1532; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1605 = 3'h5 == state ? valid_2_7 : _GEN_1533; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1606 = 3'h5 == state ? valid_2_8 : _GEN_1534; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1607 = 3'h5 == state ? valid_2_9 : _GEN_1535; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1608 = 3'h5 == state ? valid_2_10 : _GEN_1536; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1609 = 3'h5 == state ? valid_2_11 : _GEN_1537; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1610 = 3'h5 == state ? valid_2_12 : _GEN_1538; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1611 = 3'h5 == state ? valid_2_13 : _GEN_1539; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1612 = 3'h5 == state ? valid_2_14 : _GEN_1540; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1613 = 3'h5 == state ? valid_2_15 : _GEN_1541; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1614 = 3'h5 == state ? valid_3_0 : _GEN_1542; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1615 = 3'h5 == state ? valid_3_1 : _GEN_1543; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1616 = 3'h5 == state ? valid_3_2 : _GEN_1544; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1617 = 3'h5 == state ? valid_3_3 : _GEN_1545; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1618 = 3'h5 == state ? valid_3_4 : _GEN_1546; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1619 = 3'h5 == state ? valid_3_5 : _GEN_1547; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1620 = 3'h5 == state ? valid_3_6 : _GEN_1548; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1621 = 3'h5 == state ? valid_3_7 : _GEN_1549; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1622 = 3'h5 == state ? valid_3_8 : _GEN_1550; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1623 = 3'h5 == state ? valid_3_9 : _GEN_1551; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1624 = 3'h5 == state ? valid_3_10 : _GEN_1552; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1625 = 3'h5 == state ? valid_3_11 : _GEN_1553; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1626 = 3'h5 == state ? valid_3_12 : _GEN_1554; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1627 = 3'h5 == state ? valid_3_13 : _GEN_1555; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1628 = 3'h5 == state ? valid_3_14 : _GEN_1556; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1629 = 3'h5 == state ? valid_3_15 : _GEN_1557; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1630 = 3'h5 == state ? axiWaddrEn : _GEN_1558; // @[playground/src/noop/dcache.scala 205:18 199:34]
  wire [1:0] _GEN_1631 = 3'h5 == state ? _GEN_129 : _GEN_1559; // @[playground/src/noop/dcache.scala 205:18]
  wire [3:0] _GEN_1632 = 3'h5 == state ? _GEN_133 : _GEN_1560; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1633 = 3'h4 == state ? _GEN_1293 : axiWdataEn; // @[playground/src/noop/dcache.scala 205:18 202:34]
  wire [2:0] _GEN_1634 = 3'h4 == state ? _GEN_1292 : offset; // @[playground/src/noop/dcache.scala 205:18 110:34]
  wire [2:0] _GEN_1635 = 3'h4 == state ? _GEN_1294 : _GEN_1564; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1636 = 3'h4 == state ? _GEN_1295 : _GEN_1566; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1637 = 3'h4 == state ? _GEN_1296 : _GEN_1567; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1638 = 3'h4 == state ? _GEN_1297 : _GEN_1568; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1639 = 3'h4 == state ? _GEN_1298 : _GEN_1569; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1640 = 3'h4 == state ? _GEN_1299 : _GEN_1570; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1641 = 3'h4 == state ? _GEN_1300 : _GEN_1571; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1642 = 3'h4 == state ? _GEN_1301 : _GEN_1572; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1643 = 3'h4 == state ? _GEN_1302 : _GEN_1573; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1644 = 3'h4 == state ? _GEN_1303 : _GEN_1574; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1645 = 3'h4 == state ? _GEN_1304 : _GEN_1575; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1646 = 3'h4 == state ? _GEN_1305 : _GEN_1576; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1647 = 3'h4 == state ? _GEN_1306 : _GEN_1577; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1648 = 3'h4 == state ? _GEN_1307 : _GEN_1578; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1649 = 3'h4 == state ? _GEN_1308 : _GEN_1579; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1650 = 3'h4 == state ? _GEN_1309 : _GEN_1580; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1651 = 3'h4 == state ? _GEN_1310 : _GEN_1581; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1652 = 3'h4 == state ? _GEN_1311 : _GEN_1582; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1653 = 3'h4 == state ? _GEN_1312 : _GEN_1583; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1654 = 3'h4 == state ? _GEN_1313 : _GEN_1584; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1655 = 3'h4 == state ? _GEN_1314 : _GEN_1585; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1656 = 3'h4 == state ? _GEN_1315 : _GEN_1586; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1657 = 3'h4 == state ? _GEN_1316 : _GEN_1587; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1658 = 3'h4 == state ? _GEN_1317 : _GEN_1588; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1659 = 3'h4 == state ? _GEN_1318 : _GEN_1589; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1660 = 3'h4 == state ? _GEN_1319 : _GEN_1590; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1661 = 3'h4 == state ? _GEN_1320 : _GEN_1591; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1662 = 3'h4 == state ? _GEN_1321 : _GEN_1592; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1663 = 3'h4 == state ? _GEN_1322 : _GEN_1593; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1664 = 3'h4 == state ? _GEN_1323 : _GEN_1594; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1665 = 3'h4 == state ? _GEN_1324 : _GEN_1595; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1666 = 3'h4 == state ? _GEN_1325 : _GEN_1596; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1667 = 3'h4 == state ? _GEN_1326 : _GEN_1597; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1668 = 3'h4 == state ? _GEN_1327 : _GEN_1598; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1669 = 3'h4 == state ? _GEN_1328 : _GEN_1599; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1670 = 3'h4 == state ? _GEN_1329 : _GEN_1600; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1671 = 3'h4 == state ? _GEN_1330 : _GEN_1601; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1672 = 3'h4 == state ? _GEN_1331 : _GEN_1602; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1673 = 3'h4 == state ? _GEN_1332 : _GEN_1603; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1674 = 3'h4 == state ? _GEN_1333 : _GEN_1604; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1675 = 3'h4 == state ? _GEN_1334 : _GEN_1605; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1676 = 3'h4 == state ? _GEN_1335 : _GEN_1606; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1677 = 3'h4 == state ? _GEN_1336 : _GEN_1607; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1678 = 3'h4 == state ? _GEN_1337 : _GEN_1608; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1679 = 3'h4 == state ? _GEN_1338 : _GEN_1609; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1680 = 3'h4 == state ? _GEN_1339 : _GEN_1610; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1681 = 3'h4 == state ? _GEN_1340 : _GEN_1611; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1682 = 3'h4 == state ? _GEN_1341 : _GEN_1612; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1683 = 3'h4 == state ? _GEN_1342 : _GEN_1613; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1684 = 3'h4 == state ? _GEN_1343 : _GEN_1614; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1685 = 3'h4 == state ? _GEN_1344 : _GEN_1615; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1686 = 3'h4 == state ? _GEN_1345 : _GEN_1616; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1687 = 3'h4 == state ? _GEN_1346 : _GEN_1617; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1688 = 3'h4 == state ? _GEN_1347 : _GEN_1618; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1689 = 3'h4 == state ? _GEN_1348 : _GEN_1619; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1690 = 3'h4 == state ? _GEN_1349 : _GEN_1620; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1691 = 3'h4 == state ? _GEN_1350 : _GEN_1621; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1692 = 3'h4 == state ? _GEN_1351 : _GEN_1622; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1693 = 3'h4 == state ? _GEN_1352 : _GEN_1623; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1694 = 3'h4 == state ? _GEN_1353 : _GEN_1624; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1695 = 3'h4 == state ? _GEN_1354 : _GEN_1625; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1696 = 3'h4 == state ? _GEN_1355 : _GEN_1626; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1697 = 3'h4 == state ? _GEN_1356 : _GEN_1627; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1698 = 3'h4 == state ? _GEN_1357 : _GEN_1628; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1699 = 3'h4 == state ? _GEN_1358 : _GEN_1629; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1700 = 3'h4 == state ? _GEN_1359 : _GEN_414; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1701 = 3'h4 == state ? _GEN_1360 : _GEN_415; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1702 = 3'h4 == state ? _GEN_1361 : _GEN_416; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1703 = 3'h4 == state ? _GEN_1362 : _GEN_417; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1704 = 3'h4 == state ? _GEN_1363 : _GEN_418; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1705 = 3'h4 == state ? _GEN_1364 : _GEN_419; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1706 = 3'h4 == state ? _GEN_1365 : _GEN_420; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1707 = 3'h4 == state ? _GEN_1366 : _GEN_421; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1708 = 3'h4 == state ? _GEN_1367 : _GEN_422; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1709 = 3'h4 == state ? _GEN_1368 : _GEN_423; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1710 = 3'h4 == state ? _GEN_1369 : _GEN_424; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1711 = 3'h4 == state ? _GEN_1370 : _GEN_425; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1712 = 3'h4 == state ? _GEN_1371 : _GEN_426; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1713 = 3'h4 == state ? _GEN_1372 : _GEN_427; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1714 = 3'h4 == state ? _GEN_1373 : _GEN_428; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1715 = 3'h4 == state ? _GEN_1374 : _GEN_429; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1716 = 3'h4 == state ? _GEN_1375 : _GEN_430; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1717 = 3'h4 == state ? _GEN_1376 : _GEN_431; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1718 = 3'h4 == state ? _GEN_1377 : _GEN_432; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1719 = 3'h4 == state ? _GEN_1378 : _GEN_433; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1720 = 3'h4 == state ? _GEN_1379 : _GEN_434; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1721 = 3'h4 == state ? _GEN_1380 : _GEN_435; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1722 = 3'h4 == state ? _GEN_1381 : _GEN_436; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1723 = 3'h4 == state ? _GEN_1382 : _GEN_437; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1724 = 3'h4 == state ? _GEN_1383 : _GEN_438; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1725 = 3'h4 == state ? _GEN_1384 : _GEN_439; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1726 = 3'h4 == state ? _GEN_1385 : _GEN_440; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1727 = 3'h4 == state ? _GEN_1386 : _GEN_441; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1728 = 3'h4 == state ? _GEN_1387 : _GEN_442; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1729 = 3'h4 == state ? _GEN_1388 : _GEN_443; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1730 = 3'h4 == state ? _GEN_1389 : _GEN_444; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1731 = 3'h4 == state ? _GEN_1390 : _GEN_445; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1732 = 3'h4 == state ? _GEN_1391 : _GEN_446; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1733 = 3'h4 == state ? _GEN_1392 : _GEN_447; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1734 = 3'h4 == state ? _GEN_1393 : _GEN_448; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1735 = 3'h4 == state ? _GEN_1394 : _GEN_449; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1736 = 3'h4 == state ? _GEN_1395 : _GEN_450; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1737 = 3'h4 == state ? _GEN_1396 : _GEN_451; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1738 = 3'h4 == state ? _GEN_1397 : _GEN_452; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1739 = 3'h4 == state ? _GEN_1398 : _GEN_453; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1740 = 3'h4 == state ? _GEN_1399 : _GEN_454; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1741 = 3'h4 == state ? _GEN_1400 : _GEN_455; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1742 = 3'h4 == state ? _GEN_1401 : _GEN_456; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1743 = 3'h4 == state ? _GEN_1402 : _GEN_457; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1744 = 3'h4 == state ? _GEN_1403 : _GEN_458; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1745 = 3'h4 == state ? _GEN_1404 : _GEN_459; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1746 = 3'h4 == state ? _GEN_1405 : _GEN_460; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1747 = 3'h4 == state ? _GEN_1406 : _GEN_461; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1748 = 3'h4 == state ? _GEN_1407 : _GEN_462; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1749 = 3'h4 == state ? _GEN_1408 : _GEN_463; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1750 = 3'h4 == state ? _GEN_1409 : _GEN_464; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1751 = 3'h4 == state ? _GEN_1410 : _GEN_465; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1752 = 3'h4 == state ? _GEN_1411 : _GEN_466; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1753 = 3'h4 == state ? _GEN_1412 : _GEN_467; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1754 = 3'h4 == state ? _GEN_1413 : _GEN_468; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1755 = 3'h4 == state ? _GEN_1414 : _GEN_469; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1756 = 3'h4 == state ? _GEN_1415 : _GEN_470; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1757 = 3'h4 == state ? _GEN_1416 : _GEN_471; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1758 = 3'h4 == state ? _GEN_1417 : _GEN_472; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1759 = 3'h4 == state ? _GEN_1418 : _GEN_473; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1760 = 3'h4 == state ? _GEN_1419 : _GEN_474; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1761 = 3'h4 == state ? _GEN_1420 : _GEN_475; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1762 = 3'h4 == state ? _GEN_1421 : _GEN_476; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1763 = 3'h4 == state ? _GEN_1422 : _GEN_477; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1766 = 3'h4 == state ? wait_r : _GEN_1563; // @[playground/src/noop/dcache.scala 205:18 95:30]
  wire  _GEN_1767 = 3'h4 == state ? _GEN_134 : _GEN_1565; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1768 = 3'h4 == state ? axiWaddrEn : _GEN_1630; // @[playground/src/noop/dcache.scala 205:18 199:34]
  wire [1:0] _GEN_1769 = 3'h4 == state ? _GEN_129 : _GEN_1631; // @[playground/src/noop/dcache.scala 205:18]
  wire [3:0] _GEN_1770 = 3'h4 == state ? _GEN_133 : _GEN_1632; // @[playground/src/noop/dcache.scala 205:18]
  wire [2:0] _GEN_1771 = 3'h3 == state ? 3'h0 : _GEN_1634; // @[playground/src/noop/dcache.scala 205:18 259:20]
  wire [2:0] _GEN_1772 = 3'h3 == state ? _GEN_1031 : _GEN_1635; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1773 = 3'h3 == state ? _GEN_1032 : _GEN_1768; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1774 = 3'h3 == state ? _GEN_1033 : _GEN_1633; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1775 = 3'h3 == state ? valid_0_0 : _GEN_1636; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1776 = 3'h3 == state ? valid_0_1 : _GEN_1637; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1777 = 3'h3 == state ? valid_0_2 : _GEN_1638; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1778 = 3'h3 == state ? valid_0_3 : _GEN_1639; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1779 = 3'h3 == state ? valid_0_4 : _GEN_1640; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1780 = 3'h3 == state ? valid_0_5 : _GEN_1641; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1781 = 3'h3 == state ? valid_0_6 : _GEN_1642; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1782 = 3'h3 == state ? valid_0_7 : _GEN_1643; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1783 = 3'h3 == state ? valid_0_8 : _GEN_1644; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1784 = 3'h3 == state ? valid_0_9 : _GEN_1645; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1785 = 3'h3 == state ? valid_0_10 : _GEN_1646; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1786 = 3'h3 == state ? valid_0_11 : _GEN_1647; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1787 = 3'h3 == state ? valid_0_12 : _GEN_1648; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1788 = 3'h3 == state ? valid_0_13 : _GEN_1649; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1789 = 3'h3 == state ? valid_0_14 : _GEN_1650; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1790 = 3'h3 == state ? valid_0_15 : _GEN_1651; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1791 = 3'h3 == state ? valid_1_0 : _GEN_1652; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1792 = 3'h3 == state ? valid_1_1 : _GEN_1653; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1793 = 3'h3 == state ? valid_1_2 : _GEN_1654; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1794 = 3'h3 == state ? valid_1_3 : _GEN_1655; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1795 = 3'h3 == state ? valid_1_4 : _GEN_1656; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1796 = 3'h3 == state ? valid_1_5 : _GEN_1657; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1797 = 3'h3 == state ? valid_1_6 : _GEN_1658; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1798 = 3'h3 == state ? valid_1_7 : _GEN_1659; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1799 = 3'h3 == state ? valid_1_8 : _GEN_1660; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1800 = 3'h3 == state ? valid_1_9 : _GEN_1661; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1801 = 3'h3 == state ? valid_1_10 : _GEN_1662; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1802 = 3'h3 == state ? valid_1_11 : _GEN_1663; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1803 = 3'h3 == state ? valid_1_12 : _GEN_1664; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1804 = 3'h3 == state ? valid_1_13 : _GEN_1665; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1805 = 3'h3 == state ? valid_1_14 : _GEN_1666; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1806 = 3'h3 == state ? valid_1_15 : _GEN_1667; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1807 = 3'h3 == state ? valid_2_0 : _GEN_1668; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1808 = 3'h3 == state ? valid_2_1 : _GEN_1669; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1809 = 3'h3 == state ? valid_2_2 : _GEN_1670; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1810 = 3'h3 == state ? valid_2_3 : _GEN_1671; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1811 = 3'h3 == state ? valid_2_4 : _GEN_1672; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1812 = 3'h3 == state ? valid_2_5 : _GEN_1673; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1813 = 3'h3 == state ? valid_2_6 : _GEN_1674; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1814 = 3'h3 == state ? valid_2_7 : _GEN_1675; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1815 = 3'h3 == state ? valid_2_8 : _GEN_1676; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1816 = 3'h3 == state ? valid_2_9 : _GEN_1677; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1817 = 3'h3 == state ? valid_2_10 : _GEN_1678; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1818 = 3'h3 == state ? valid_2_11 : _GEN_1679; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1819 = 3'h3 == state ? valid_2_12 : _GEN_1680; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1820 = 3'h3 == state ? valid_2_13 : _GEN_1681; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1821 = 3'h3 == state ? valid_2_14 : _GEN_1682; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1822 = 3'h3 == state ? valid_2_15 : _GEN_1683; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1823 = 3'h3 == state ? valid_3_0 : _GEN_1684; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1824 = 3'h3 == state ? valid_3_1 : _GEN_1685; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1825 = 3'h3 == state ? valid_3_2 : _GEN_1686; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1826 = 3'h3 == state ? valid_3_3 : _GEN_1687; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1827 = 3'h3 == state ? valid_3_4 : _GEN_1688; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1828 = 3'h3 == state ? valid_3_5 : _GEN_1689; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1829 = 3'h3 == state ? valid_3_6 : _GEN_1690; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1830 = 3'h3 == state ? valid_3_7 : _GEN_1691; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1831 = 3'h3 == state ? valid_3_8 : _GEN_1692; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1832 = 3'h3 == state ? valid_3_9 : _GEN_1693; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1833 = 3'h3 == state ? valid_3_10 : _GEN_1694; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1834 = 3'h3 == state ? valid_3_11 : _GEN_1695; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1835 = 3'h3 == state ? valid_3_12 : _GEN_1696; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1836 = 3'h3 == state ? valid_3_13 : _GEN_1697; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1837 = 3'h3 == state ? valid_3_14 : _GEN_1698; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1838 = 3'h3 == state ? valid_3_15 : _GEN_1699; // @[playground/src/noop/dcache.scala 205:18 89:26]
  wire  _GEN_1839 = 3'h3 == state ? _GEN_414 : _GEN_1700; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1840 = 3'h3 == state ? _GEN_415 : _GEN_1701; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1841 = 3'h3 == state ? _GEN_416 : _GEN_1702; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1842 = 3'h3 == state ? _GEN_417 : _GEN_1703; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1843 = 3'h3 == state ? _GEN_418 : _GEN_1704; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1844 = 3'h3 == state ? _GEN_419 : _GEN_1705; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1845 = 3'h3 == state ? _GEN_420 : _GEN_1706; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1846 = 3'h3 == state ? _GEN_421 : _GEN_1707; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1847 = 3'h3 == state ? _GEN_422 : _GEN_1708; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1848 = 3'h3 == state ? _GEN_423 : _GEN_1709; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1849 = 3'h3 == state ? _GEN_424 : _GEN_1710; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1850 = 3'h3 == state ? _GEN_425 : _GEN_1711; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1851 = 3'h3 == state ? _GEN_426 : _GEN_1712; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1852 = 3'h3 == state ? _GEN_427 : _GEN_1713; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1853 = 3'h3 == state ? _GEN_428 : _GEN_1714; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1854 = 3'h3 == state ? _GEN_429 : _GEN_1715; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1855 = 3'h3 == state ? _GEN_430 : _GEN_1716; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1856 = 3'h3 == state ? _GEN_431 : _GEN_1717; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1857 = 3'h3 == state ? _GEN_432 : _GEN_1718; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1858 = 3'h3 == state ? _GEN_433 : _GEN_1719; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1859 = 3'h3 == state ? _GEN_434 : _GEN_1720; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1860 = 3'h3 == state ? _GEN_435 : _GEN_1721; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1861 = 3'h3 == state ? _GEN_436 : _GEN_1722; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1862 = 3'h3 == state ? _GEN_437 : _GEN_1723; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1863 = 3'h3 == state ? _GEN_438 : _GEN_1724; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1864 = 3'h3 == state ? _GEN_439 : _GEN_1725; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1865 = 3'h3 == state ? _GEN_440 : _GEN_1726; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1866 = 3'h3 == state ? _GEN_441 : _GEN_1727; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1867 = 3'h3 == state ? _GEN_442 : _GEN_1728; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1868 = 3'h3 == state ? _GEN_443 : _GEN_1729; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1869 = 3'h3 == state ? _GEN_444 : _GEN_1730; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1870 = 3'h3 == state ? _GEN_445 : _GEN_1731; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1871 = 3'h3 == state ? _GEN_446 : _GEN_1732; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1872 = 3'h3 == state ? _GEN_447 : _GEN_1733; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1873 = 3'h3 == state ? _GEN_448 : _GEN_1734; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1874 = 3'h3 == state ? _GEN_449 : _GEN_1735; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1875 = 3'h3 == state ? _GEN_450 : _GEN_1736; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1876 = 3'h3 == state ? _GEN_451 : _GEN_1737; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1877 = 3'h3 == state ? _GEN_452 : _GEN_1738; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1878 = 3'h3 == state ? _GEN_453 : _GEN_1739; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1879 = 3'h3 == state ? _GEN_454 : _GEN_1740; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1880 = 3'h3 == state ? _GEN_455 : _GEN_1741; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1881 = 3'h3 == state ? _GEN_456 : _GEN_1742; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1882 = 3'h3 == state ? _GEN_457 : _GEN_1743; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1883 = 3'h3 == state ? _GEN_458 : _GEN_1744; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1884 = 3'h3 == state ? _GEN_459 : _GEN_1745; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1885 = 3'h3 == state ? _GEN_460 : _GEN_1746; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1886 = 3'h3 == state ? _GEN_461 : _GEN_1747; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1887 = 3'h3 == state ? _GEN_462 : _GEN_1748; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1888 = 3'h3 == state ? _GEN_463 : _GEN_1749; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1889 = 3'h3 == state ? _GEN_464 : _GEN_1750; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1890 = 3'h3 == state ? _GEN_465 : _GEN_1751; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1891 = 3'h3 == state ? _GEN_466 : _GEN_1752; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1892 = 3'h3 == state ? _GEN_467 : _GEN_1753; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1893 = 3'h3 == state ? _GEN_468 : _GEN_1754; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1894 = 3'h3 == state ? _GEN_469 : _GEN_1755; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1895 = 3'h3 == state ? _GEN_470 : _GEN_1756; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1896 = 3'h3 == state ? _GEN_471 : _GEN_1757; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1897 = 3'h3 == state ? _GEN_472 : _GEN_1758; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1898 = 3'h3 == state ? _GEN_473 : _GEN_1759; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1899 = 3'h3 == state ? _GEN_474 : _GEN_1760; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1900 = 3'h3 == state ? _GEN_475 : _GEN_1761; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1901 = 3'h3 == state ? _GEN_476 : _GEN_1762; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1902 = 3'h3 == state ? _GEN_477 : _GEN_1763; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_1905 = 3'h3 == state ? wait_r : _GEN_1766; // @[playground/src/noop/dcache.scala 205:18 95:30]
  wire  _GEN_1906 = 3'h3 == state ? _GEN_134 : _GEN_1767; // @[playground/src/noop/dcache.scala 205:18]
  wire [1:0] _GEN_1907 = 3'h3 == state ? _GEN_129 : _GEN_1769; // @[playground/src/noop/dcache.scala 205:18]
  wire [3:0] _GEN_1908 = 3'h3 == state ? _GEN_133 : _GEN_1770; // @[playground/src/noop/dcache.scala 205:18]
  wire  _GEN_2319 = 3'h0 == state & _GEN_629; // @[playground/src/noop/dcache.scala 101:13 205:18]
  Ram_bw Ram_bw ( // @[playground/src/noop/dcache.scala 91:57]
    .clock(Ram_bw_clock),
    .reset(Ram_bw_reset),
    .io_cen(Ram_bw_io_cen),
    .io_wen(Ram_bw_io_wen),
    .io_addr(Ram_bw_io_addr),
    .io_rdata(Ram_bw_io_rdata),
    .io_wdata(Ram_bw_io_wdata),
    .io_mask(Ram_bw_io_mask)
  );
  Ram_bw Ram_bw_1 ( // @[playground/src/noop/dcache.scala 91:57]
    .clock(Ram_bw_1_clock),
    .reset(Ram_bw_1_reset),
    .io_cen(Ram_bw_1_io_cen),
    .io_wen(Ram_bw_1_io_wen),
    .io_addr(Ram_bw_1_io_addr),
    .io_rdata(Ram_bw_1_io_rdata),
    .io_wdata(Ram_bw_1_io_wdata),
    .io_mask(Ram_bw_1_io_mask)
  );
  Ram_bw Ram_bw_2 ( // @[playground/src/noop/dcache.scala 91:57]
    .clock(Ram_bw_2_clock),
    .reset(Ram_bw_2_reset),
    .io_cen(Ram_bw_2_io_cen),
    .io_wen(Ram_bw_2_io_wen),
    .io_addr(Ram_bw_2_io_addr),
    .io_rdata(Ram_bw_2_io_rdata),
    .io_wdata(Ram_bw_2_io_wdata),
    .io_mask(Ram_bw_2_io_mask)
  );
  Ram_bw Ram_bw_3 ( // @[playground/src/noop/dcache.scala 91:57]
    .clock(Ram_bw_3_clock),
    .reset(Ram_bw_3_reset),
    .io_cen(Ram_bw_3_io_cen),
    .io_wen(Ram_bw_3_io_wen),
    .io_addr(Ram_bw_3_io_addr),
    .io_rdata(Ram_bw_3_io_rdata),
    .io_wdata(Ram_bw_3_io_wdata),
    .io_mask(Ram_bw_3_io_mask)
  );
  MaxPeriodFibonacciLFSR matchWay_prng ( // @[src/main/scala/chisel3/util/random/PRNG.scala 91:22]
    .clock(matchWay_prng_clock),
    .reset(matchWay_prng_reset),
    .io_out_0(matchWay_prng_io_out_0),
    .io_out_1(matchWay_prng_io_out_1)
  );
  assign io_dataAxi_wa_valid = axiWaddrEn; // @[playground/src/noop/dcache.scala 308:30]
  assign io_dataAxi_wa_bits_addr = {axiWaddr_hi,6'h0}; // @[playground/src/noop/dcache.scala 200:30]
  assign io_dataAxi_wd_valid = axiWdataEn; // @[playground/src/noop/dcache.scala 314:30]
  assign io_dataAxi_wd_bits_data = offset[0] ? _GEN_329[127:64] : _GEN_329[63:0]; // @[playground/src/noop/dcache.scala 201:30]
  assign io_dataAxi_wd_bits_last = offset == 3'h7; // @[playground/src/noop/dcache.scala 203:34]
  assign io_dataAxi_ra_valid = axiRaddrEn; // @[playground/src/noop/dcache.scala 300:30]
  assign io_dataAxi_ra_bits_addr = cur_addr & 32'hffffffc0; // @[playground/src/noop/dcache.scala 197:36]
  assign io_dcRW_rdata = _io_dcRW_rdata_T_40[63:0]; // @[playground/src/noop/dcache.scala 154:19]
  assign io_dcRW_rvalid = valid_r; // @[playground/src/noop/dcache.scala 105:20]
  assign io_dcRW_ready = valid_in & ~wait_r; // @[playground/src/noop/dcache.scala 104:31]
  assign io_flush_out = flush_r; // @[playground/src/noop/dcache.scala 106:18]
  assign Ram_bw_clock = clock;
  assign Ram_bw_reset = reset;
  assign Ram_bw_io_cen = 2'h0 == _GEN_129 & (wait_r | hs_in | flush_r); // @[playground/src/noop/dcache.scala 184:{25,25} playground/src/ram/ram.scala 41:17]
  assign Ram_bw_io_wen = _GEN_2524 & wen; // @[playground/src/noop/dcache.scala 185:{25,25} playground/src/ram/ram.scala 42:17]
  assign Ram_bw_io_addr = 2'h0 == _GEN_129 ? _data_addr_T_3 : 6'h0; // @[playground/src/noop/dcache.scala 183:{25,25} playground/src/ram/ram.scala 43:17]
  assign Ram_bw_io_wdata = 2'h0 == _GEN_129 ? _data_wdata_T_4[127:0] : 128'h0; // @[playground/src/noop/dcache.scala 186:{25,25} playground/src/ram/ram.scala 44:17]
  assign Ram_bw_io_mask = 2'h0 == _GEN_129 ? mask : 128'h0; // @[playground/src/noop/dcache.scala 188:{25,25} playground/src/ram/ram.scala 45:17]
  assign Ram_bw_1_clock = clock;
  assign Ram_bw_1_reset = reset;
  assign Ram_bw_1_io_cen = 2'h1 == _GEN_129 & (wait_r | hs_in | flush_r); // @[playground/src/noop/dcache.scala 184:{25,25} playground/src/ram/ram.scala 41:17]
  assign Ram_bw_1_io_wen = _GEN_2525 & wen; // @[playground/src/noop/dcache.scala 185:{25,25} playground/src/ram/ram.scala 42:17]
  assign Ram_bw_1_io_addr = 2'h1 == _GEN_129 ? _data_addr_T_3 : 6'h0; // @[playground/src/noop/dcache.scala 183:{25,25} playground/src/ram/ram.scala 43:17]
  assign Ram_bw_1_io_wdata = 2'h1 == _GEN_129 ? _data_wdata_T_4[127:0] : 128'h0; // @[playground/src/noop/dcache.scala 186:{25,25} playground/src/ram/ram.scala 44:17]
  assign Ram_bw_1_io_mask = 2'h1 == _GEN_129 ? mask : 128'h0; // @[playground/src/noop/dcache.scala 188:{25,25} playground/src/ram/ram.scala 45:17]
  assign Ram_bw_2_clock = clock;
  assign Ram_bw_2_reset = reset;
  assign Ram_bw_2_io_cen = 2'h2 == _GEN_129 & (wait_r | hs_in | flush_r); // @[playground/src/noop/dcache.scala 184:{25,25} playground/src/ram/ram.scala 41:17]
  assign Ram_bw_2_io_wen = _GEN_2526 & wen; // @[playground/src/noop/dcache.scala 185:{25,25} playground/src/ram/ram.scala 42:17]
  assign Ram_bw_2_io_addr = 2'h2 == _GEN_129 ? _data_addr_T_3 : 6'h0; // @[playground/src/noop/dcache.scala 183:{25,25} playground/src/ram/ram.scala 43:17]
  assign Ram_bw_2_io_wdata = 2'h2 == _GEN_129 ? _data_wdata_T_4[127:0] : 128'h0; // @[playground/src/noop/dcache.scala 186:{25,25} playground/src/ram/ram.scala 44:17]
  assign Ram_bw_2_io_mask = 2'h2 == _GEN_129 ? mask : 128'h0; // @[playground/src/noop/dcache.scala 188:{25,25} playground/src/ram/ram.scala 45:17]
  assign Ram_bw_3_clock = clock;
  assign Ram_bw_3_reset = reset;
  assign Ram_bw_3_io_cen = 2'h3 == _GEN_129 & (wait_r | hs_in | flush_r); // @[playground/src/noop/dcache.scala 184:{25,25} playground/src/ram/ram.scala 41:17]
  assign Ram_bw_3_io_wen = _GEN_2527 & wen; // @[playground/src/noop/dcache.scala 185:{25,25} playground/src/ram/ram.scala 42:17]
  assign Ram_bw_3_io_addr = 2'h3 == _GEN_129 ? _data_addr_T_3 : 6'h0; // @[playground/src/noop/dcache.scala 183:{25,25} playground/src/ram/ram.scala 43:17]
  assign Ram_bw_3_io_wdata = 2'h3 == _GEN_129 ? _data_wdata_T_4[127:0] : 128'h0; // @[playground/src/noop/dcache.scala 186:{25,25} playground/src/ram/ram.scala 44:17]
  assign Ram_bw_3_io_mask = 2'h3 == _GEN_129 ? mask : 128'h0; // @[playground/src/noop/dcache.scala 188:{25,25} playground/src/ram/ram.scala 45:17]
  assign matchWay_prng_clock = clock;
  assign matchWay_prng_reset = reset;
  always @(posedge clock) begin
    if (reset) begin // @[playground/src/noop/dcache.scala 88:26]
      tag_0_0 <= 22'h0; // @[playground/src/noop/dcache.scala 88:26]
    end else if (!(3'h0 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
      if (!(3'h1 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
        if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
          tag_0_0 <= _GEN_902;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 88:26]
      tag_0_1 <= 22'h0; // @[playground/src/noop/dcache.scala 88:26]
    end else if (!(3'h0 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
      if (!(3'h1 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
        if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
          tag_0_1 <= _GEN_903;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 88:26]
      tag_0_2 <= 22'h0; // @[playground/src/noop/dcache.scala 88:26]
    end else if (!(3'h0 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
      if (!(3'h1 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
        if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
          tag_0_2 <= _GEN_904;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 88:26]
      tag_0_3 <= 22'h0; // @[playground/src/noop/dcache.scala 88:26]
    end else if (!(3'h0 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
      if (!(3'h1 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
        if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
          tag_0_3 <= _GEN_905;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 88:26]
      tag_0_4 <= 22'h0; // @[playground/src/noop/dcache.scala 88:26]
    end else if (!(3'h0 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
      if (!(3'h1 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
        if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
          tag_0_4 <= _GEN_906;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 88:26]
      tag_0_5 <= 22'h0; // @[playground/src/noop/dcache.scala 88:26]
    end else if (!(3'h0 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
      if (!(3'h1 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
        if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
          tag_0_5 <= _GEN_907;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 88:26]
      tag_0_6 <= 22'h0; // @[playground/src/noop/dcache.scala 88:26]
    end else if (!(3'h0 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
      if (!(3'h1 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
        if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
          tag_0_6 <= _GEN_908;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 88:26]
      tag_0_7 <= 22'h0; // @[playground/src/noop/dcache.scala 88:26]
    end else if (!(3'h0 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
      if (!(3'h1 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
        if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
          tag_0_7 <= _GEN_909;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 88:26]
      tag_0_8 <= 22'h0; // @[playground/src/noop/dcache.scala 88:26]
    end else if (!(3'h0 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
      if (!(3'h1 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
        if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
          tag_0_8 <= _GEN_910;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 88:26]
      tag_0_9 <= 22'h0; // @[playground/src/noop/dcache.scala 88:26]
    end else if (!(3'h0 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
      if (!(3'h1 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
        if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
          tag_0_9 <= _GEN_911;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 88:26]
      tag_0_10 <= 22'h0; // @[playground/src/noop/dcache.scala 88:26]
    end else if (!(3'h0 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
      if (!(3'h1 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
        if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
          tag_0_10 <= _GEN_912;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 88:26]
      tag_0_11 <= 22'h0; // @[playground/src/noop/dcache.scala 88:26]
    end else if (!(3'h0 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
      if (!(3'h1 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
        if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
          tag_0_11 <= _GEN_913;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 88:26]
      tag_0_12 <= 22'h0; // @[playground/src/noop/dcache.scala 88:26]
    end else if (!(3'h0 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
      if (!(3'h1 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
        if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
          tag_0_12 <= _GEN_914;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 88:26]
      tag_0_13 <= 22'h0; // @[playground/src/noop/dcache.scala 88:26]
    end else if (!(3'h0 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
      if (!(3'h1 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
        if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
          tag_0_13 <= _GEN_915;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 88:26]
      tag_0_14 <= 22'h0; // @[playground/src/noop/dcache.scala 88:26]
    end else if (!(3'h0 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
      if (!(3'h1 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
        if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
          tag_0_14 <= _GEN_916;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 88:26]
      tag_0_15 <= 22'h0; // @[playground/src/noop/dcache.scala 88:26]
    end else if (!(3'h0 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
      if (!(3'h1 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
        if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
          tag_0_15 <= _GEN_917;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 88:26]
      tag_1_0 <= 22'h0; // @[playground/src/noop/dcache.scala 88:26]
    end else if (!(3'h0 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
      if (!(3'h1 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
        if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
          tag_1_0 <= _GEN_918;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 88:26]
      tag_1_1 <= 22'h0; // @[playground/src/noop/dcache.scala 88:26]
    end else if (!(3'h0 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
      if (!(3'h1 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
        if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
          tag_1_1 <= _GEN_919;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 88:26]
      tag_1_2 <= 22'h0; // @[playground/src/noop/dcache.scala 88:26]
    end else if (!(3'h0 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
      if (!(3'h1 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
        if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
          tag_1_2 <= _GEN_920;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 88:26]
      tag_1_3 <= 22'h0; // @[playground/src/noop/dcache.scala 88:26]
    end else if (!(3'h0 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
      if (!(3'h1 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
        if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
          tag_1_3 <= _GEN_921;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 88:26]
      tag_1_4 <= 22'h0; // @[playground/src/noop/dcache.scala 88:26]
    end else if (!(3'h0 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
      if (!(3'h1 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
        if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
          tag_1_4 <= _GEN_922;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 88:26]
      tag_1_5 <= 22'h0; // @[playground/src/noop/dcache.scala 88:26]
    end else if (!(3'h0 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
      if (!(3'h1 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
        if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
          tag_1_5 <= _GEN_923;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 88:26]
      tag_1_6 <= 22'h0; // @[playground/src/noop/dcache.scala 88:26]
    end else if (!(3'h0 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
      if (!(3'h1 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
        if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
          tag_1_6 <= _GEN_924;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 88:26]
      tag_1_7 <= 22'h0; // @[playground/src/noop/dcache.scala 88:26]
    end else if (!(3'h0 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
      if (!(3'h1 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
        if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
          tag_1_7 <= _GEN_925;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 88:26]
      tag_1_8 <= 22'h0; // @[playground/src/noop/dcache.scala 88:26]
    end else if (!(3'h0 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
      if (!(3'h1 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
        if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
          tag_1_8 <= _GEN_926;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 88:26]
      tag_1_9 <= 22'h0; // @[playground/src/noop/dcache.scala 88:26]
    end else if (!(3'h0 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
      if (!(3'h1 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
        if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
          tag_1_9 <= _GEN_927;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 88:26]
      tag_1_10 <= 22'h0; // @[playground/src/noop/dcache.scala 88:26]
    end else if (!(3'h0 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
      if (!(3'h1 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
        if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
          tag_1_10 <= _GEN_928;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 88:26]
      tag_1_11 <= 22'h0; // @[playground/src/noop/dcache.scala 88:26]
    end else if (!(3'h0 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
      if (!(3'h1 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
        if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
          tag_1_11 <= _GEN_929;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 88:26]
      tag_1_12 <= 22'h0; // @[playground/src/noop/dcache.scala 88:26]
    end else if (!(3'h0 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
      if (!(3'h1 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
        if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
          tag_1_12 <= _GEN_930;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 88:26]
      tag_1_13 <= 22'h0; // @[playground/src/noop/dcache.scala 88:26]
    end else if (!(3'h0 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
      if (!(3'h1 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
        if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
          tag_1_13 <= _GEN_931;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 88:26]
      tag_1_14 <= 22'h0; // @[playground/src/noop/dcache.scala 88:26]
    end else if (!(3'h0 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
      if (!(3'h1 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
        if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
          tag_1_14 <= _GEN_932;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 88:26]
      tag_1_15 <= 22'h0; // @[playground/src/noop/dcache.scala 88:26]
    end else if (!(3'h0 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
      if (!(3'h1 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
        if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
          tag_1_15 <= _GEN_933;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 88:26]
      tag_2_0 <= 22'h0; // @[playground/src/noop/dcache.scala 88:26]
    end else if (!(3'h0 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
      if (!(3'h1 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
        if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
          tag_2_0 <= _GEN_934;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 88:26]
      tag_2_1 <= 22'h0; // @[playground/src/noop/dcache.scala 88:26]
    end else if (!(3'h0 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
      if (!(3'h1 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
        if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
          tag_2_1 <= _GEN_935;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 88:26]
      tag_2_2 <= 22'h0; // @[playground/src/noop/dcache.scala 88:26]
    end else if (!(3'h0 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
      if (!(3'h1 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
        if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
          tag_2_2 <= _GEN_936;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 88:26]
      tag_2_3 <= 22'h0; // @[playground/src/noop/dcache.scala 88:26]
    end else if (!(3'h0 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
      if (!(3'h1 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
        if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
          tag_2_3 <= _GEN_937;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 88:26]
      tag_2_4 <= 22'h0; // @[playground/src/noop/dcache.scala 88:26]
    end else if (!(3'h0 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
      if (!(3'h1 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
        if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
          tag_2_4 <= _GEN_938;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 88:26]
      tag_2_5 <= 22'h0; // @[playground/src/noop/dcache.scala 88:26]
    end else if (!(3'h0 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
      if (!(3'h1 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
        if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
          tag_2_5 <= _GEN_939;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 88:26]
      tag_2_6 <= 22'h0; // @[playground/src/noop/dcache.scala 88:26]
    end else if (!(3'h0 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
      if (!(3'h1 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
        if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
          tag_2_6 <= _GEN_940;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 88:26]
      tag_2_7 <= 22'h0; // @[playground/src/noop/dcache.scala 88:26]
    end else if (!(3'h0 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
      if (!(3'h1 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
        if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
          tag_2_7 <= _GEN_941;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 88:26]
      tag_2_8 <= 22'h0; // @[playground/src/noop/dcache.scala 88:26]
    end else if (!(3'h0 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
      if (!(3'h1 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
        if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
          tag_2_8 <= _GEN_942;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 88:26]
      tag_2_9 <= 22'h0; // @[playground/src/noop/dcache.scala 88:26]
    end else if (!(3'h0 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
      if (!(3'h1 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
        if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
          tag_2_9 <= _GEN_943;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 88:26]
      tag_2_10 <= 22'h0; // @[playground/src/noop/dcache.scala 88:26]
    end else if (!(3'h0 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
      if (!(3'h1 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
        if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
          tag_2_10 <= _GEN_944;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 88:26]
      tag_2_11 <= 22'h0; // @[playground/src/noop/dcache.scala 88:26]
    end else if (!(3'h0 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
      if (!(3'h1 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
        if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
          tag_2_11 <= _GEN_945;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 88:26]
      tag_2_12 <= 22'h0; // @[playground/src/noop/dcache.scala 88:26]
    end else if (!(3'h0 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
      if (!(3'h1 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
        if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
          tag_2_12 <= _GEN_946;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 88:26]
      tag_2_13 <= 22'h0; // @[playground/src/noop/dcache.scala 88:26]
    end else if (!(3'h0 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
      if (!(3'h1 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
        if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
          tag_2_13 <= _GEN_947;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 88:26]
      tag_2_14 <= 22'h0; // @[playground/src/noop/dcache.scala 88:26]
    end else if (!(3'h0 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
      if (!(3'h1 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
        if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
          tag_2_14 <= _GEN_948;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 88:26]
      tag_2_15 <= 22'h0; // @[playground/src/noop/dcache.scala 88:26]
    end else if (!(3'h0 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
      if (!(3'h1 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
        if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
          tag_2_15 <= _GEN_949;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 88:26]
      tag_3_0 <= 22'h0; // @[playground/src/noop/dcache.scala 88:26]
    end else if (!(3'h0 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
      if (!(3'h1 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
        if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
          tag_3_0 <= _GEN_950;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 88:26]
      tag_3_1 <= 22'h0; // @[playground/src/noop/dcache.scala 88:26]
    end else if (!(3'h0 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
      if (!(3'h1 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
        if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
          tag_3_1 <= _GEN_951;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 88:26]
      tag_3_2 <= 22'h0; // @[playground/src/noop/dcache.scala 88:26]
    end else if (!(3'h0 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
      if (!(3'h1 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
        if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
          tag_3_2 <= _GEN_952;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 88:26]
      tag_3_3 <= 22'h0; // @[playground/src/noop/dcache.scala 88:26]
    end else if (!(3'h0 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
      if (!(3'h1 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
        if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
          tag_3_3 <= _GEN_953;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 88:26]
      tag_3_4 <= 22'h0; // @[playground/src/noop/dcache.scala 88:26]
    end else if (!(3'h0 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
      if (!(3'h1 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
        if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
          tag_3_4 <= _GEN_954;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 88:26]
      tag_3_5 <= 22'h0; // @[playground/src/noop/dcache.scala 88:26]
    end else if (!(3'h0 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
      if (!(3'h1 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
        if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
          tag_3_5 <= _GEN_955;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 88:26]
      tag_3_6 <= 22'h0; // @[playground/src/noop/dcache.scala 88:26]
    end else if (!(3'h0 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
      if (!(3'h1 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
        if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
          tag_3_6 <= _GEN_956;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 88:26]
      tag_3_7 <= 22'h0; // @[playground/src/noop/dcache.scala 88:26]
    end else if (!(3'h0 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
      if (!(3'h1 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
        if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
          tag_3_7 <= _GEN_957;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 88:26]
      tag_3_8 <= 22'h0; // @[playground/src/noop/dcache.scala 88:26]
    end else if (!(3'h0 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
      if (!(3'h1 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
        if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
          tag_3_8 <= _GEN_958;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 88:26]
      tag_3_9 <= 22'h0; // @[playground/src/noop/dcache.scala 88:26]
    end else if (!(3'h0 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
      if (!(3'h1 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
        if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
          tag_3_9 <= _GEN_959;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 88:26]
      tag_3_10 <= 22'h0; // @[playground/src/noop/dcache.scala 88:26]
    end else if (!(3'h0 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
      if (!(3'h1 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
        if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
          tag_3_10 <= _GEN_960;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 88:26]
      tag_3_11 <= 22'h0; // @[playground/src/noop/dcache.scala 88:26]
    end else if (!(3'h0 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
      if (!(3'h1 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
        if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
          tag_3_11 <= _GEN_961;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 88:26]
      tag_3_12 <= 22'h0; // @[playground/src/noop/dcache.scala 88:26]
    end else if (!(3'h0 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
      if (!(3'h1 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
        if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
          tag_3_12 <= _GEN_962;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 88:26]
      tag_3_13 <= 22'h0; // @[playground/src/noop/dcache.scala 88:26]
    end else if (!(3'h0 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
      if (!(3'h1 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
        if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
          tag_3_13 <= _GEN_963;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 88:26]
      tag_3_14 <= 22'h0; // @[playground/src/noop/dcache.scala 88:26]
    end else if (!(3'h0 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
      if (!(3'h1 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
        if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
          tag_3_14 <= _GEN_964;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 88:26]
      tag_3_15 <= 22'h0; // @[playground/src/noop/dcache.scala 88:26]
    end else if (!(3'h0 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
      if (!(3'h1 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
        if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
          tag_3_15 <= _GEN_965;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 89:26]
      valid_0_0 <= 1'h0; // @[playground/src/noop/dcache.scala 89:26]
    end else if (!(3'h0 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
      if (!(3'h1 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
        if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
          valid_0_0 <= _GEN_966;
        end else begin
          valid_0_0 <= _GEN_1775;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 89:26]
      valid_0_1 <= 1'h0; // @[playground/src/noop/dcache.scala 89:26]
    end else if (!(3'h0 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
      if (!(3'h1 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
        if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
          valid_0_1 <= _GEN_967;
        end else begin
          valid_0_1 <= _GEN_1776;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 89:26]
      valid_0_2 <= 1'h0; // @[playground/src/noop/dcache.scala 89:26]
    end else if (!(3'h0 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
      if (!(3'h1 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
        if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
          valid_0_2 <= _GEN_968;
        end else begin
          valid_0_2 <= _GEN_1777;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 89:26]
      valid_0_3 <= 1'h0; // @[playground/src/noop/dcache.scala 89:26]
    end else if (!(3'h0 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
      if (!(3'h1 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
        if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
          valid_0_3 <= _GEN_969;
        end else begin
          valid_0_3 <= _GEN_1778;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 89:26]
      valid_0_4 <= 1'h0; // @[playground/src/noop/dcache.scala 89:26]
    end else if (!(3'h0 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
      if (!(3'h1 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
        if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
          valid_0_4 <= _GEN_970;
        end else begin
          valid_0_4 <= _GEN_1779;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 89:26]
      valid_0_5 <= 1'h0; // @[playground/src/noop/dcache.scala 89:26]
    end else if (!(3'h0 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
      if (!(3'h1 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
        if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
          valid_0_5 <= _GEN_971;
        end else begin
          valid_0_5 <= _GEN_1780;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 89:26]
      valid_0_6 <= 1'h0; // @[playground/src/noop/dcache.scala 89:26]
    end else if (!(3'h0 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
      if (!(3'h1 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
        if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
          valid_0_6 <= _GEN_972;
        end else begin
          valid_0_6 <= _GEN_1781;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 89:26]
      valid_0_7 <= 1'h0; // @[playground/src/noop/dcache.scala 89:26]
    end else if (!(3'h0 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
      if (!(3'h1 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
        if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
          valid_0_7 <= _GEN_973;
        end else begin
          valid_0_7 <= _GEN_1782;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 89:26]
      valid_0_8 <= 1'h0; // @[playground/src/noop/dcache.scala 89:26]
    end else if (!(3'h0 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
      if (!(3'h1 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
        if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
          valid_0_8 <= _GEN_974;
        end else begin
          valid_0_8 <= _GEN_1783;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 89:26]
      valid_0_9 <= 1'h0; // @[playground/src/noop/dcache.scala 89:26]
    end else if (!(3'h0 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
      if (!(3'h1 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
        if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
          valid_0_9 <= _GEN_975;
        end else begin
          valid_0_9 <= _GEN_1784;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 89:26]
      valid_0_10 <= 1'h0; // @[playground/src/noop/dcache.scala 89:26]
    end else if (!(3'h0 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
      if (!(3'h1 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
        if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
          valid_0_10 <= _GEN_976;
        end else begin
          valid_0_10 <= _GEN_1785;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 89:26]
      valid_0_11 <= 1'h0; // @[playground/src/noop/dcache.scala 89:26]
    end else if (!(3'h0 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
      if (!(3'h1 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
        if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
          valid_0_11 <= _GEN_977;
        end else begin
          valid_0_11 <= _GEN_1786;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 89:26]
      valid_0_12 <= 1'h0; // @[playground/src/noop/dcache.scala 89:26]
    end else if (!(3'h0 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
      if (!(3'h1 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
        if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
          valid_0_12 <= _GEN_978;
        end else begin
          valid_0_12 <= _GEN_1787;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 89:26]
      valid_0_13 <= 1'h0; // @[playground/src/noop/dcache.scala 89:26]
    end else if (!(3'h0 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
      if (!(3'h1 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
        if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
          valid_0_13 <= _GEN_979;
        end else begin
          valid_0_13 <= _GEN_1788;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 89:26]
      valid_0_14 <= 1'h0; // @[playground/src/noop/dcache.scala 89:26]
    end else if (!(3'h0 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
      if (!(3'h1 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
        if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
          valid_0_14 <= _GEN_980;
        end else begin
          valid_0_14 <= _GEN_1789;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 89:26]
      valid_0_15 <= 1'h0; // @[playground/src/noop/dcache.scala 89:26]
    end else if (!(3'h0 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
      if (!(3'h1 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
        if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
          valid_0_15 <= _GEN_981;
        end else begin
          valid_0_15 <= _GEN_1790;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 89:26]
      valid_1_0 <= 1'h0; // @[playground/src/noop/dcache.scala 89:26]
    end else if (!(3'h0 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
      if (!(3'h1 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
        if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
          valid_1_0 <= _GEN_982;
        end else begin
          valid_1_0 <= _GEN_1791;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 89:26]
      valid_1_1 <= 1'h0; // @[playground/src/noop/dcache.scala 89:26]
    end else if (!(3'h0 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
      if (!(3'h1 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
        if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
          valid_1_1 <= _GEN_983;
        end else begin
          valid_1_1 <= _GEN_1792;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 89:26]
      valid_1_2 <= 1'h0; // @[playground/src/noop/dcache.scala 89:26]
    end else if (!(3'h0 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
      if (!(3'h1 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
        if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
          valid_1_2 <= _GEN_984;
        end else begin
          valid_1_2 <= _GEN_1793;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 89:26]
      valid_1_3 <= 1'h0; // @[playground/src/noop/dcache.scala 89:26]
    end else if (!(3'h0 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
      if (!(3'h1 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
        if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
          valid_1_3 <= _GEN_985;
        end else begin
          valid_1_3 <= _GEN_1794;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 89:26]
      valid_1_4 <= 1'h0; // @[playground/src/noop/dcache.scala 89:26]
    end else if (!(3'h0 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
      if (!(3'h1 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
        if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
          valid_1_4 <= _GEN_986;
        end else begin
          valid_1_4 <= _GEN_1795;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 89:26]
      valid_1_5 <= 1'h0; // @[playground/src/noop/dcache.scala 89:26]
    end else if (!(3'h0 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
      if (!(3'h1 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
        if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
          valid_1_5 <= _GEN_987;
        end else begin
          valid_1_5 <= _GEN_1796;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 89:26]
      valid_1_6 <= 1'h0; // @[playground/src/noop/dcache.scala 89:26]
    end else if (!(3'h0 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
      if (!(3'h1 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
        if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
          valid_1_6 <= _GEN_988;
        end else begin
          valid_1_6 <= _GEN_1797;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 89:26]
      valid_1_7 <= 1'h0; // @[playground/src/noop/dcache.scala 89:26]
    end else if (!(3'h0 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
      if (!(3'h1 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
        if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
          valid_1_7 <= _GEN_989;
        end else begin
          valid_1_7 <= _GEN_1798;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 89:26]
      valid_1_8 <= 1'h0; // @[playground/src/noop/dcache.scala 89:26]
    end else if (!(3'h0 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
      if (!(3'h1 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
        if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
          valid_1_8 <= _GEN_990;
        end else begin
          valid_1_8 <= _GEN_1799;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 89:26]
      valid_1_9 <= 1'h0; // @[playground/src/noop/dcache.scala 89:26]
    end else if (!(3'h0 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
      if (!(3'h1 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
        if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
          valid_1_9 <= _GEN_991;
        end else begin
          valid_1_9 <= _GEN_1800;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 89:26]
      valid_1_10 <= 1'h0; // @[playground/src/noop/dcache.scala 89:26]
    end else if (!(3'h0 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
      if (!(3'h1 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
        if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
          valid_1_10 <= _GEN_992;
        end else begin
          valid_1_10 <= _GEN_1801;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 89:26]
      valid_1_11 <= 1'h0; // @[playground/src/noop/dcache.scala 89:26]
    end else if (!(3'h0 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
      if (!(3'h1 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
        if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
          valid_1_11 <= _GEN_993;
        end else begin
          valid_1_11 <= _GEN_1802;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 89:26]
      valid_1_12 <= 1'h0; // @[playground/src/noop/dcache.scala 89:26]
    end else if (!(3'h0 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
      if (!(3'h1 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
        if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
          valid_1_12 <= _GEN_994;
        end else begin
          valid_1_12 <= _GEN_1803;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 89:26]
      valid_1_13 <= 1'h0; // @[playground/src/noop/dcache.scala 89:26]
    end else if (!(3'h0 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
      if (!(3'h1 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
        if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
          valid_1_13 <= _GEN_995;
        end else begin
          valid_1_13 <= _GEN_1804;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 89:26]
      valid_1_14 <= 1'h0; // @[playground/src/noop/dcache.scala 89:26]
    end else if (!(3'h0 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
      if (!(3'h1 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
        if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
          valid_1_14 <= _GEN_996;
        end else begin
          valid_1_14 <= _GEN_1805;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 89:26]
      valid_1_15 <= 1'h0; // @[playground/src/noop/dcache.scala 89:26]
    end else if (!(3'h0 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
      if (!(3'h1 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
        if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
          valid_1_15 <= _GEN_997;
        end else begin
          valid_1_15 <= _GEN_1806;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 89:26]
      valid_2_0 <= 1'h0; // @[playground/src/noop/dcache.scala 89:26]
    end else if (!(3'h0 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
      if (!(3'h1 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
        if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
          valid_2_0 <= _GEN_998;
        end else begin
          valid_2_0 <= _GEN_1807;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 89:26]
      valid_2_1 <= 1'h0; // @[playground/src/noop/dcache.scala 89:26]
    end else if (!(3'h0 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
      if (!(3'h1 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
        if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
          valid_2_1 <= _GEN_999;
        end else begin
          valid_2_1 <= _GEN_1808;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 89:26]
      valid_2_2 <= 1'h0; // @[playground/src/noop/dcache.scala 89:26]
    end else if (!(3'h0 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
      if (!(3'h1 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
        if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
          valid_2_2 <= _GEN_1000;
        end else begin
          valid_2_2 <= _GEN_1809;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 89:26]
      valid_2_3 <= 1'h0; // @[playground/src/noop/dcache.scala 89:26]
    end else if (!(3'h0 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
      if (!(3'h1 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
        if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
          valid_2_3 <= _GEN_1001;
        end else begin
          valid_2_3 <= _GEN_1810;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 89:26]
      valid_2_4 <= 1'h0; // @[playground/src/noop/dcache.scala 89:26]
    end else if (!(3'h0 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
      if (!(3'h1 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
        if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
          valid_2_4 <= _GEN_1002;
        end else begin
          valid_2_4 <= _GEN_1811;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 89:26]
      valid_2_5 <= 1'h0; // @[playground/src/noop/dcache.scala 89:26]
    end else if (!(3'h0 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
      if (!(3'h1 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
        if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
          valid_2_5 <= _GEN_1003;
        end else begin
          valid_2_5 <= _GEN_1812;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 89:26]
      valid_2_6 <= 1'h0; // @[playground/src/noop/dcache.scala 89:26]
    end else if (!(3'h0 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
      if (!(3'h1 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
        if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
          valid_2_6 <= _GEN_1004;
        end else begin
          valid_2_6 <= _GEN_1813;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 89:26]
      valid_2_7 <= 1'h0; // @[playground/src/noop/dcache.scala 89:26]
    end else if (!(3'h0 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
      if (!(3'h1 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
        if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
          valid_2_7 <= _GEN_1005;
        end else begin
          valid_2_7 <= _GEN_1814;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 89:26]
      valid_2_8 <= 1'h0; // @[playground/src/noop/dcache.scala 89:26]
    end else if (!(3'h0 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
      if (!(3'h1 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
        if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
          valid_2_8 <= _GEN_1006;
        end else begin
          valid_2_8 <= _GEN_1815;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 89:26]
      valid_2_9 <= 1'h0; // @[playground/src/noop/dcache.scala 89:26]
    end else if (!(3'h0 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
      if (!(3'h1 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
        if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
          valid_2_9 <= _GEN_1007;
        end else begin
          valid_2_9 <= _GEN_1816;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 89:26]
      valid_2_10 <= 1'h0; // @[playground/src/noop/dcache.scala 89:26]
    end else if (!(3'h0 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
      if (!(3'h1 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
        if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
          valid_2_10 <= _GEN_1008;
        end else begin
          valid_2_10 <= _GEN_1817;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 89:26]
      valid_2_11 <= 1'h0; // @[playground/src/noop/dcache.scala 89:26]
    end else if (!(3'h0 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
      if (!(3'h1 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
        if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
          valid_2_11 <= _GEN_1009;
        end else begin
          valid_2_11 <= _GEN_1818;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 89:26]
      valid_2_12 <= 1'h0; // @[playground/src/noop/dcache.scala 89:26]
    end else if (!(3'h0 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
      if (!(3'h1 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
        if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
          valid_2_12 <= _GEN_1010;
        end else begin
          valid_2_12 <= _GEN_1819;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 89:26]
      valid_2_13 <= 1'h0; // @[playground/src/noop/dcache.scala 89:26]
    end else if (!(3'h0 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
      if (!(3'h1 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
        if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
          valid_2_13 <= _GEN_1011;
        end else begin
          valid_2_13 <= _GEN_1820;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 89:26]
      valid_2_14 <= 1'h0; // @[playground/src/noop/dcache.scala 89:26]
    end else if (!(3'h0 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
      if (!(3'h1 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
        if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
          valid_2_14 <= _GEN_1012;
        end else begin
          valid_2_14 <= _GEN_1821;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 89:26]
      valid_2_15 <= 1'h0; // @[playground/src/noop/dcache.scala 89:26]
    end else if (!(3'h0 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
      if (!(3'h1 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
        if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
          valid_2_15 <= _GEN_1013;
        end else begin
          valid_2_15 <= _GEN_1822;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 89:26]
      valid_3_0 <= 1'h0; // @[playground/src/noop/dcache.scala 89:26]
    end else if (!(3'h0 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
      if (!(3'h1 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
        if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
          valid_3_0 <= _GEN_1014;
        end else begin
          valid_3_0 <= _GEN_1823;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 89:26]
      valid_3_1 <= 1'h0; // @[playground/src/noop/dcache.scala 89:26]
    end else if (!(3'h0 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
      if (!(3'h1 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
        if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
          valid_3_1 <= _GEN_1015;
        end else begin
          valid_3_1 <= _GEN_1824;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 89:26]
      valid_3_2 <= 1'h0; // @[playground/src/noop/dcache.scala 89:26]
    end else if (!(3'h0 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
      if (!(3'h1 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
        if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
          valid_3_2 <= _GEN_1016;
        end else begin
          valid_3_2 <= _GEN_1825;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 89:26]
      valid_3_3 <= 1'h0; // @[playground/src/noop/dcache.scala 89:26]
    end else if (!(3'h0 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
      if (!(3'h1 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
        if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
          valid_3_3 <= _GEN_1017;
        end else begin
          valid_3_3 <= _GEN_1826;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 89:26]
      valid_3_4 <= 1'h0; // @[playground/src/noop/dcache.scala 89:26]
    end else if (!(3'h0 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
      if (!(3'h1 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
        if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
          valid_3_4 <= _GEN_1018;
        end else begin
          valid_3_4 <= _GEN_1827;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 89:26]
      valid_3_5 <= 1'h0; // @[playground/src/noop/dcache.scala 89:26]
    end else if (!(3'h0 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
      if (!(3'h1 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
        if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
          valid_3_5 <= _GEN_1019;
        end else begin
          valid_3_5 <= _GEN_1828;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 89:26]
      valid_3_6 <= 1'h0; // @[playground/src/noop/dcache.scala 89:26]
    end else if (!(3'h0 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
      if (!(3'h1 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
        if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
          valid_3_6 <= _GEN_1020;
        end else begin
          valid_3_6 <= _GEN_1829;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 89:26]
      valid_3_7 <= 1'h0; // @[playground/src/noop/dcache.scala 89:26]
    end else if (!(3'h0 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
      if (!(3'h1 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
        if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
          valid_3_7 <= _GEN_1021;
        end else begin
          valid_3_7 <= _GEN_1830;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 89:26]
      valid_3_8 <= 1'h0; // @[playground/src/noop/dcache.scala 89:26]
    end else if (!(3'h0 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
      if (!(3'h1 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
        if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
          valid_3_8 <= _GEN_1022;
        end else begin
          valid_3_8 <= _GEN_1831;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 89:26]
      valid_3_9 <= 1'h0; // @[playground/src/noop/dcache.scala 89:26]
    end else if (!(3'h0 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
      if (!(3'h1 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
        if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
          valid_3_9 <= _GEN_1023;
        end else begin
          valid_3_9 <= _GEN_1832;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 89:26]
      valid_3_10 <= 1'h0; // @[playground/src/noop/dcache.scala 89:26]
    end else if (!(3'h0 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
      if (!(3'h1 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
        if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
          valid_3_10 <= _GEN_1024;
        end else begin
          valid_3_10 <= _GEN_1833;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 89:26]
      valid_3_11 <= 1'h0; // @[playground/src/noop/dcache.scala 89:26]
    end else if (!(3'h0 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
      if (!(3'h1 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
        if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
          valid_3_11 <= _GEN_1025;
        end else begin
          valid_3_11 <= _GEN_1834;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 89:26]
      valid_3_12 <= 1'h0; // @[playground/src/noop/dcache.scala 89:26]
    end else if (!(3'h0 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
      if (!(3'h1 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
        if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
          valid_3_12 <= _GEN_1026;
        end else begin
          valid_3_12 <= _GEN_1835;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 89:26]
      valid_3_13 <= 1'h0; // @[playground/src/noop/dcache.scala 89:26]
    end else if (!(3'h0 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
      if (!(3'h1 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
        if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
          valid_3_13 <= _GEN_1027;
        end else begin
          valid_3_13 <= _GEN_1836;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 89:26]
      valid_3_14 <= 1'h0; // @[playground/src/noop/dcache.scala 89:26]
    end else if (!(3'h0 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
      if (!(3'h1 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
        if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
          valid_3_14 <= _GEN_1028;
        end else begin
          valid_3_14 <= _GEN_1837;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 89:26]
      valid_3_15 <= 1'h0; // @[playground/src/noop/dcache.scala 89:26]
    end else if (!(3'h0 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
      if (!(3'h1 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
        if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
          valid_3_15 <= _GEN_1029;
        end else begin
          valid_3_15 <= _GEN_1838;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 90:26]
      dirty_0_0 <= 1'h0; // @[playground/src/noop/dcache.scala 90:26]
    end else if (3'h0 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_0_0 <= _GEN_414;
    end else if (3'h1 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_0_0 <= _GEN_414;
    end else if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_0_0 <= _GEN_414;
    end else begin
      dirty_0_0 <= _GEN_1839;
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 90:26]
      dirty_0_1 <= 1'h0; // @[playground/src/noop/dcache.scala 90:26]
    end else if (3'h0 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_0_1 <= _GEN_415;
    end else if (3'h1 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_0_1 <= _GEN_415;
    end else if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_0_1 <= _GEN_415;
    end else begin
      dirty_0_1 <= _GEN_1840;
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 90:26]
      dirty_0_2 <= 1'h0; // @[playground/src/noop/dcache.scala 90:26]
    end else if (3'h0 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_0_2 <= _GEN_416;
    end else if (3'h1 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_0_2 <= _GEN_416;
    end else if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_0_2 <= _GEN_416;
    end else begin
      dirty_0_2 <= _GEN_1841;
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 90:26]
      dirty_0_3 <= 1'h0; // @[playground/src/noop/dcache.scala 90:26]
    end else if (3'h0 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_0_3 <= _GEN_417;
    end else if (3'h1 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_0_3 <= _GEN_417;
    end else if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_0_3 <= _GEN_417;
    end else begin
      dirty_0_3 <= _GEN_1842;
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 90:26]
      dirty_0_4 <= 1'h0; // @[playground/src/noop/dcache.scala 90:26]
    end else if (3'h0 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_0_4 <= _GEN_418;
    end else if (3'h1 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_0_4 <= _GEN_418;
    end else if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_0_4 <= _GEN_418;
    end else begin
      dirty_0_4 <= _GEN_1843;
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 90:26]
      dirty_0_5 <= 1'h0; // @[playground/src/noop/dcache.scala 90:26]
    end else if (3'h0 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_0_5 <= _GEN_419;
    end else if (3'h1 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_0_5 <= _GEN_419;
    end else if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_0_5 <= _GEN_419;
    end else begin
      dirty_0_5 <= _GEN_1844;
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 90:26]
      dirty_0_6 <= 1'h0; // @[playground/src/noop/dcache.scala 90:26]
    end else if (3'h0 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_0_6 <= _GEN_420;
    end else if (3'h1 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_0_6 <= _GEN_420;
    end else if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_0_6 <= _GEN_420;
    end else begin
      dirty_0_6 <= _GEN_1845;
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 90:26]
      dirty_0_7 <= 1'h0; // @[playground/src/noop/dcache.scala 90:26]
    end else if (3'h0 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_0_7 <= _GEN_421;
    end else if (3'h1 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_0_7 <= _GEN_421;
    end else if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_0_7 <= _GEN_421;
    end else begin
      dirty_0_7 <= _GEN_1846;
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 90:26]
      dirty_0_8 <= 1'h0; // @[playground/src/noop/dcache.scala 90:26]
    end else if (3'h0 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_0_8 <= _GEN_422;
    end else if (3'h1 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_0_8 <= _GEN_422;
    end else if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_0_8 <= _GEN_422;
    end else begin
      dirty_0_8 <= _GEN_1847;
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 90:26]
      dirty_0_9 <= 1'h0; // @[playground/src/noop/dcache.scala 90:26]
    end else if (3'h0 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_0_9 <= _GEN_423;
    end else if (3'h1 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_0_9 <= _GEN_423;
    end else if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_0_9 <= _GEN_423;
    end else begin
      dirty_0_9 <= _GEN_1848;
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 90:26]
      dirty_0_10 <= 1'h0; // @[playground/src/noop/dcache.scala 90:26]
    end else if (3'h0 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_0_10 <= _GEN_424;
    end else if (3'h1 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_0_10 <= _GEN_424;
    end else if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_0_10 <= _GEN_424;
    end else begin
      dirty_0_10 <= _GEN_1849;
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 90:26]
      dirty_0_11 <= 1'h0; // @[playground/src/noop/dcache.scala 90:26]
    end else if (3'h0 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_0_11 <= _GEN_425;
    end else if (3'h1 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_0_11 <= _GEN_425;
    end else if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_0_11 <= _GEN_425;
    end else begin
      dirty_0_11 <= _GEN_1850;
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 90:26]
      dirty_0_12 <= 1'h0; // @[playground/src/noop/dcache.scala 90:26]
    end else if (3'h0 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_0_12 <= _GEN_426;
    end else if (3'h1 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_0_12 <= _GEN_426;
    end else if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_0_12 <= _GEN_426;
    end else begin
      dirty_0_12 <= _GEN_1851;
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 90:26]
      dirty_0_13 <= 1'h0; // @[playground/src/noop/dcache.scala 90:26]
    end else if (3'h0 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_0_13 <= _GEN_427;
    end else if (3'h1 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_0_13 <= _GEN_427;
    end else if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_0_13 <= _GEN_427;
    end else begin
      dirty_0_13 <= _GEN_1852;
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 90:26]
      dirty_0_14 <= 1'h0; // @[playground/src/noop/dcache.scala 90:26]
    end else if (3'h0 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_0_14 <= _GEN_428;
    end else if (3'h1 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_0_14 <= _GEN_428;
    end else if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_0_14 <= _GEN_428;
    end else begin
      dirty_0_14 <= _GEN_1853;
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 90:26]
      dirty_0_15 <= 1'h0; // @[playground/src/noop/dcache.scala 90:26]
    end else if (3'h0 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_0_15 <= _GEN_429;
    end else if (3'h1 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_0_15 <= _GEN_429;
    end else if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_0_15 <= _GEN_429;
    end else begin
      dirty_0_15 <= _GEN_1854;
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 90:26]
      dirty_1_0 <= 1'h0; // @[playground/src/noop/dcache.scala 90:26]
    end else if (3'h0 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_1_0 <= _GEN_430;
    end else if (3'h1 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_1_0 <= _GEN_430;
    end else if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_1_0 <= _GEN_430;
    end else begin
      dirty_1_0 <= _GEN_1855;
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 90:26]
      dirty_1_1 <= 1'h0; // @[playground/src/noop/dcache.scala 90:26]
    end else if (3'h0 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_1_1 <= _GEN_431;
    end else if (3'h1 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_1_1 <= _GEN_431;
    end else if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_1_1 <= _GEN_431;
    end else begin
      dirty_1_1 <= _GEN_1856;
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 90:26]
      dirty_1_2 <= 1'h0; // @[playground/src/noop/dcache.scala 90:26]
    end else if (3'h0 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_1_2 <= _GEN_432;
    end else if (3'h1 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_1_2 <= _GEN_432;
    end else if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_1_2 <= _GEN_432;
    end else begin
      dirty_1_2 <= _GEN_1857;
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 90:26]
      dirty_1_3 <= 1'h0; // @[playground/src/noop/dcache.scala 90:26]
    end else if (3'h0 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_1_3 <= _GEN_433;
    end else if (3'h1 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_1_3 <= _GEN_433;
    end else if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_1_3 <= _GEN_433;
    end else begin
      dirty_1_3 <= _GEN_1858;
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 90:26]
      dirty_1_4 <= 1'h0; // @[playground/src/noop/dcache.scala 90:26]
    end else if (3'h0 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_1_4 <= _GEN_434;
    end else if (3'h1 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_1_4 <= _GEN_434;
    end else if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_1_4 <= _GEN_434;
    end else begin
      dirty_1_4 <= _GEN_1859;
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 90:26]
      dirty_1_5 <= 1'h0; // @[playground/src/noop/dcache.scala 90:26]
    end else if (3'h0 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_1_5 <= _GEN_435;
    end else if (3'h1 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_1_5 <= _GEN_435;
    end else if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_1_5 <= _GEN_435;
    end else begin
      dirty_1_5 <= _GEN_1860;
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 90:26]
      dirty_1_6 <= 1'h0; // @[playground/src/noop/dcache.scala 90:26]
    end else if (3'h0 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_1_6 <= _GEN_436;
    end else if (3'h1 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_1_6 <= _GEN_436;
    end else if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_1_6 <= _GEN_436;
    end else begin
      dirty_1_6 <= _GEN_1861;
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 90:26]
      dirty_1_7 <= 1'h0; // @[playground/src/noop/dcache.scala 90:26]
    end else if (3'h0 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_1_7 <= _GEN_437;
    end else if (3'h1 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_1_7 <= _GEN_437;
    end else if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_1_7 <= _GEN_437;
    end else begin
      dirty_1_7 <= _GEN_1862;
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 90:26]
      dirty_1_8 <= 1'h0; // @[playground/src/noop/dcache.scala 90:26]
    end else if (3'h0 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_1_8 <= _GEN_438;
    end else if (3'h1 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_1_8 <= _GEN_438;
    end else if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_1_8 <= _GEN_438;
    end else begin
      dirty_1_8 <= _GEN_1863;
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 90:26]
      dirty_1_9 <= 1'h0; // @[playground/src/noop/dcache.scala 90:26]
    end else if (3'h0 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_1_9 <= _GEN_439;
    end else if (3'h1 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_1_9 <= _GEN_439;
    end else if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_1_9 <= _GEN_439;
    end else begin
      dirty_1_9 <= _GEN_1864;
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 90:26]
      dirty_1_10 <= 1'h0; // @[playground/src/noop/dcache.scala 90:26]
    end else if (3'h0 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_1_10 <= _GEN_440;
    end else if (3'h1 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_1_10 <= _GEN_440;
    end else if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_1_10 <= _GEN_440;
    end else begin
      dirty_1_10 <= _GEN_1865;
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 90:26]
      dirty_1_11 <= 1'h0; // @[playground/src/noop/dcache.scala 90:26]
    end else if (3'h0 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_1_11 <= _GEN_441;
    end else if (3'h1 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_1_11 <= _GEN_441;
    end else if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_1_11 <= _GEN_441;
    end else begin
      dirty_1_11 <= _GEN_1866;
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 90:26]
      dirty_1_12 <= 1'h0; // @[playground/src/noop/dcache.scala 90:26]
    end else if (3'h0 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_1_12 <= _GEN_442;
    end else if (3'h1 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_1_12 <= _GEN_442;
    end else if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_1_12 <= _GEN_442;
    end else begin
      dirty_1_12 <= _GEN_1867;
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 90:26]
      dirty_1_13 <= 1'h0; // @[playground/src/noop/dcache.scala 90:26]
    end else if (3'h0 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_1_13 <= _GEN_443;
    end else if (3'h1 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_1_13 <= _GEN_443;
    end else if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_1_13 <= _GEN_443;
    end else begin
      dirty_1_13 <= _GEN_1868;
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 90:26]
      dirty_1_14 <= 1'h0; // @[playground/src/noop/dcache.scala 90:26]
    end else if (3'h0 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_1_14 <= _GEN_444;
    end else if (3'h1 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_1_14 <= _GEN_444;
    end else if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_1_14 <= _GEN_444;
    end else begin
      dirty_1_14 <= _GEN_1869;
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 90:26]
      dirty_1_15 <= 1'h0; // @[playground/src/noop/dcache.scala 90:26]
    end else if (3'h0 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_1_15 <= _GEN_445;
    end else if (3'h1 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_1_15 <= _GEN_445;
    end else if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_1_15 <= _GEN_445;
    end else begin
      dirty_1_15 <= _GEN_1870;
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 90:26]
      dirty_2_0 <= 1'h0; // @[playground/src/noop/dcache.scala 90:26]
    end else if (3'h0 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_2_0 <= _GEN_446;
    end else if (3'h1 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_2_0 <= _GEN_446;
    end else if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_2_0 <= _GEN_446;
    end else begin
      dirty_2_0 <= _GEN_1871;
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 90:26]
      dirty_2_1 <= 1'h0; // @[playground/src/noop/dcache.scala 90:26]
    end else if (3'h0 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_2_1 <= _GEN_447;
    end else if (3'h1 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_2_1 <= _GEN_447;
    end else if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_2_1 <= _GEN_447;
    end else begin
      dirty_2_1 <= _GEN_1872;
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 90:26]
      dirty_2_2 <= 1'h0; // @[playground/src/noop/dcache.scala 90:26]
    end else if (3'h0 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_2_2 <= _GEN_448;
    end else if (3'h1 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_2_2 <= _GEN_448;
    end else if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_2_2 <= _GEN_448;
    end else begin
      dirty_2_2 <= _GEN_1873;
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 90:26]
      dirty_2_3 <= 1'h0; // @[playground/src/noop/dcache.scala 90:26]
    end else if (3'h0 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_2_3 <= _GEN_449;
    end else if (3'h1 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_2_3 <= _GEN_449;
    end else if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_2_3 <= _GEN_449;
    end else begin
      dirty_2_3 <= _GEN_1874;
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 90:26]
      dirty_2_4 <= 1'h0; // @[playground/src/noop/dcache.scala 90:26]
    end else if (3'h0 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_2_4 <= _GEN_450;
    end else if (3'h1 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_2_4 <= _GEN_450;
    end else if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_2_4 <= _GEN_450;
    end else begin
      dirty_2_4 <= _GEN_1875;
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 90:26]
      dirty_2_5 <= 1'h0; // @[playground/src/noop/dcache.scala 90:26]
    end else if (3'h0 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_2_5 <= _GEN_451;
    end else if (3'h1 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_2_5 <= _GEN_451;
    end else if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_2_5 <= _GEN_451;
    end else begin
      dirty_2_5 <= _GEN_1876;
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 90:26]
      dirty_2_6 <= 1'h0; // @[playground/src/noop/dcache.scala 90:26]
    end else if (3'h0 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_2_6 <= _GEN_452;
    end else if (3'h1 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_2_6 <= _GEN_452;
    end else if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_2_6 <= _GEN_452;
    end else begin
      dirty_2_6 <= _GEN_1877;
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 90:26]
      dirty_2_7 <= 1'h0; // @[playground/src/noop/dcache.scala 90:26]
    end else if (3'h0 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_2_7 <= _GEN_453;
    end else if (3'h1 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_2_7 <= _GEN_453;
    end else if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_2_7 <= _GEN_453;
    end else begin
      dirty_2_7 <= _GEN_1878;
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 90:26]
      dirty_2_8 <= 1'h0; // @[playground/src/noop/dcache.scala 90:26]
    end else if (3'h0 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_2_8 <= _GEN_454;
    end else if (3'h1 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_2_8 <= _GEN_454;
    end else if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_2_8 <= _GEN_454;
    end else begin
      dirty_2_8 <= _GEN_1879;
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 90:26]
      dirty_2_9 <= 1'h0; // @[playground/src/noop/dcache.scala 90:26]
    end else if (3'h0 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_2_9 <= _GEN_455;
    end else if (3'h1 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_2_9 <= _GEN_455;
    end else if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_2_9 <= _GEN_455;
    end else begin
      dirty_2_9 <= _GEN_1880;
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 90:26]
      dirty_2_10 <= 1'h0; // @[playground/src/noop/dcache.scala 90:26]
    end else if (3'h0 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_2_10 <= _GEN_456;
    end else if (3'h1 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_2_10 <= _GEN_456;
    end else if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_2_10 <= _GEN_456;
    end else begin
      dirty_2_10 <= _GEN_1881;
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 90:26]
      dirty_2_11 <= 1'h0; // @[playground/src/noop/dcache.scala 90:26]
    end else if (3'h0 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_2_11 <= _GEN_457;
    end else if (3'h1 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_2_11 <= _GEN_457;
    end else if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_2_11 <= _GEN_457;
    end else begin
      dirty_2_11 <= _GEN_1882;
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 90:26]
      dirty_2_12 <= 1'h0; // @[playground/src/noop/dcache.scala 90:26]
    end else if (3'h0 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_2_12 <= _GEN_458;
    end else if (3'h1 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_2_12 <= _GEN_458;
    end else if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_2_12 <= _GEN_458;
    end else begin
      dirty_2_12 <= _GEN_1883;
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 90:26]
      dirty_2_13 <= 1'h0; // @[playground/src/noop/dcache.scala 90:26]
    end else if (3'h0 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_2_13 <= _GEN_459;
    end else if (3'h1 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_2_13 <= _GEN_459;
    end else if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_2_13 <= _GEN_459;
    end else begin
      dirty_2_13 <= _GEN_1884;
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 90:26]
      dirty_2_14 <= 1'h0; // @[playground/src/noop/dcache.scala 90:26]
    end else if (3'h0 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_2_14 <= _GEN_460;
    end else if (3'h1 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_2_14 <= _GEN_460;
    end else if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_2_14 <= _GEN_460;
    end else begin
      dirty_2_14 <= _GEN_1885;
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 90:26]
      dirty_2_15 <= 1'h0; // @[playground/src/noop/dcache.scala 90:26]
    end else if (3'h0 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_2_15 <= _GEN_461;
    end else if (3'h1 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_2_15 <= _GEN_461;
    end else if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_2_15 <= _GEN_461;
    end else begin
      dirty_2_15 <= _GEN_1886;
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 90:26]
      dirty_3_0 <= 1'h0; // @[playground/src/noop/dcache.scala 90:26]
    end else if (3'h0 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_3_0 <= _GEN_462;
    end else if (3'h1 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_3_0 <= _GEN_462;
    end else if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_3_0 <= _GEN_462;
    end else begin
      dirty_3_0 <= _GEN_1887;
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 90:26]
      dirty_3_1 <= 1'h0; // @[playground/src/noop/dcache.scala 90:26]
    end else if (3'h0 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_3_1 <= _GEN_463;
    end else if (3'h1 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_3_1 <= _GEN_463;
    end else if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_3_1 <= _GEN_463;
    end else begin
      dirty_3_1 <= _GEN_1888;
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 90:26]
      dirty_3_2 <= 1'h0; // @[playground/src/noop/dcache.scala 90:26]
    end else if (3'h0 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_3_2 <= _GEN_464;
    end else if (3'h1 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_3_2 <= _GEN_464;
    end else if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_3_2 <= _GEN_464;
    end else begin
      dirty_3_2 <= _GEN_1889;
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 90:26]
      dirty_3_3 <= 1'h0; // @[playground/src/noop/dcache.scala 90:26]
    end else if (3'h0 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_3_3 <= _GEN_465;
    end else if (3'h1 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_3_3 <= _GEN_465;
    end else if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_3_3 <= _GEN_465;
    end else begin
      dirty_3_3 <= _GEN_1890;
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 90:26]
      dirty_3_4 <= 1'h0; // @[playground/src/noop/dcache.scala 90:26]
    end else if (3'h0 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_3_4 <= _GEN_466;
    end else if (3'h1 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_3_4 <= _GEN_466;
    end else if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_3_4 <= _GEN_466;
    end else begin
      dirty_3_4 <= _GEN_1891;
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 90:26]
      dirty_3_5 <= 1'h0; // @[playground/src/noop/dcache.scala 90:26]
    end else if (3'h0 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_3_5 <= _GEN_467;
    end else if (3'h1 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_3_5 <= _GEN_467;
    end else if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_3_5 <= _GEN_467;
    end else begin
      dirty_3_5 <= _GEN_1892;
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 90:26]
      dirty_3_6 <= 1'h0; // @[playground/src/noop/dcache.scala 90:26]
    end else if (3'h0 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_3_6 <= _GEN_468;
    end else if (3'h1 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_3_6 <= _GEN_468;
    end else if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_3_6 <= _GEN_468;
    end else begin
      dirty_3_6 <= _GEN_1893;
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 90:26]
      dirty_3_7 <= 1'h0; // @[playground/src/noop/dcache.scala 90:26]
    end else if (3'h0 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_3_7 <= _GEN_469;
    end else if (3'h1 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_3_7 <= _GEN_469;
    end else if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_3_7 <= _GEN_469;
    end else begin
      dirty_3_7 <= _GEN_1894;
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 90:26]
      dirty_3_8 <= 1'h0; // @[playground/src/noop/dcache.scala 90:26]
    end else if (3'h0 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_3_8 <= _GEN_470;
    end else if (3'h1 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_3_8 <= _GEN_470;
    end else if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_3_8 <= _GEN_470;
    end else begin
      dirty_3_8 <= _GEN_1895;
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 90:26]
      dirty_3_9 <= 1'h0; // @[playground/src/noop/dcache.scala 90:26]
    end else if (3'h0 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_3_9 <= _GEN_471;
    end else if (3'h1 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_3_9 <= _GEN_471;
    end else if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_3_9 <= _GEN_471;
    end else begin
      dirty_3_9 <= _GEN_1896;
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 90:26]
      dirty_3_10 <= 1'h0; // @[playground/src/noop/dcache.scala 90:26]
    end else if (3'h0 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_3_10 <= _GEN_472;
    end else if (3'h1 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_3_10 <= _GEN_472;
    end else if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_3_10 <= _GEN_472;
    end else begin
      dirty_3_10 <= _GEN_1897;
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 90:26]
      dirty_3_11 <= 1'h0; // @[playground/src/noop/dcache.scala 90:26]
    end else if (3'h0 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_3_11 <= _GEN_473;
    end else if (3'h1 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_3_11 <= _GEN_473;
    end else if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_3_11 <= _GEN_473;
    end else begin
      dirty_3_11 <= _GEN_1898;
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 90:26]
      dirty_3_12 <= 1'h0; // @[playground/src/noop/dcache.scala 90:26]
    end else if (3'h0 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_3_12 <= _GEN_474;
    end else if (3'h1 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_3_12 <= _GEN_474;
    end else if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_3_12 <= _GEN_474;
    end else begin
      dirty_3_12 <= _GEN_1899;
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 90:26]
      dirty_3_13 <= 1'h0; // @[playground/src/noop/dcache.scala 90:26]
    end else if (3'h0 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_3_13 <= _GEN_475;
    end else if (3'h1 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_3_13 <= _GEN_475;
    end else if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_3_13 <= _GEN_475;
    end else begin
      dirty_3_13 <= _GEN_1900;
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 90:26]
      dirty_3_14 <= 1'h0; // @[playground/src/noop/dcache.scala 90:26]
    end else if (3'h0 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_3_14 <= _GEN_476;
    end else if (3'h1 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_3_14 <= _GEN_476;
    end else if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_3_14 <= _GEN_476;
    end else begin
      dirty_3_14 <= _GEN_1901;
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 90:26]
      dirty_3_15 <= 1'h0; // @[playground/src/noop/dcache.scala 90:26]
    end else if (3'h0 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_3_15 <= _GEN_477;
    end else if (3'h1 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_3_15 <= _GEN_477;
    end else if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      dirty_3_15 <= _GEN_477;
    end else begin
      dirty_3_15 <= _GEN_1902;
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 95:30]
      wait_r <= 1'h0; // @[playground/src/noop/dcache.scala 95:30]
    end else if (3'h0 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      if (!(flush_r | io_flush)) begin // @[playground/src/noop/dcache.scala 207:38]
        if (!(~hs_in & _io_dcRW_ready_T)) begin // @[playground/src/noop/dcache.scala 209:42]
          wait_r <= _GEN_616;
        end
      end
    end else if (!(3'h1 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
      if (!(3'h2 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
        wait_r <= _GEN_1905;
      end
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 96:30]
      valid_r <= 1'h0; // @[playground/src/noop/dcache.scala 96:30]
    end else begin
      valid_r <= _GEN_2319;
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 97:30]
      flush_r <= 1'h0; // @[playground/src/noop/dcache.scala 97:30]
    end else if (3'h0 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      flush_r <= _GEN_134;
    end else if (3'h1 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      flush_r <= _GEN_134;
    end else if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      flush_r <= _GEN_134;
    end else begin
      flush_r <= _GEN_1906;
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 98:30]
      mode_r <= 5'h0; // @[playground/src/noop/dcache.scala 98:30]
    end else if (hs_in) begin // @[playground/src/noop/dcache.scala 119:16]
      mode_r <= io_dcRW_dc_mode; // @[playground/src/noop/dcache.scala 122:17]
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 99:30]
      wdata_r <= 64'h0; // @[playground/src/noop/dcache.scala 99:30]
    end else if (hs_in) begin // @[playground/src/noop/dcache.scala 119:16]
      wdata_r <= io_dcRW_wdata; // @[playground/src/noop/dcache.scala 123:17]
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 100:30]
      amo_r <= 5'h0; // @[playground/src/noop/dcache.scala 100:30]
    end else if (hs_in) begin // @[playground/src/noop/dcache.scala 119:16]
      amo_r <= io_dcRW_amo; // @[playground/src/noop/dcache.scala 124:17]
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 107:34]
      addr_r <= 32'h0; // @[playground/src/noop/dcache.scala 107:34]
    end else if (hs_in) begin // @[playground/src/noop/dcache.scala 108:30]
      addr_r <= io_dcRW_addr;
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 109:34]
      matchWay_r <= 2'h0; // @[playground/src/noop/dcache.scala 109:34]
    end else if (3'h0 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      matchWay_r <= _GEN_129;
    end else if (3'h1 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      matchWay_r <= _GEN_129;
    end else if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      matchWay_r <= _GEN_129;
    end else begin
      matchWay_r <= _GEN_1907;
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 110:34]
      offset <= 3'h0; // @[playground/src/noop/dcache.scala 110:34]
    end else if (!(3'h0 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
      if (3'h1 == state) begin // @[playground/src/noop/dcache.scala 205:18]
        offset <= 3'h0; // @[playground/src/noop/dcache.scala 235:20]
      end else if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
        offset <= _GEN_898;
      end else begin
        offset <= _GEN_1771;
      end
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 111:34]
      rdatabuf <= 64'h0; // @[playground/src/noop/dcache.scala 111:34]
    end else if (!(3'h0 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
      if (!(3'h1 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
        if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
          rdatabuf <= _GEN_900;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 113:34]
      blockIdx_r <= 4'h0; // @[playground/src/noop/dcache.scala 113:34]
    end else if (3'h0 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      blockIdx_r <= _GEN_133;
    end else if (3'h1 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      blockIdx_r <= _GEN_133;
    end else if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      blockIdx_r <= _GEN_133;
    end else begin
      blockIdx_r <= _GEN_1908;
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 152:24]
      state <= 3'h0; // @[playground/src/noop/dcache.scala 152:24]
    end else if (3'h0 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      if (flush_r | io_flush) begin // @[playground/src/noop/dcache.scala 207:38]
        state <= 3'h6; // @[playground/src/noop/dcache.scala 208:23]
      end else if (!(~hs_in & _io_dcRW_ready_T)) begin // @[playground/src/noop/dcache.scala 209:42]
        state <= _GEN_614;
      end
    end else if (3'h1 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      if (axiRaddrEn & io_dataAxi_ra_ready) begin // @[playground/src/noop/dcache.scala 236:52]
        state <= 3'h2; // @[playground/src/noop/dcache.scala 237:25]
      end
    end else if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      state <= _GEN_1030;
    end else begin
      state <= _GEN_1772;
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 198:34]
      axiRdataEn <= 1'h0; // @[playground/src/noop/dcache.scala 198:34]
    end else if (!(3'h0 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
      if (3'h1 == state) begin // @[playground/src/noop/dcache.scala 205:18]
        axiRdataEn <= _GEN_637;
      end else if (3'h2 == state) begin // @[playground/src/noop/dcache.scala 205:18]
        axiRdataEn <= _GEN_901;
      end
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 196:34]
      axiRaddrEn <= 1'h0; // @[playground/src/noop/dcache.scala 196:34]
    end else if (3'h0 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      if (!(flush_r | io_flush)) begin // @[playground/src/noop/dcache.scala 207:38]
        if (!(~hs_in & _io_dcRW_ready_T)) begin // @[playground/src/noop/dcache.scala 209:42]
          axiRaddrEn <= _GEN_620;
        end
      end
    end else if (3'h1 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      if (axiRaddrEn & io_dataAxi_ra_ready) begin // @[playground/src/noop/dcache.scala 236:52]
        axiRaddrEn <= 1'h0; // @[playground/src/noop/dcache.scala 238:28]
      end
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 199:34]
      axiWaddrEn <= 1'h0; // @[playground/src/noop/dcache.scala 199:34]
    end else if (3'h0 == state) begin // @[playground/src/noop/dcache.scala 205:18]
      if (!(flush_r | io_flush)) begin // @[playground/src/noop/dcache.scala 207:38]
        if (!(~hs_in & _io_dcRW_ready_T)) begin // @[playground/src/noop/dcache.scala 209:42]
          axiWaddrEn <= _GEN_619;
        end
      end
    end else if (!(3'h1 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
      if (!(3'h2 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
        axiWaddrEn <= _GEN_1773;
      end
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 202:34]
      axiWdataEn <= 1'h0; // @[playground/src/noop/dcache.scala 202:34]
    end else if (!(3'h0 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
      if (!(3'h1 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
        if (!(3'h2 == state)) begin // @[playground/src/noop/dcache.scala 205:18]
          axiWdataEn <= _GEN_1774;
        end
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  tag_0_0 = _RAND_0[21:0];
  _RAND_1 = {1{`RANDOM}};
  tag_0_1 = _RAND_1[21:0];
  _RAND_2 = {1{`RANDOM}};
  tag_0_2 = _RAND_2[21:0];
  _RAND_3 = {1{`RANDOM}};
  tag_0_3 = _RAND_3[21:0];
  _RAND_4 = {1{`RANDOM}};
  tag_0_4 = _RAND_4[21:0];
  _RAND_5 = {1{`RANDOM}};
  tag_0_5 = _RAND_5[21:0];
  _RAND_6 = {1{`RANDOM}};
  tag_0_6 = _RAND_6[21:0];
  _RAND_7 = {1{`RANDOM}};
  tag_0_7 = _RAND_7[21:0];
  _RAND_8 = {1{`RANDOM}};
  tag_0_8 = _RAND_8[21:0];
  _RAND_9 = {1{`RANDOM}};
  tag_0_9 = _RAND_9[21:0];
  _RAND_10 = {1{`RANDOM}};
  tag_0_10 = _RAND_10[21:0];
  _RAND_11 = {1{`RANDOM}};
  tag_0_11 = _RAND_11[21:0];
  _RAND_12 = {1{`RANDOM}};
  tag_0_12 = _RAND_12[21:0];
  _RAND_13 = {1{`RANDOM}};
  tag_0_13 = _RAND_13[21:0];
  _RAND_14 = {1{`RANDOM}};
  tag_0_14 = _RAND_14[21:0];
  _RAND_15 = {1{`RANDOM}};
  tag_0_15 = _RAND_15[21:0];
  _RAND_16 = {1{`RANDOM}};
  tag_1_0 = _RAND_16[21:0];
  _RAND_17 = {1{`RANDOM}};
  tag_1_1 = _RAND_17[21:0];
  _RAND_18 = {1{`RANDOM}};
  tag_1_2 = _RAND_18[21:0];
  _RAND_19 = {1{`RANDOM}};
  tag_1_3 = _RAND_19[21:0];
  _RAND_20 = {1{`RANDOM}};
  tag_1_4 = _RAND_20[21:0];
  _RAND_21 = {1{`RANDOM}};
  tag_1_5 = _RAND_21[21:0];
  _RAND_22 = {1{`RANDOM}};
  tag_1_6 = _RAND_22[21:0];
  _RAND_23 = {1{`RANDOM}};
  tag_1_7 = _RAND_23[21:0];
  _RAND_24 = {1{`RANDOM}};
  tag_1_8 = _RAND_24[21:0];
  _RAND_25 = {1{`RANDOM}};
  tag_1_9 = _RAND_25[21:0];
  _RAND_26 = {1{`RANDOM}};
  tag_1_10 = _RAND_26[21:0];
  _RAND_27 = {1{`RANDOM}};
  tag_1_11 = _RAND_27[21:0];
  _RAND_28 = {1{`RANDOM}};
  tag_1_12 = _RAND_28[21:0];
  _RAND_29 = {1{`RANDOM}};
  tag_1_13 = _RAND_29[21:0];
  _RAND_30 = {1{`RANDOM}};
  tag_1_14 = _RAND_30[21:0];
  _RAND_31 = {1{`RANDOM}};
  tag_1_15 = _RAND_31[21:0];
  _RAND_32 = {1{`RANDOM}};
  tag_2_0 = _RAND_32[21:0];
  _RAND_33 = {1{`RANDOM}};
  tag_2_1 = _RAND_33[21:0];
  _RAND_34 = {1{`RANDOM}};
  tag_2_2 = _RAND_34[21:0];
  _RAND_35 = {1{`RANDOM}};
  tag_2_3 = _RAND_35[21:0];
  _RAND_36 = {1{`RANDOM}};
  tag_2_4 = _RAND_36[21:0];
  _RAND_37 = {1{`RANDOM}};
  tag_2_5 = _RAND_37[21:0];
  _RAND_38 = {1{`RANDOM}};
  tag_2_6 = _RAND_38[21:0];
  _RAND_39 = {1{`RANDOM}};
  tag_2_7 = _RAND_39[21:0];
  _RAND_40 = {1{`RANDOM}};
  tag_2_8 = _RAND_40[21:0];
  _RAND_41 = {1{`RANDOM}};
  tag_2_9 = _RAND_41[21:0];
  _RAND_42 = {1{`RANDOM}};
  tag_2_10 = _RAND_42[21:0];
  _RAND_43 = {1{`RANDOM}};
  tag_2_11 = _RAND_43[21:0];
  _RAND_44 = {1{`RANDOM}};
  tag_2_12 = _RAND_44[21:0];
  _RAND_45 = {1{`RANDOM}};
  tag_2_13 = _RAND_45[21:0];
  _RAND_46 = {1{`RANDOM}};
  tag_2_14 = _RAND_46[21:0];
  _RAND_47 = {1{`RANDOM}};
  tag_2_15 = _RAND_47[21:0];
  _RAND_48 = {1{`RANDOM}};
  tag_3_0 = _RAND_48[21:0];
  _RAND_49 = {1{`RANDOM}};
  tag_3_1 = _RAND_49[21:0];
  _RAND_50 = {1{`RANDOM}};
  tag_3_2 = _RAND_50[21:0];
  _RAND_51 = {1{`RANDOM}};
  tag_3_3 = _RAND_51[21:0];
  _RAND_52 = {1{`RANDOM}};
  tag_3_4 = _RAND_52[21:0];
  _RAND_53 = {1{`RANDOM}};
  tag_3_5 = _RAND_53[21:0];
  _RAND_54 = {1{`RANDOM}};
  tag_3_6 = _RAND_54[21:0];
  _RAND_55 = {1{`RANDOM}};
  tag_3_7 = _RAND_55[21:0];
  _RAND_56 = {1{`RANDOM}};
  tag_3_8 = _RAND_56[21:0];
  _RAND_57 = {1{`RANDOM}};
  tag_3_9 = _RAND_57[21:0];
  _RAND_58 = {1{`RANDOM}};
  tag_3_10 = _RAND_58[21:0];
  _RAND_59 = {1{`RANDOM}};
  tag_3_11 = _RAND_59[21:0];
  _RAND_60 = {1{`RANDOM}};
  tag_3_12 = _RAND_60[21:0];
  _RAND_61 = {1{`RANDOM}};
  tag_3_13 = _RAND_61[21:0];
  _RAND_62 = {1{`RANDOM}};
  tag_3_14 = _RAND_62[21:0];
  _RAND_63 = {1{`RANDOM}};
  tag_3_15 = _RAND_63[21:0];
  _RAND_64 = {1{`RANDOM}};
  valid_0_0 = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  valid_0_1 = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  valid_0_2 = _RAND_66[0:0];
  _RAND_67 = {1{`RANDOM}};
  valid_0_3 = _RAND_67[0:0];
  _RAND_68 = {1{`RANDOM}};
  valid_0_4 = _RAND_68[0:0];
  _RAND_69 = {1{`RANDOM}};
  valid_0_5 = _RAND_69[0:0];
  _RAND_70 = {1{`RANDOM}};
  valid_0_6 = _RAND_70[0:0];
  _RAND_71 = {1{`RANDOM}};
  valid_0_7 = _RAND_71[0:0];
  _RAND_72 = {1{`RANDOM}};
  valid_0_8 = _RAND_72[0:0];
  _RAND_73 = {1{`RANDOM}};
  valid_0_9 = _RAND_73[0:0];
  _RAND_74 = {1{`RANDOM}};
  valid_0_10 = _RAND_74[0:0];
  _RAND_75 = {1{`RANDOM}};
  valid_0_11 = _RAND_75[0:0];
  _RAND_76 = {1{`RANDOM}};
  valid_0_12 = _RAND_76[0:0];
  _RAND_77 = {1{`RANDOM}};
  valid_0_13 = _RAND_77[0:0];
  _RAND_78 = {1{`RANDOM}};
  valid_0_14 = _RAND_78[0:0];
  _RAND_79 = {1{`RANDOM}};
  valid_0_15 = _RAND_79[0:0];
  _RAND_80 = {1{`RANDOM}};
  valid_1_0 = _RAND_80[0:0];
  _RAND_81 = {1{`RANDOM}};
  valid_1_1 = _RAND_81[0:0];
  _RAND_82 = {1{`RANDOM}};
  valid_1_2 = _RAND_82[0:0];
  _RAND_83 = {1{`RANDOM}};
  valid_1_3 = _RAND_83[0:0];
  _RAND_84 = {1{`RANDOM}};
  valid_1_4 = _RAND_84[0:0];
  _RAND_85 = {1{`RANDOM}};
  valid_1_5 = _RAND_85[0:0];
  _RAND_86 = {1{`RANDOM}};
  valid_1_6 = _RAND_86[0:0];
  _RAND_87 = {1{`RANDOM}};
  valid_1_7 = _RAND_87[0:0];
  _RAND_88 = {1{`RANDOM}};
  valid_1_8 = _RAND_88[0:0];
  _RAND_89 = {1{`RANDOM}};
  valid_1_9 = _RAND_89[0:0];
  _RAND_90 = {1{`RANDOM}};
  valid_1_10 = _RAND_90[0:0];
  _RAND_91 = {1{`RANDOM}};
  valid_1_11 = _RAND_91[0:0];
  _RAND_92 = {1{`RANDOM}};
  valid_1_12 = _RAND_92[0:0];
  _RAND_93 = {1{`RANDOM}};
  valid_1_13 = _RAND_93[0:0];
  _RAND_94 = {1{`RANDOM}};
  valid_1_14 = _RAND_94[0:0];
  _RAND_95 = {1{`RANDOM}};
  valid_1_15 = _RAND_95[0:0];
  _RAND_96 = {1{`RANDOM}};
  valid_2_0 = _RAND_96[0:0];
  _RAND_97 = {1{`RANDOM}};
  valid_2_1 = _RAND_97[0:0];
  _RAND_98 = {1{`RANDOM}};
  valid_2_2 = _RAND_98[0:0];
  _RAND_99 = {1{`RANDOM}};
  valid_2_3 = _RAND_99[0:0];
  _RAND_100 = {1{`RANDOM}};
  valid_2_4 = _RAND_100[0:0];
  _RAND_101 = {1{`RANDOM}};
  valid_2_5 = _RAND_101[0:0];
  _RAND_102 = {1{`RANDOM}};
  valid_2_6 = _RAND_102[0:0];
  _RAND_103 = {1{`RANDOM}};
  valid_2_7 = _RAND_103[0:0];
  _RAND_104 = {1{`RANDOM}};
  valid_2_8 = _RAND_104[0:0];
  _RAND_105 = {1{`RANDOM}};
  valid_2_9 = _RAND_105[0:0];
  _RAND_106 = {1{`RANDOM}};
  valid_2_10 = _RAND_106[0:0];
  _RAND_107 = {1{`RANDOM}};
  valid_2_11 = _RAND_107[0:0];
  _RAND_108 = {1{`RANDOM}};
  valid_2_12 = _RAND_108[0:0];
  _RAND_109 = {1{`RANDOM}};
  valid_2_13 = _RAND_109[0:0];
  _RAND_110 = {1{`RANDOM}};
  valid_2_14 = _RAND_110[0:0];
  _RAND_111 = {1{`RANDOM}};
  valid_2_15 = _RAND_111[0:0];
  _RAND_112 = {1{`RANDOM}};
  valid_3_0 = _RAND_112[0:0];
  _RAND_113 = {1{`RANDOM}};
  valid_3_1 = _RAND_113[0:0];
  _RAND_114 = {1{`RANDOM}};
  valid_3_2 = _RAND_114[0:0];
  _RAND_115 = {1{`RANDOM}};
  valid_3_3 = _RAND_115[0:0];
  _RAND_116 = {1{`RANDOM}};
  valid_3_4 = _RAND_116[0:0];
  _RAND_117 = {1{`RANDOM}};
  valid_3_5 = _RAND_117[0:0];
  _RAND_118 = {1{`RANDOM}};
  valid_3_6 = _RAND_118[0:0];
  _RAND_119 = {1{`RANDOM}};
  valid_3_7 = _RAND_119[0:0];
  _RAND_120 = {1{`RANDOM}};
  valid_3_8 = _RAND_120[0:0];
  _RAND_121 = {1{`RANDOM}};
  valid_3_9 = _RAND_121[0:0];
  _RAND_122 = {1{`RANDOM}};
  valid_3_10 = _RAND_122[0:0];
  _RAND_123 = {1{`RANDOM}};
  valid_3_11 = _RAND_123[0:0];
  _RAND_124 = {1{`RANDOM}};
  valid_3_12 = _RAND_124[0:0];
  _RAND_125 = {1{`RANDOM}};
  valid_3_13 = _RAND_125[0:0];
  _RAND_126 = {1{`RANDOM}};
  valid_3_14 = _RAND_126[0:0];
  _RAND_127 = {1{`RANDOM}};
  valid_3_15 = _RAND_127[0:0];
  _RAND_128 = {1{`RANDOM}};
  dirty_0_0 = _RAND_128[0:0];
  _RAND_129 = {1{`RANDOM}};
  dirty_0_1 = _RAND_129[0:0];
  _RAND_130 = {1{`RANDOM}};
  dirty_0_2 = _RAND_130[0:0];
  _RAND_131 = {1{`RANDOM}};
  dirty_0_3 = _RAND_131[0:0];
  _RAND_132 = {1{`RANDOM}};
  dirty_0_4 = _RAND_132[0:0];
  _RAND_133 = {1{`RANDOM}};
  dirty_0_5 = _RAND_133[0:0];
  _RAND_134 = {1{`RANDOM}};
  dirty_0_6 = _RAND_134[0:0];
  _RAND_135 = {1{`RANDOM}};
  dirty_0_7 = _RAND_135[0:0];
  _RAND_136 = {1{`RANDOM}};
  dirty_0_8 = _RAND_136[0:0];
  _RAND_137 = {1{`RANDOM}};
  dirty_0_9 = _RAND_137[0:0];
  _RAND_138 = {1{`RANDOM}};
  dirty_0_10 = _RAND_138[0:0];
  _RAND_139 = {1{`RANDOM}};
  dirty_0_11 = _RAND_139[0:0];
  _RAND_140 = {1{`RANDOM}};
  dirty_0_12 = _RAND_140[0:0];
  _RAND_141 = {1{`RANDOM}};
  dirty_0_13 = _RAND_141[0:0];
  _RAND_142 = {1{`RANDOM}};
  dirty_0_14 = _RAND_142[0:0];
  _RAND_143 = {1{`RANDOM}};
  dirty_0_15 = _RAND_143[0:0];
  _RAND_144 = {1{`RANDOM}};
  dirty_1_0 = _RAND_144[0:0];
  _RAND_145 = {1{`RANDOM}};
  dirty_1_1 = _RAND_145[0:0];
  _RAND_146 = {1{`RANDOM}};
  dirty_1_2 = _RAND_146[0:0];
  _RAND_147 = {1{`RANDOM}};
  dirty_1_3 = _RAND_147[0:0];
  _RAND_148 = {1{`RANDOM}};
  dirty_1_4 = _RAND_148[0:0];
  _RAND_149 = {1{`RANDOM}};
  dirty_1_5 = _RAND_149[0:0];
  _RAND_150 = {1{`RANDOM}};
  dirty_1_6 = _RAND_150[0:0];
  _RAND_151 = {1{`RANDOM}};
  dirty_1_7 = _RAND_151[0:0];
  _RAND_152 = {1{`RANDOM}};
  dirty_1_8 = _RAND_152[0:0];
  _RAND_153 = {1{`RANDOM}};
  dirty_1_9 = _RAND_153[0:0];
  _RAND_154 = {1{`RANDOM}};
  dirty_1_10 = _RAND_154[0:0];
  _RAND_155 = {1{`RANDOM}};
  dirty_1_11 = _RAND_155[0:0];
  _RAND_156 = {1{`RANDOM}};
  dirty_1_12 = _RAND_156[0:0];
  _RAND_157 = {1{`RANDOM}};
  dirty_1_13 = _RAND_157[0:0];
  _RAND_158 = {1{`RANDOM}};
  dirty_1_14 = _RAND_158[0:0];
  _RAND_159 = {1{`RANDOM}};
  dirty_1_15 = _RAND_159[0:0];
  _RAND_160 = {1{`RANDOM}};
  dirty_2_0 = _RAND_160[0:0];
  _RAND_161 = {1{`RANDOM}};
  dirty_2_1 = _RAND_161[0:0];
  _RAND_162 = {1{`RANDOM}};
  dirty_2_2 = _RAND_162[0:0];
  _RAND_163 = {1{`RANDOM}};
  dirty_2_3 = _RAND_163[0:0];
  _RAND_164 = {1{`RANDOM}};
  dirty_2_4 = _RAND_164[0:0];
  _RAND_165 = {1{`RANDOM}};
  dirty_2_5 = _RAND_165[0:0];
  _RAND_166 = {1{`RANDOM}};
  dirty_2_6 = _RAND_166[0:0];
  _RAND_167 = {1{`RANDOM}};
  dirty_2_7 = _RAND_167[0:0];
  _RAND_168 = {1{`RANDOM}};
  dirty_2_8 = _RAND_168[0:0];
  _RAND_169 = {1{`RANDOM}};
  dirty_2_9 = _RAND_169[0:0];
  _RAND_170 = {1{`RANDOM}};
  dirty_2_10 = _RAND_170[0:0];
  _RAND_171 = {1{`RANDOM}};
  dirty_2_11 = _RAND_171[0:0];
  _RAND_172 = {1{`RANDOM}};
  dirty_2_12 = _RAND_172[0:0];
  _RAND_173 = {1{`RANDOM}};
  dirty_2_13 = _RAND_173[0:0];
  _RAND_174 = {1{`RANDOM}};
  dirty_2_14 = _RAND_174[0:0];
  _RAND_175 = {1{`RANDOM}};
  dirty_2_15 = _RAND_175[0:0];
  _RAND_176 = {1{`RANDOM}};
  dirty_3_0 = _RAND_176[0:0];
  _RAND_177 = {1{`RANDOM}};
  dirty_3_1 = _RAND_177[0:0];
  _RAND_178 = {1{`RANDOM}};
  dirty_3_2 = _RAND_178[0:0];
  _RAND_179 = {1{`RANDOM}};
  dirty_3_3 = _RAND_179[0:0];
  _RAND_180 = {1{`RANDOM}};
  dirty_3_4 = _RAND_180[0:0];
  _RAND_181 = {1{`RANDOM}};
  dirty_3_5 = _RAND_181[0:0];
  _RAND_182 = {1{`RANDOM}};
  dirty_3_6 = _RAND_182[0:0];
  _RAND_183 = {1{`RANDOM}};
  dirty_3_7 = _RAND_183[0:0];
  _RAND_184 = {1{`RANDOM}};
  dirty_3_8 = _RAND_184[0:0];
  _RAND_185 = {1{`RANDOM}};
  dirty_3_9 = _RAND_185[0:0];
  _RAND_186 = {1{`RANDOM}};
  dirty_3_10 = _RAND_186[0:0];
  _RAND_187 = {1{`RANDOM}};
  dirty_3_11 = _RAND_187[0:0];
  _RAND_188 = {1{`RANDOM}};
  dirty_3_12 = _RAND_188[0:0];
  _RAND_189 = {1{`RANDOM}};
  dirty_3_13 = _RAND_189[0:0];
  _RAND_190 = {1{`RANDOM}};
  dirty_3_14 = _RAND_190[0:0];
  _RAND_191 = {1{`RANDOM}};
  dirty_3_15 = _RAND_191[0:0];
  _RAND_192 = {1{`RANDOM}};
  wait_r = _RAND_192[0:0];
  _RAND_193 = {1{`RANDOM}};
  valid_r = _RAND_193[0:0];
  _RAND_194 = {1{`RANDOM}};
  flush_r = _RAND_194[0:0];
  _RAND_195 = {1{`RANDOM}};
  mode_r = _RAND_195[4:0];
  _RAND_196 = {2{`RANDOM}};
  wdata_r = _RAND_196[63:0];
  _RAND_197 = {1{`RANDOM}};
  amo_r = _RAND_197[4:0];
  _RAND_198 = {1{`RANDOM}};
  addr_r = _RAND_198[31:0];
  _RAND_199 = {1{`RANDOM}};
  matchWay_r = _RAND_199[1:0];
  _RAND_200 = {1{`RANDOM}};
  offset = _RAND_200[2:0];
  _RAND_201 = {2{`RANDOM}};
  rdatabuf = _RAND_201[63:0];
  _RAND_202 = {1{`RANDOM}};
  blockIdx_r = _RAND_202[3:0];
  _RAND_203 = {1{`RANDOM}};
  state = _RAND_203[2:0];
  _RAND_204 = {1{`RANDOM}};
  axiRdataEn = _RAND_204[0:0];
  _RAND_205 = {1{`RANDOM}};
  axiRaddrEn = _RAND_205[0:0];
  _RAND_206 = {1{`RANDOM}};
  axiWaddrEn = _RAND_206[0:0];
  _RAND_207 = {1{`RANDOM}};
  axiWdataEn = _RAND_207[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ToAXI(
  input         clock,
  input         reset,
  input  [31:0] io_dataIO_addr, // @[playground/src/axi/toaxi.scala 61:16]
  output [63:0] io_dataIO_rdata, // @[playground/src/axi/toaxi.scala 61:16]
  output        io_dataIO_rvalid, // @[playground/src/axi/toaxi.scala 61:16]
  input  [63:0] io_dataIO_wdata, // @[playground/src/axi/toaxi.scala 61:16]
  input  [4:0]  io_dataIO_dc_mode, // @[playground/src/axi/toaxi.scala 61:16]
  output        io_dataIO_ready, // @[playground/src/axi/toaxi.scala 61:16]
  input         io_outAxi_wa_ready, // @[playground/src/axi/toaxi.scala 61:16]
  output        io_outAxi_wa_valid, // @[playground/src/axi/toaxi.scala 61:16]
  output [3:0]  io_outAxi_wa_bits_id, // @[playground/src/axi/toaxi.scala 61:16]
  output [31:0] io_outAxi_wa_bits_addr, // @[playground/src/axi/toaxi.scala 61:16]
  output [7:0]  io_outAxi_wa_bits_len, // @[playground/src/axi/toaxi.scala 61:16]
  output [2:0]  io_outAxi_wa_bits_size, // @[playground/src/axi/toaxi.scala 61:16]
  output [1:0]  io_outAxi_wa_bits_burst, // @[playground/src/axi/toaxi.scala 61:16]
  input         io_outAxi_wd_ready, // @[playground/src/axi/toaxi.scala 61:16]
  output        io_outAxi_wd_valid, // @[playground/src/axi/toaxi.scala 61:16]
  output [63:0] io_outAxi_wd_bits_data, // @[playground/src/axi/toaxi.scala 61:16]
  output [7:0]  io_outAxi_wd_bits_strb, // @[playground/src/axi/toaxi.scala 61:16]
  output        io_outAxi_wd_bits_last, // @[playground/src/axi/toaxi.scala 61:16]
  output        io_outAxi_wr_ready, // @[playground/src/axi/toaxi.scala 61:16]
  input         io_outAxi_wr_valid, // @[playground/src/axi/toaxi.scala 61:16]
  input  [3:0]  io_outAxi_wr_bits_id, // @[playground/src/axi/toaxi.scala 61:16]
  input  [1:0]  io_outAxi_wr_bits_resp, // @[playground/src/axi/toaxi.scala 61:16]
  input         io_outAxi_ra_ready, // @[playground/src/axi/toaxi.scala 61:16]
  output        io_outAxi_ra_valid, // @[playground/src/axi/toaxi.scala 61:16]
  output [3:0]  io_outAxi_ra_bits_id, // @[playground/src/axi/toaxi.scala 61:16]
  output [31:0] io_outAxi_ra_bits_addr, // @[playground/src/axi/toaxi.scala 61:16]
  output [7:0]  io_outAxi_ra_bits_len, // @[playground/src/axi/toaxi.scala 61:16]
  output [2:0]  io_outAxi_ra_bits_size, // @[playground/src/axi/toaxi.scala 61:16]
  output [1:0]  io_outAxi_ra_bits_burst, // @[playground/src/axi/toaxi.scala 61:16]
  output        io_outAxi_rd_ready, // @[playground/src/axi/toaxi.scala 61:16]
  input         io_outAxi_rd_valid, // @[playground/src/axi/toaxi.scala 61:16]
  input  [3:0]  io_outAxi_rd_bits_id, // @[playground/src/axi/toaxi.scala 61:16]
  input  [63:0] io_outAxi_rd_bits_data, // @[playground/src/axi/toaxi.scala 61:16]
  input  [1:0]  io_outAxi_rd_bits_resp, // @[playground/src/axi/toaxi.scala 61:16]
  input         io_outAxi_rd_bits_last // @[playground/src/axi/toaxi.scala 61:16]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [63:0] _RAND_14;
  reg [31:0] _RAND_15;
`endif // RANDOMIZE_REG_INIT
  reg  waddrEn; // @[playground/src/axi/toaxi.scala 66:26]
  reg [31:0] waddr; // @[playground/src/axi/toaxi.scala 67:26]
  reg [2:0] wsize; // @[playground/src/axi/toaxi.scala 68:26]
  reg  wdataEn; // @[playground/src/axi/toaxi.scala 71:26]
  reg [63:0] wdata; // @[playground/src/axi/toaxi.scala 72:26]
  reg [7:0] wstrb; // @[playground/src/axi/toaxi.scala 73:26]
  reg [2:0] rsize; // @[playground/src/axi/toaxi.scala 75:26]
  reg  raddrEn; // @[playground/src/axi/toaxi.scala 76:26]
  reg [31:0] raddr; // @[playground/src/axi/toaxi.scala 77:26]
  reg  rdataEn; // @[playground/src/axi/toaxi.scala 78:26]
  reg [63:0] rdata; // @[playground/src/axi/toaxi.scala 79:26]
  reg [31:0] pre_addr; // @[playground/src/axi/toaxi.scala 81:27]
  reg [4:0] mode; // @[playground/src/axi/toaxi.scala 85:23]
  reg [2:0] state; // @[playground/src/axi/toaxi.scala 92:25]
  wire  _wtype_T_1 = 5'h8 == io_dataIO_dc_mode; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _wtype_T_3 = 5'h9 == io_dataIO_dc_mode; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _wtype_T_5 = 5'ha == io_dataIO_dc_mode; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _wtype_T_7 = 5'hb == io_dataIO_dc_mode; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire [2:0] _wtype_T_8 = _wtype_T_7 ? 3'h3 : 3'h0; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _wtype_T_9 = _wtype_T_5 ? 3'h2 : _wtype_T_8; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _wtype_T_10 = _wtype_T_3 ? 3'h1 : _wtype_T_9; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [7:0] _wtype_T_11 = _wtype_T_7 ? 8'hff : 8'h0; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [7:0] _wtype_T_12 = _wtype_T_5 ? 8'hf : _wtype_T_11; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [7:0] _wtype_T_13 = _wtype_T_3 ? 8'h3 : _wtype_T_12; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [7:0] wtype_1 = _wtype_T_1 ? 8'h1 : _wtype_T_13; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [14:0] _GEN_69 = {{7'd0}, wtype_1}; // @[playground/src/axi/toaxi.scala 113:37]
  wire [14:0] _wstrb_T_1 = _GEN_69 << io_dataIO_addr[2:0]; // @[playground/src/axi/toaxi.scala 113:37]
  wire [6:0] _wdata_T_1 = io_dataIO_addr[2:0] * 4'h8; // @[playground/src/axi/toaxi.scala 114:55]
  wire [190:0] _GEN_84 = {{127'd0}, io_dataIO_wdata}; // @[playground/src/axi/toaxi.scala 114:38]
  wire [190:0] _wdata_T_2 = _GEN_84 << _wdata_T_1; // @[playground/src/axi/toaxi.scala 114:38]
  wire [2:0] _rsize_T_5 = 5'h5 == io_dataIO_dc_mode ? 3'h1 : 3'h0; // @[src/main/scala/chisel3/util/Mux.scala 81:58]
  wire [2:0] _rsize_T_7 = 5'h15 == io_dataIO_dc_mode ? 3'h1 : _rsize_T_5; // @[src/main/scala/chisel3/util/Mux.scala 81:58]
  wire [2:0] _rsize_T_9 = 5'h6 == io_dataIO_dc_mode ? 3'h2 : _rsize_T_7; // @[src/main/scala/chisel3/util/Mux.scala 81:58]
  wire [2:0] _rsize_T_11 = 5'h16 == io_dataIO_dc_mode ? 3'h2 : _rsize_T_9; // @[src/main/scala/chisel3/util/Mux.scala 81:58]
  wire [2:0] _rsize_T_13 = 5'h7 == io_dataIO_dc_mode ? 3'h3 : _rsize_T_11; // @[src/main/scala/chisel3/util/Mux.scala 81:58]
  wire  _GEN_4 = io_dataIO_dc_mode[2] | raddrEn; // @[playground/src/axi/toaxi.scala 116:43 130:25 76:26]
  wire  _GEN_8 = io_dataIO_dc_mode[3] | waddrEn; // @[playground/src/axi/toaxi.scala 101:37 105:25 66:26]
  wire [14:0] _GEN_10 = io_dataIO_dc_mode[3] ? _wstrb_T_1 : {{7'd0}, wstrb}; // @[playground/src/axi/toaxi.scala 101:37 113:25 73:26]
  wire [2:0] _GEN_21 = io_outAxi_wd_ready ? 3'h3 : state; // @[playground/src/axi/toaxi.scala 144:37 92:25]
  wire  _GEN_22 = raddrEn & io_outAxi_ra_ready ? 1'h0 : raddrEn; // @[playground/src/axi/toaxi.scala 157:48 158:25 76:26]
  wire [2:0] _GEN_24 = raddrEn & io_outAxi_ra_ready ? 3'h5 : state; // @[playground/src/axi/toaxi.scala 157:48 160:25 92:25]
  wire [2:0] strb_offset = pre_addr[2:0]; // @[playground/src/axi/toaxi.scala 169:43]
  wire [6:0] _tem_rdata_T = 4'h8 * strb_offset; // @[playground/src/axi/toaxi.scala 172:72]
  wire [63:0] _tem_rdata_T_1 = io_outAxi_rd_bits_data >> _tem_rdata_T; // @[playground/src/axi/toaxi.scala 172:64]
  wire [7:0] _tem_rdata_T_3 = _tem_rdata_T_1[7:0]; // @[playground/src/axi/toaxi.scala 172:94]
  wire [15:0] _tem_rdata_T_7 = _tem_rdata_T_1[15:0]; // @[playground/src/axi/toaxi.scala 176:95]
  wire [31:0] _tem_rdata_T_11 = _tem_rdata_T_1[31:0]; // @[playground/src/axi/toaxi.scala 180:95]
  wire [31:0] _GEN_29 = 5'h6 == mode ? $signed(_tem_rdata_T_11) : $signed(32'sh0); // @[playground/src/axi/toaxi.scala 168:29 170:29 180:37]
  wire [31:0] _GEN_31 = 5'h5 == mode ? $signed({{16{_tem_rdata_T_7[15]}},_tem_rdata_T_7}) : $signed(_GEN_29); // @[playground/src/axi/toaxi.scala 170:29 176:37]
  wire [31:0] _GEN_33 = 5'h4 == mode ? $signed({{24{_tem_rdata_T_3[7]}},_tem_rdata_T_3}) : $signed(_GEN_31); // @[playground/src/axi/toaxi.scala 170:29 172:37]
  wire [63:0] _rdata_T = {{32{_GEN_33[31]}},_GEN_33}; // @[playground/src/axi/toaxi.scala 173:50]
  wire [63:0] _GEN_25 = 5'h16 == mode ? {{32'd0}, _tem_rdata_T_1[31:0]} : rdata; // @[playground/src/axi/toaxi.scala 170:29 193:33 79:26]
  wire [63:0] _GEN_26 = 5'h15 == mode ? {{48'd0}, _tem_rdata_T_1[15:0]} : _GEN_25; // @[playground/src/axi/toaxi.scala 170:29 190:33]
  wire [63:0] _GEN_27 = 5'h14 == mode ? {{56'd0}, _tem_rdata_T_1[7:0]} : _GEN_26; // @[playground/src/axi/toaxi.scala 170:29 187:33]
  wire [63:0] _GEN_28 = 5'h7 == mode ? io_outAxi_rd_bits_data : _GEN_27; // @[playground/src/axi/toaxi.scala 170:29 184:37]
  wire [63:0] _GEN_30 = 5'h6 == mode ? _rdata_T : _GEN_28; // @[playground/src/axi/toaxi.scala 170:29 181:37]
  wire [63:0] _GEN_32 = 5'h5 == mode ? _rdata_T : _GEN_30; // @[playground/src/axi/toaxi.scala 170:29 177:37]
  wire [63:0] _GEN_34 = 5'h4 == mode ? _rdata_T : _GEN_32; // @[playground/src/axi/toaxi.scala 170:29 173:37]
  wire [63:0] _GEN_35 = rdataEn & io_outAxi_rd_valid ? _GEN_34 : rdata; // @[playground/src/axi/toaxi.scala 166:48 79:26]
  wire  _GEN_37 = rdataEn & io_outAxi_rd_valid ? 1'h0 : 1'h1; // @[playground/src/axi/toaxi.scala 164:21 166:48 198:25]
  wire [2:0] _GEN_38 = rdataEn & io_outAxi_rd_valid ? 3'h6 : state; // @[playground/src/axi/toaxi.scala 166:48 199:25 92:25]
  wire [2:0] _GEN_39 = 3'h6 == state ? 3'h0 : state; // @[playground/src/axi/toaxi.scala 95:18 203:19 92:25]
  wire  _GEN_40 = 3'h5 == state ? _GEN_37 : rdataEn; // @[playground/src/axi/toaxi.scala 95:18 78:26]
  wire [63:0] _GEN_41 = 3'h5 == state ? _GEN_35 : rdata; // @[playground/src/axi/toaxi.scala 95:18 79:26]
  wire [2:0] _GEN_43 = 3'h5 == state ? _GEN_38 : _GEN_39; // @[playground/src/axi/toaxi.scala 95:18]
  wire  _GEN_44 = 3'h4 == state ? _GEN_22 : raddrEn; // @[playground/src/axi/toaxi.scala 95:18 76:26]
  wire [2:0] _GEN_46 = 3'h4 == state ? _GEN_24 : _GEN_43; // @[playground/src/axi/toaxi.scala 95:18]
  wire  _GEN_47 = 3'h4 == state ? rdataEn : _GEN_40; // @[playground/src/axi/toaxi.scala 95:18 78:26]
  wire [63:0] _GEN_48 = 3'h4 == state ? rdata : _GEN_41; // @[playground/src/axi/toaxi.scala 95:18 79:26]
  wire  _GEN_49 = 3'h3 == state ? 1'h0 : wdataEn; // @[playground/src/axi/toaxi.scala 95:18 152:21 71:26]
  wire [2:0] _GEN_50 = 3'h3 == state ? 3'h0 : _GEN_46; // @[playground/src/axi/toaxi.scala 95:18 153:21]
  wire  _GEN_51 = 3'h3 == state ? raddrEn : _GEN_44; // @[playground/src/axi/toaxi.scala 95:18 76:26]
  wire  _GEN_53 = 3'h3 == state ? rdataEn : _GEN_47; // @[playground/src/axi/toaxi.scala 95:18 78:26]
  wire [63:0] _GEN_54 = 3'h3 == state ? rdata : _GEN_48; // @[playground/src/axi/toaxi.scala 95:18 79:26]
  wire  _GEN_55 = 3'h2 == state | _GEN_49; // @[playground/src/axi/toaxi.scala 95:18 143:21]
  wire [14:0] _GEN_74 = 3'h0 == state ? _GEN_10 : {{7'd0}, wstrb}; // @[playground/src/axi/toaxi.scala 95:18 73:26]
  reg [63:0] out_rdata; // @[playground/src/axi/toaxi.scala 208:28]
  reg  out_valid; // @[playground/src/axi/toaxi.scala 209:28]
  wire [14:0] _GEN_0 = reset ? 15'h0 : _GEN_74; // @[playground/src/axi/toaxi.scala 73:{26,26}]
  assign io_dataIO_rdata = out_rdata; // @[playground/src/axi/toaxi.scala 213:25]
  assign io_dataIO_rvalid = out_valid; // @[playground/src/axi/toaxi.scala 212:25]
  assign io_dataIO_ready = state == 3'h0; // @[playground/src/axi/toaxi.scala 206:31]
  assign io_outAxi_wa_valid = waddrEn; // @[playground/src/axi/toaxi.scala 217:31]
  assign io_outAxi_wa_bits_id = 4'h0; // @[playground/src/axi/axi.scala 41:{38,38}]
  assign io_outAxi_wa_bits_addr = waddr; // @[playground/src/axi/toaxi.scala 218:31]
  assign io_outAxi_wa_bits_len = 8'h0; // @[playground/src/axi/toaxi.scala 219:31]
  assign io_outAxi_wa_bits_size = wsize; // @[playground/src/axi/toaxi.scala 220:31]
  assign io_outAxi_wa_bits_burst = 2'h1; // @[playground/src/axi/toaxi.scala 221:31]
  assign io_outAxi_wd_valid = wdataEn; // @[playground/src/axi/toaxi.scala 223:31]
  assign io_outAxi_wd_bits_data = wdata; // @[playground/src/axi/toaxi.scala 224:31]
  assign io_outAxi_wd_bits_strb = wstrb; // @[playground/src/axi/toaxi.scala 225:31]
  assign io_outAxi_wd_bits_last = 1'h1; // @[playground/src/axi/toaxi.scala 70:27]
  assign io_outAxi_wr_ready = 1'h1; // @[playground/src/axi/toaxi.scala 228:31]
  assign io_outAxi_ra_valid = raddrEn; // @[playground/src/axi/toaxi.scala 230:31]
  assign io_outAxi_ra_bits_id = 4'h0; // @[playground/src/axi/axi.scala 41:{38,38}]
  assign io_outAxi_ra_bits_addr = raddr; // @[playground/src/axi/toaxi.scala 231:31]
  assign io_outAxi_ra_bits_len = 8'h0; // @[playground/src/axi/toaxi.scala 232:31]
  assign io_outAxi_ra_bits_size = rsize; // @[playground/src/axi/toaxi.scala 233:31]
  assign io_outAxi_ra_bits_burst = 2'h1; // @[playground/src/axi/toaxi.scala 234:31]
  assign io_outAxi_rd_ready = rdataEn; // @[playground/src/axi/toaxi.scala 236:31]
  always @(posedge clock) begin
    if (reset) begin // @[playground/src/axi/toaxi.scala 66:26]
      waddrEn <= 1'h0; // @[playground/src/axi/toaxi.scala 66:26]
    end else if (3'h0 == state) begin // @[playground/src/axi/toaxi.scala 95:18]
      waddrEn <= _GEN_8;
    end else if (3'h1 == state) begin // @[playground/src/axi/toaxi.scala 95:18]
      if (waddrEn & io_outAxi_wa_ready) begin // @[playground/src/axi/toaxi.scala 136:48]
        waddrEn <= 1'h0; // @[playground/src/axi/toaxi.scala 137:25]
      end
    end
    if (reset) begin // @[playground/src/axi/toaxi.scala 67:26]
      waddr <= 32'h0; // @[playground/src/axi/toaxi.scala 67:26]
    end else if (3'h0 == state) begin // @[playground/src/axi/toaxi.scala 95:18]
      if (io_dataIO_dc_mode[3]) begin // @[playground/src/axi/toaxi.scala 101:37]
        waddr <= io_dataIO_addr; // @[playground/src/axi/toaxi.scala 103:25]
      end
    end
    if (reset) begin // @[playground/src/axi/toaxi.scala 68:26]
      wsize <= 3'h0; // @[playground/src/axi/toaxi.scala 68:26]
    end else if (3'h0 == state) begin // @[playground/src/axi/toaxi.scala 95:18]
      if (io_dataIO_dc_mode[3]) begin // @[playground/src/axi/toaxi.scala 101:37]
        if (_wtype_T_1) begin // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
          wsize <= 3'h0;
        end else begin
          wsize <= _wtype_T_10;
        end
      end
    end
    if (reset) begin // @[playground/src/axi/toaxi.scala 71:26]
      wdataEn <= 1'h0; // @[playground/src/axi/toaxi.scala 71:26]
    end else if (!(3'h0 == state)) begin // @[playground/src/axi/toaxi.scala 95:18]
      if (!(3'h1 == state)) begin // @[playground/src/axi/toaxi.scala 95:18]
        wdataEn <= _GEN_55;
      end
    end
    if (reset) begin // @[playground/src/axi/toaxi.scala 72:26]
      wdata <= 64'h0; // @[playground/src/axi/toaxi.scala 72:26]
    end else if (3'h0 == state) begin // @[playground/src/axi/toaxi.scala 95:18]
      if (io_dataIO_dc_mode[3]) begin // @[playground/src/axi/toaxi.scala 101:37]
        wdata <= _wdata_T_2[63:0]; // @[playground/src/axi/toaxi.scala 114:25]
      end
    end
    wstrb <= _GEN_0[7:0]; // @[playground/src/axi/toaxi.scala 73:{26,26}]
    if (reset) begin // @[playground/src/axi/toaxi.scala 75:26]
      rsize <= 3'h0; // @[playground/src/axi/toaxi.scala 75:26]
    end else if (3'h0 == state) begin // @[playground/src/axi/toaxi.scala 95:18]
      if (!(io_dataIO_dc_mode[3])) begin // @[playground/src/axi/toaxi.scala 101:37]
        if (io_dataIO_dc_mode[2]) begin // @[playground/src/axi/toaxi.scala 116:43]
          rsize <= _rsize_T_13; // @[playground/src/axi/toaxi.scala 118:23]
        end
      end
    end
    if (reset) begin // @[playground/src/axi/toaxi.scala 76:26]
      raddrEn <= 1'h0; // @[playground/src/axi/toaxi.scala 76:26]
    end else if (3'h0 == state) begin // @[playground/src/axi/toaxi.scala 95:18]
      if (!(io_dataIO_dc_mode[3])) begin // @[playground/src/axi/toaxi.scala 101:37]
        raddrEn <= _GEN_4;
      end
    end else if (!(3'h1 == state)) begin // @[playground/src/axi/toaxi.scala 95:18]
      if (!(3'h2 == state)) begin // @[playground/src/axi/toaxi.scala 95:18]
        raddrEn <= _GEN_51;
      end
    end
    if (reset) begin // @[playground/src/axi/toaxi.scala 77:26]
      raddr <= 32'h0; // @[playground/src/axi/toaxi.scala 77:26]
    end else if (3'h0 == state) begin // @[playground/src/axi/toaxi.scala 95:18]
      if (!(io_dataIO_dc_mode[3])) begin // @[playground/src/axi/toaxi.scala 101:37]
        if (io_dataIO_dc_mode[2]) begin // @[playground/src/axi/toaxi.scala 116:43]
          raddr <= io_dataIO_addr; // @[playground/src/axi/toaxi.scala 129:23]
        end
      end
    end
    if (reset) begin // @[playground/src/axi/toaxi.scala 78:26]
      rdataEn <= 1'h0; // @[playground/src/axi/toaxi.scala 78:26]
    end else if (!(3'h0 == state)) begin // @[playground/src/axi/toaxi.scala 95:18]
      if (!(3'h1 == state)) begin // @[playground/src/axi/toaxi.scala 95:18]
        if (!(3'h2 == state)) begin // @[playground/src/axi/toaxi.scala 95:18]
          rdataEn <= _GEN_53;
        end
      end
    end
    if (reset) begin // @[playground/src/axi/toaxi.scala 79:26]
      rdata <= 64'h0; // @[playground/src/axi/toaxi.scala 79:26]
    end else if (!(3'h0 == state)) begin // @[playground/src/axi/toaxi.scala 95:18]
      if (!(3'h1 == state)) begin // @[playground/src/axi/toaxi.scala 95:18]
        if (!(3'h2 == state)) begin // @[playground/src/axi/toaxi.scala 95:18]
          rdata <= _GEN_54;
        end
      end
    end
    if (reset) begin // @[playground/src/axi/toaxi.scala 81:27]
      pre_addr <= 32'h0; // @[playground/src/axi/toaxi.scala 81:27]
    end else if (3'h0 == state) begin // @[playground/src/axi/toaxi.scala 95:18]
      if (io_dataIO_dc_mode[3]) begin // @[playground/src/axi/toaxi.scala 101:37]
        pre_addr <= io_dataIO_addr; // @[playground/src/axi/toaxi.scala 115:26]
      end else if (io_dataIO_dc_mode[2]) begin // @[playground/src/axi/toaxi.scala 116:43]
        pre_addr <= io_dataIO_addr; // @[playground/src/axi/toaxi.scala 131:26]
      end
    end
    if (reset) begin // @[playground/src/axi/toaxi.scala 85:23]
      mode <= 5'h0; // @[playground/src/axi/toaxi.scala 85:23]
    end else if (3'h0 == state) begin // @[playground/src/axi/toaxi.scala 95:18]
      mode <= io_dataIO_dc_mode; // @[playground/src/axi/toaxi.scala 97:21]
    end
    if (reset) begin // @[playground/src/axi/toaxi.scala 92:25]
      state <= 3'h0; // @[playground/src/axi/toaxi.scala 92:25]
    end else if (3'h0 == state) begin // @[playground/src/axi/toaxi.scala 95:18]
      if (io_dataIO_dc_mode[3]) begin // @[playground/src/axi/toaxi.scala 101:37]
        state <= 3'h1; // @[playground/src/axi/toaxi.scala 102:25]
      end else if (io_dataIO_dc_mode[2]) begin // @[playground/src/axi/toaxi.scala 116:43]
        state <= 3'h4; // @[playground/src/axi/toaxi.scala 117:23]
      end
    end else if (3'h1 == state) begin // @[playground/src/axi/toaxi.scala 95:18]
      if (waddrEn & io_outAxi_wa_ready) begin // @[playground/src/axi/toaxi.scala 136:48]
        state <= 3'h2; // @[playground/src/axi/toaxi.scala 139:25]
      end
    end else if (3'h2 == state) begin // @[playground/src/axi/toaxi.scala 95:18]
      state <= _GEN_21;
    end else begin
      state <= _GEN_50;
    end
    if (reset) begin // @[playground/src/axi/toaxi.scala 208:28]
      out_rdata <= 64'h0; // @[playground/src/axi/toaxi.scala 208:28]
    end else begin
      out_rdata <= rdata; // @[playground/src/axi/toaxi.scala 211:15]
    end
    if (reset) begin // @[playground/src/axi/toaxi.scala 209:28]
      out_valid <= 1'h0; // @[playground/src/axi/toaxi.scala 209:28]
    end else begin
      out_valid <= state == 3'h6 | state == 3'h3; // @[playground/src/axi/toaxi.scala 210:15]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  waddrEn = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  waddr = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  wsize = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  wdataEn = _RAND_3[0:0];
  _RAND_4 = {2{`RANDOM}};
  wdata = _RAND_4[63:0];
  _RAND_5 = {1{`RANDOM}};
  wstrb = _RAND_5[7:0];
  _RAND_6 = {1{`RANDOM}};
  rsize = _RAND_6[2:0];
  _RAND_7 = {1{`RANDOM}};
  raddrEn = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  raddr = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  rdataEn = _RAND_9[0:0];
  _RAND_10 = {2{`RANDOM}};
  rdata = _RAND_10[63:0];
  _RAND_11 = {1{`RANDOM}};
  pre_addr = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  mode = _RAND_12[4:0];
  _RAND_13 = {1{`RANDOM}};
  state = _RAND_13[2:0];
  _RAND_14 = {2{`RANDOM}};
  out_rdata = _RAND_14[63:0];
  _RAND_15 = {1{`RANDOM}};
  out_valid = _RAND_15[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module CrossBar(
  input         clock,
  input         reset,
  output        io_icAxi_ra_ready, // @[playground/src/noop/crossbar.scala 18:16]
  input         io_icAxi_ra_valid, // @[playground/src/noop/crossbar.scala 18:16]
  input  [31:0] io_icAxi_ra_bits_addr, // @[playground/src/noop/crossbar.scala 18:16]
  output        io_icAxi_rd_valid, // @[playground/src/noop/crossbar.scala 18:16]
  output [63:0] io_icAxi_rd_bits_data, // @[playground/src/noop/crossbar.scala 18:16]
  output        io_icAxi_rd_bits_last, // @[playground/src/noop/crossbar.scala 18:16]
  output        io_flashAxi_wa_ready, // @[playground/src/noop/crossbar.scala 18:16]
  input         io_flashAxi_wa_valid, // @[playground/src/noop/crossbar.scala 18:16]
  input  [3:0]  io_flashAxi_wa_bits_id, // @[playground/src/noop/crossbar.scala 18:16]
  input  [31:0] io_flashAxi_wa_bits_addr, // @[playground/src/noop/crossbar.scala 18:16]
  input  [7:0]  io_flashAxi_wa_bits_len, // @[playground/src/noop/crossbar.scala 18:16]
  input  [2:0]  io_flashAxi_wa_bits_size, // @[playground/src/noop/crossbar.scala 18:16]
  input  [1:0]  io_flashAxi_wa_bits_burst, // @[playground/src/noop/crossbar.scala 18:16]
  output        io_flashAxi_wd_ready, // @[playground/src/noop/crossbar.scala 18:16]
  input         io_flashAxi_wd_valid, // @[playground/src/noop/crossbar.scala 18:16]
  input  [63:0] io_flashAxi_wd_bits_data, // @[playground/src/noop/crossbar.scala 18:16]
  input  [7:0]  io_flashAxi_wd_bits_strb, // @[playground/src/noop/crossbar.scala 18:16]
  input         io_flashAxi_wd_bits_last, // @[playground/src/noop/crossbar.scala 18:16]
  input         io_flashAxi_wr_ready, // @[playground/src/noop/crossbar.scala 18:16]
  output        io_flashAxi_wr_valid, // @[playground/src/noop/crossbar.scala 18:16]
  output [3:0]  io_flashAxi_wr_bits_id, // @[playground/src/noop/crossbar.scala 18:16]
  output [1:0]  io_flashAxi_wr_bits_resp, // @[playground/src/noop/crossbar.scala 18:16]
  output        io_flashAxi_ra_ready, // @[playground/src/noop/crossbar.scala 18:16]
  input         io_flashAxi_ra_valid, // @[playground/src/noop/crossbar.scala 18:16]
  input  [3:0]  io_flashAxi_ra_bits_id, // @[playground/src/noop/crossbar.scala 18:16]
  input  [31:0] io_flashAxi_ra_bits_addr, // @[playground/src/noop/crossbar.scala 18:16]
  input  [7:0]  io_flashAxi_ra_bits_len, // @[playground/src/noop/crossbar.scala 18:16]
  input  [2:0]  io_flashAxi_ra_bits_size, // @[playground/src/noop/crossbar.scala 18:16]
  input  [1:0]  io_flashAxi_ra_bits_burst, // @[playground/src/noop/crossbar.scala 18:16]
  input         io_flashAxi_rd_ready, // @[playground/src/noop/crossbar.scala 18:16]
  output        io_flashAxi_rd_valid, // @[playground/src/noop/crossbar.scala 18:16]
  output [3:0]  io_flashAxi_rd_bits_id, // @[playground/src/noop/crossbar.scala 18:16]
  output [63:0] io_flashAxi_rd_bits_data, // @[playground/src/noop/crossbar.scala 18:16]
  output [1:0]  io_flashAxi_rd_bits_resp, // @[playground/src/noop/crossbar.scala 18:16]
  output        io_flashAxi_rd_bits_last, // @[playground/src/noop/crossbar.scala 18:16]
  output        io_memAxi_wa_ready, // @[playground/src/noop/crossbar.scala 18:16]
  input         io_memAxi_wa_valid, // @[playground/src/noop/crossbar.scala 18:16]
  input  [31:0] io_memAxi_wa_bits_addr, // @[playground/src/noop/crossbar.scala 18:16]
  output        io_memAxi_wd_ready, // @[playground/src/noop/crossbar.scala 18:16]
  input         io_memAxi_wd_valid, // @[playground/src/noop/crossbar.scala 18:16]
  input  [63:0] io_memAxi_wd_bits_data, // @[playground/src/noop/crossbar.scala 18:16]
  input         io_memAxi_wd_bits_last, // @[playground/src/noop/crossbar.scala 18:16]
  output        io_memAxi_ra_ready, // @[playground/src/noop/crossbar.scala 18:16]
  input         io_memAxi_ra_valid, // @[playground/src/noop/crossbar.scala 18:16]
  input  [31:0] io_memAxi_ra_bits_addr, // @[playground/src/noop/crossbar.scala 18:16]
  output        io_memAxi_rd_valid, // @[playground/src/noop/crossbar.scala 18:16]
  output [63:0] io_memAxi_rd_bits_data, // @[playground/src/noop/crossbar.scala 18:16]
  output        io_memAxi_rd_bits_last, // @[playground/src/noop/crossbar.scala 18:16]
  output        io_mmioAxi_wa_ready, // @[playground/src/noop/crossbar.scala 18:16]
  input         io_mmioAxi_wa_valid, // @[playground/src/noop/crossbar.scala 18:16]
  input  [3:0]  io_mmioAxi_wa_bits_id, // @[playground/src/noop/crossbar.scala 18:16]
  input  [31:0] io_mmioAxi_wa_bits_addr, // @[playground/src/noop/crossbar.scala 18:16]
  input  [7:0]  io_mmioAxi_wa_bits_len, // @[playground/src/noop/crossbar.scala 18:16]
  input  [2:0]  io_mmioAxi_wa_bits_size, // @[playground/src/noop/crossbar.scala 18:16]
  input  [1:0]  io_mmioAxi_wa_bits_burst, // @[playground/src/noop/crossbar.scala 18:16]
  output        io_mmioAxi_wd_ready, // @[playground/src/noop/crossbar.scala 18:16]
  input         io_mmioAxi_wd_valid, // @[playground/src/noop/crossbar.scala 18:16]
  input  [63:0] io_mmioAxi_wd_bits_data, // @[playground/src/noop/crossbar.scala 18:16]
  input  [7:0]  io_mmioAxi_wd_bits_strb, // @[playground/src/noop/crossbar.scala 18:16]
  input         io_mmioAxi_wd_bits_last, // @[playground/src/noop/crossbar.scala 18:16]
  input         io_mmioAxi_wr_ready, // @[playground/src/noop/crossbar.scala 18:16]
  output        io_mmioAxi_wr_valid, // @[playground/src/noop/crossbar.scala 18:16]
  output [3:0]  io_mmioAxi_wr_bits_id, // @[playground/src/noop/crossbar.scala 18:16]
  output [1:0]  io_mmioAxi_wr_bits_resp, // @[playground/src/noop/crossbar.scala 18:16]
  output        io_mmioAxi_ra_ready, // @[playground/src/noop/crossbar.scala 18:16]
  input         io_mmioAxi_ra_valid, // @[playground/src/noop/crossbar.scala 18:16]
  input  [3:0]  io_mmioAxi_ra_bits_id, // @[playground/src/noop/crossbar.scala 18:16]
  input  [31:0] io_mmioAxi_ra_bits_addr, // @[playground/src/noop/crossbar.scala 18:16]
  input  [7:0]  io_mmioAxi_ra_bits_len, // @[playground/src/noop/crossbar.scala 18:16]
  input  [2:0]  io_mmioAxi_ra_bits_size, // @[playground/src/noop/crossbar.scala 18:16]
  input  [1:0]  io_mmioAxi_ra_bits_burst, // @[playground/src/noop/crossbar.scala 18:16]
  input         io_mmioAxi_rd_ready, // @[playground/src/noop/crossbar.scala 18:16]
  output        io_mmioAxi_rd_valid, // @[playground/src/noop/crossbar.scala 18:16]
  output [3:0]  io_mmioAxi_rd_bits_id, // @[playground/src/noop/crossbar.scala 18:16]
  output [63:0] io_mmioAxi_rd_bits_data, // @[playground/src/noop/crossbar.scala 18:16]
  output [1:0]  io_mmioAxi_rd_bits_resp, // @[playground/src/noop/crossbar.scala 18:16]
  output        io_mmioAxi_rd_bits_last, // @[playground/src/noop/crossbar.scala 18:16]
  input         io_outAxi_wa_ready, // @[playground/src/noop/crossbar.scala 18:16]
  output        io_outAxi_wa_valid, // @[playground/src/noop/crossbar.scala 18:16]
  output [3:0]  io_outAxi_wa_bits_id, // @[playground/src/noop/crossbar.scala 18:16]
  output [31:0] io_outAxi_wa_bits_addr, // @[playground/src/noop/crossbar.scala 18:16]
  output [7:0]  io_outAxi_wa_bits_len, // @[playground/src/noop/crossbar.scala 18:16]
  output [2:0]  io_outAxi_wa_bits_size, // @[playground/src/noop/crossbar.scala 18:16]
  output [1:0]  io_outAxi_wa_bits_burst, // @[playground/src/noop/crossbar.scala 18:16]
  input         io_outAxi_wd_ready, // @[playground/src/noop/crossbar.scala 18:16]
  output        io_outAxi_wd_valid, // @[playground/src/noop/crossbar.scala 18:16]
  output [63:0] io_outAxi_wd_bits_data, // @[playground/src/noop/crossbar.scala 18:16]
  output [7:0]  io_outAxi_wd_bits_strb, // @[playground/src/noop/crossbar.scala 18:16]
  output        io_outAxi_wd_bits_last, // @[playground/src/noop/crossbar.scala 18:16]
  output        io_outAxi_wr_ready, // @[playground/src/noop/crossbar.scala 18:16]
  input         io_outAxi_wr_valid, // @[playground/src/noop/crossbar.scala 18:16]
  input  [3:0]  io_outAxi_wr_bits_id, // @[playground/src/noop/crossbar.scala 18:16]
  input  [1:0]  io_outAxi_wr_bits_resp, // @[playground/src/noop/crossbar.scala 18:16]
  input         io_outAxi_ra_ready, // @[playground/src/noop/crossbar.scala 18:16]
  output        io_outAxi_ra_valid, // @[playground/src/noop/crossbar.scala 18:16]
  output [3:0]  io_outAxi_ra_bits_id, // @[playground/src/noop/crossbar.scala 18:16]
  output [31:0] io_outAxi_ra_bits_addr, // @[playground/src/noop/crossbar.scala 18:16]
  output [7:0]  io_outAxi_ra_bits_len, // @[playground/src/noop/crossbar.scala 18:16]
  output [2:0]  io_outAxi_ra_bits_size, // @[playground/src/noop/crossbar.scala 18:16]
  output [1:0]  io_outAxi_ra_bits_burst, // @[playground/src/noop/crossbar.scala 18:16]
  output        io_outAxi_rd_ready, // @[playground/src/noop/crossbar.scala 18:16]
  input         io_outAxi_rd_valid, // @[playground/src/noop/crossbar.scala 18:16]
  input  [3:0]  io_outAxi_rd_bits_id, // @[playground/src/noop/crossbar.scala 18:16]
  input  [63:0] io_outAxi_rd_bits_data, // @[playground/src/noop/crossbar.scala 18:16]
  input  [1:0]  io_outAxi_rd_bits_resp, // @[playground/src/noop/crossbar.scala 18:16]
  input         io_outAxi_rd_bits_last, // @[playground/src/noop/crossbar.scala 18:16]
  input         io_selectMem // @[playground/src/noop/crossbar.scala 18:16]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg [3:0] state; // @[playground/src/noop/crossbar.scala 20:24]
  reg  selectMem_r; // @[playground/src/noop/crossbar.scala 22:30]
  wire  memTrans = io_memAxi_ra_valid & io_memAxi_ra_ready | io_memAxi_wa_valid & io_memAxi_wa_ready; // @[playground/src/noop/crossbar.scala 31:63]
  wire  memDone = io_memAxi_rd_valid & io_memAxi_rd_bits_last | io_memAxi_wd_valid & io_memAxi_wd_ready &
    io_memAxi_wd_bits_last; // @[playground/src/noop/crossbar.scala 32:88]
  wire  instTrans = io_icAxi_ra_valid & io_icAxi_ra_ready; // @[playground/src/noop/crossbar.scala 33:40]
  wire  instDone = io_icAxi_rd_valid & io_icAxi_rd_bits_last; // @[playground/src/noop/crossbar.scala 34:60]
  wire  flashTrans = io_flashAxi_ra_valid & io_flashAxi_ra_ready; // @[playground/src/noop/crossbar.scala 35:44]
  wire  flashDone = io_flashAxi_rd_valid & io_flashAxi_rd_ready & io_flashAxi_rd_bits_last; // @[playground/src/noop/crossbar.scala 36:67]
  wire  mmioTrans = io_mmioAxi_ra_valid & io_mmioAxi_ra_ready | io_mmioAxi_wa_valid & io_mmioAxi_wa_ready; // @[playground/src/noop/crossbar.scala 37:67]
  wire  mmioDone = io_mmioAxi_rd_valid & io_mmioAxi_rd_ready & io_mmioAxi_rd_bits_last | io_mmioAxi_wd_valid &
    io_mmioAxi_wd_ready & io_mmioAxi_wd_bits_last; // @[playground/src/noop/crossbar.scala 38:93]
  wire [3:0] _GEN_0 = io_icAxi_ra_valid ? 4'h2 : state; // @[playground/src/noop/crossbar.scala 51:42 52:23 20:24]
  wire [3:0] _GEN_1 = io_flashAxi_ra_valid ? 4'h5 : _GEN_0; // @[playground/src/noop/crossbar.scala 49:45 50:23]
  wire [3:0] _GEN_2 = io_mmioAxi_ra_valid | io_mmioAxi_wa_valid ? 4'h7 : _GEN_1; // @[playground/src/noop/crossbar.scala 47:67 48:23]
  wire  _GEN_5 = io_selectMem | selectMem_r; // @[playground/src/noop/crossbar.scala 42:31 44:29 22:30]
  wire [3:0] _GEN_6 = memTrans ? 4'h3 : state; // @[playground/src/noop/crossbar.scala 20:24 61:31 62:27]
  wire  _GEN_9 = selectMem_r & ~io_selectMem ? 1'h0 : 1'h1; // @[playground/src/noop/crossbar.scala 56:47 playground/src/axi/axi.scala 87:18 playground/src/noop/crossbar.scala 60:27]
  wire  _GEN_10 = selectMem_r & ~io_selectMem ? 1'h0 : io_outAxi_rd_valid; // @[playground/src/axi/axi.scala 105:18 playground/src/noop/crossbar.scala 56:47 60:27]
  wire [63:0] _GEN_12 = selectMem_r & ~io_selectMem ? 64'h0 : io_outAxi_rd_bits_data; // @[playground/src/noop/crossbar.scala 56:47 playground/src/axi/axi.scala 68:23 playground/src/noop/crossbar.scala 60:27]
  wire  _GEN_14 = selectMem_r & ~io_selectMem ? 1'h0 : io_outAxi_rd_bits_last; // @[playground/src/noop/crossbar.scala 56:47 playground/src/axi/axi.scala 68:23 playground/src/noop/crossbar.scala 60:27]
  wire  _GEN_15 = selectMem_r & ~io_selectMem ? 1'h0 : io_outAxi_ra_ready; // @[playground/src/axi/axi.scala 104:18 playground/src/noop/crossbar.scala 56:47 60:27]
  wire  _GEN_16 = selectMem_r & ~io_selectMem ? 1'h0 : io_memAxi_ra_valid; // @[playground/src/noop/crossbar.scala 56:47 playground/src/axi/axi.scala 86:18 playground/src/noop/crossbar.scala 60:27]
  wire [31:0] _GEN_18 = selectMem_r & ~io_selectMem ? 32'h0 : io_memAxi_ra_bits_addr; // @[playground/src/axi/axi.scala 41:23 playground/src/noop/crossbar.scala 56:47 60:27]
  wire [7:0] _GEN_19 = selectMem_r & ~io_selectMem ? 8'h0 : 8'h7; // @[playground/src/axi/axi.scala 41:23 playground/src/noop/crossbar.scala 56:47 60:27]
  wire [2:0] _GEN_20 = selectMem_r & ~io_selectMem ? 3'h0 : 3'h3; // @[playground/src/axi/axi.scala 41:23 playground/src/noop/crossbar.scala 56:47 60:27]
  wire [1:0] _GEN_21 = selectMem_r & ~io_selectMem ? 2'h0 : 2'h1; // @[playground/src/axi/axi.scala 41:23 playground/src/noop/crossbar.scala 56:47 60:27]
  wire  _GEN_26 = selectMem_r & ~io_selectMem ? 1'h0 : io_outAxi_wd_ready; // @[playground/src/axi/axi.scala 102:18 playground/src/noop/crossbar.scala 56:47 60:27]
  wire  _GEN_27 = selectMem_r & ~io_selectMem ? 1'h0 : io_memAxi_wd_valid; // @[playground/src/noop/crossbar.scala 56:47 playground/src/axi/axi.scala 84:18 playground/src/noop/crossbar.scala 60:27]
  wire [63:0] _GEN_28 = selectMem_r & ~io_selectMem ? 64'h0 : io_memAxi_wd_bits_data; // @[playground/src/axi/axi.scala 50:23 playground/src/noop/crossbar.scala 56:47 60:27]
  wire [7:0] _GEN_29 = selectMem_r & ~io_selectMem ? 8'h0 : 8'hff; // @[playground/src/axi/axi.scala 50:23 playground/src/noop/crossbar.scala 56:47 60:27]
  wire  _GEN_30 = selectMem_r & ~io_selectMem ? 1'h0 : io_memAxi_wd_bits_last; // @[playground/src/axi/axi.scala 50:23 playground/src/noop/crossbar.scala 56:47 60:27]
  wire  _GEN_31 = selectMem_r & ~io_selectMem ? 1'h0 : io_outAxi_wa_ready; // @[playground/src/axi/axi.scala 101:18 playground/src/noop/crossbar.scala 56:47 60:27]
  wire  _GEN_32 = selectMem_r & ~io_selectMem ? 1'h0 : io_memAxi_wa_valid; // @[playground/src/noop/crossbar.scala 56:47 playground/src/axi/axi.scala 83:18 playground/src/noop/crossbar.scala 60:27]
  wire [31:0] _GEN_34 = selectMem_r & ~io_selectMem ? 32'h0 : io_memAxi_wa_bits_addr; // @[playground/src/axi/axi.scala 41:23 playground/src/noop/crossbar.scala 56:47 60:27]
  wire [3:0] _GEN_38 = memDone ? 4'h0 : state; // @[playground/src/noop/crossbar.scala 68:26 69:23 20:24]
  wire  _GEN_39 = memDone ? 1'h0 : selectMem_r; // @[playground/src/noop/crossbar.scala 68:26 70:29 22:30]
  wire [3:0] _GEN_40 = instTrans ? 4'h4 : state; // @[playground/src/noop/crossbar.scala 75:28 76:23 20:24]
  wire [3:0] _GEN_41 = instDone ? 4'h0 : state; // @[playground/src/noop/crossbar.scala 81:27 82:23 20:24]
  wire [3:0] _GEN_42 = flashTrans ? 4'h6 : state; // @[playground/src/noop/crossbar.scala 87:29 88:23 20:24]
  wire [3:0] _GEN_43 = flashDone ? 4'h0 : state; // @[playground/src/noop/crossbar.scala 93:28 94:23 20:24]
  wire [3:0] _GEN_44 = mmioTrans ? 4'h8 : state; // @[playground/src/noop/crossbar.scala 100:23 20:24 99:28]
  wire [3:0] _GEN_45 = mmioDone ? 4'h0 : state; // @[playground/src/noop/crossbar.scala 105:27 106:23 20:24]
  wire  _GEN_46 = 4'h8 == state & io_mmioAxi_rd_ready; // @[playground/src/noop/crossbar.scala 40:18 104:23 playground/src/axi/axi.scala 87:18]
  wire  _GEN_47 = 4'h8 == state & io_outAxi_rd_valid; // @[playground/src/noop/crossbar.scala 40:18 104:23 playground/src/axi/axi.scala 105:18]
  wire [3:0] _GEN_48 = 4'h8 == state ? io_outAxi_rd_bits_id : 4'h0; // @[playground/src/noop/crossbar.scala 40:18 104:23 playground/src/axi/axi.scala 68:23]
  wire [63:0] _GEN_49 = 4'h8 == state ? io_outAxi_rd_bits_data : 64'h0; // @[playground/src/noop/crossbar.scala 40:18 104:23 playground/src/axi/axi.scala 68:23]
  wire [1:0] _GEN_50 = 4'h8 == state ? io_outAxi_rd_bits_resp : 2'h0; // @[playground/src/noop/crossbar.scala 40:18 104:23 playground/src/axi/axi.scala 68:23]
  wire  _GEN_51 = 4'h8 == state & io_outAxi_rd_bits_last; // @[playground/src/noop/crossbar.scala 40:18 104:23 playground/src/axi/axi.scala 68:23]
  wire  _GEN_52 = 4'h8 == state & io_outAxi_ra_ready; // @[playground/src/axi/axi.scala 104:18 playground/src/noop/crossbar.scala 40:18 104:23]
  wire  _GEN_53 = 4'h8 == state & io_mmioAxi_ra_valid; // @[playground/src/noop/crossbar.scala 40:18 104:23 playground/src/axi/axi.scala 86:18]
  wire [3:0] _GEN_54 = 4'h8 == state ? io_mmioAxi_ra_bits_id : 4'h0; // @[playground/src/noop/crossbar.scala 40:18 104:23 playground/src/axi/axi.scala 41:23]
  wire [31:0] _GEN_55 = 4'h8 == state ? io_mmioAxi_ra_bits_addr : 32'h0; // @[playground/src/noop/crossbar.scala 40:18 104:23 playground/src/axi/axi.scala 41:23]
  wire [7:0] _GEN_56 = 4'h8 == state ? io_mmioAxi_ra_bits_len : 8'h0; // @[playground/src/noop/crossbar.scala 40:18 104:23 playground/src/axi/axi.scala 41:23]
  wire [2:0] _GEN_57 = 4'h8 == state ? io_mmioAxi_ra_bits_size : 3'h0; // @[playground/src/noop/crossbar.scala 40:18 104:23 playground/src/axi/axi.scala 41:23]
  wire [1:0] _GEN_58 = 4'h8 == state ? io_mmioAxi_ra_bits_burst : 2'h0; // @[playground/src/noop/crossbar.scala 40:18 104:23 playground/src/axi/axi.scala 41:23]
  wire  _GEN_59 = 4'h8 == state ? io_mmioAxi_wr_ready : 1'h1; // @[playground/src/noop/crossbar.scala 40:18 104:23 29:24]
  wire  _GEN_60 = 4'h8 == state & io_outAxi_wr_valid; // @[playground/src/axi/axi.scala 103:18 playground/src/noop/crossbar.scala 40:18 104:23]
  wire [3:0] _GEN_61 = 4'h8 == state ? io_outAxi_wr_bits_id : 4'h0; // @[playground/src/noop/crossbar.scala 40:18 104:23 playground/src/axi/axi.scala 58:23]
  wire [1:0] _GEN_62 = 4'h8 == state ? io_outAxi_wr_bits_resp : 2'h0; // @[playground/src/noop/crossbar.scala 40:18 104:23 playground/src/axi/axi.scala 58:23]
  wire  _GEN_63 = 4'h8 == state & io_outAxi_wd_ready; // @[playground/src/axi/axi.scala 102:18 playground/src/noop/crossbar.scala 40:18 104:23]
  wire  _GEN_64 = 4'h8 == state & io_mmioAxi_wd_valid; // @[playground/src/noop/crossbar.scala 40:18 104:23 playground/src/axi/axi.scala 84:18]
  wire [63:0] _GEN_65 = 4'h8 == state ? io_mmioAxi_wd_bits_data : 64'h0; // @[playground/src/noop/crossbar.scala 40:18 104:23 playground/src/axi/axi.scala 50:23]
  wire [7:0] _GEN_66 = 4'h8 == state ? io_mmioAxi_wd_bits_strb : 8'h0; // @[playground/src/noop/crossbar.scala 40:18 104:23 playground/src/axi/axi.scala 50:23]
  wire  _GEN_67 = 4'h8 == state & io_mmioAxi_wd_bits_last; // @[playground/src/noop/crossbar.scala 40:18 104:23 playground/src/axi/axi.scala 50:23]
  wire  _GEN_68 = 4'h8 == state & io_outAxi_wa_ready; // @[playground/src/axi/axi.scala 101:18 playground/src/noop/crossbar.scala 40:18 104:23]
  wire  _GEN_69 = 4'h8 == state & io_mmioAxi_wa_valid; // @[playground/src/noop/crossbar.scala 40:18 104:23 playground/src/axi/axi.scala 83:18]
  wire [3:0] _GEN_70 = 4'h8 == state ? io_mmioAxi_wa_bits_id : 4'h0; // @[playground/src/noop/crossbar.scala 40:18 104:23 playground/src/axi/axi.scala 41:23]
  wire [31:0] _GEN_71 = 4'h8 == state ? io_mmioAxi_wa_bits_addr : 32'h0; // @[playground/src/noop/crossbar.scala 40:18 104:23 playground/src/axi/axi.scala 41:23]
  wire [7:0] _GEN_72 = 4'h8 == state ? io_mmioAxi_wa_bits_len : 8'h0; // @[playground/src/noop/crossbar.scala 40:18 104:23 playground/src/axi/axi.scala 41:23]
  wire [2:0] _GEN_73 = 4'h8 == state ? io_mmioAxi_wa_bits_size : 3'h0; // @[playground/src/noop/crossbar.scala 40:18 104:23 playground/src/axi/axi.scala 41:23]
  wire [1:0] _GEN_74 = 4'h8 == state ? io_mmioAxi_wa_bits_burst : 2'h0; // @[playground/src/noop/crossbar.scala 40:18 104:23 playground/src/axi/axi.scala 41:23]
  wire [3:0] _GEN_75 = 4'h8 == state ? _GEN_45 : state; // @[playground/src/noop/crossbar.scala 40:18 20:24]
  wire  _GEN_76 = 4'h7 == state ? io_mmioAxi_rd_ready : _GEN_46; // @[playground/src/noop/crossbar.scala 40:18 98:23]
  wire  _GEN_77 = 4'h7 == state ? io_outAxi_rd_valid : _GEN_47; // @[playground/src/noop/crossbar.scala 40:18 98:23]
  wire [3:0] _GEN_78 = 4'h7 == state ? io_outAxi_rd_bits_id : _GEN_48; // @[playground/src/noop/crossbar.scala 40:18 98:23]
  wire [63:0] _GEN_79 = 4'h7 == state ? io_outAxi_rd_bits_data : _GEN_49; // @[playground/src/noop/crossbar.scala 40:18 98:23]
  wire [1:0] _GEN_80 = 4'h7 == state ? io_outAxi_rd_bits_resp : _GEN_50; // @[playground/src/noop/crossbar.scala 40:18 98:23]
  wire  _GEN_81 = 4'h7 == state ? io_outAxi_rd_bits_last : _GEN_51; // @[playground/src/noop/crossbar.scala 40:18 98:23]
  wire  _GEN_82 = 4'h7 == state ? io_outAxi_ra_ready : _GEN_52; // @[playground/src/noop/crossbar.scala 40:18 98:23]
  wire  _GEN_83 = 4'h7 == state ? io_mmioAxi_ra_valid : _GEN_53; // @[playground/src/noop/crossbar.scala 40:18 98:23]
  wire [3:0] _GEN_84 = 4'h7 == state ? io_mmioAxi_ra_bits_id : _GEN_54; // @[playground/src/noop/crossbar.scala 40:18 98:23]
  wire [31:0] _GEN_85 = 4'h7 == state ? io_mmioAxi_ra_bits_addr : _GEN_55; // @[playground/src/noop/crossbar.scala 40:18 98:23]
  wire [7:0] _GEN_86 = 4'h7 == state ? io_mmioAxi_ra_bits_len : _GEN_56; // @[playground/src/noop/crossbar.scala 40:18 98:23]
  wire [2:0] _GEN_87 = 4'h7 == state ? io_mmioAxi_ra_bits_size : _GEN_57; // @[playground/src/noop/crossbar.scala 40:18 98:23]
  wire [1:0] _GEN_88 = 4'h7 == state ? io_mmioAxi_ra_bits_burst : _GEN_58; // @[playground/src/noop/crossbar.scala 40:18 98:23]
  wire  _GEN_89 = 4'h7 == state ? io_mmioAxi_wr_ready : _GEN_59; // @[playground/src/noop/crossbar.scala 40:18 98:23]
  wire  _GEN_90 = 4'h7 == state ? io_outAxi_wr_valid : _GEN_60; // @[playground/src/noop/crossbar.scala 40:18 98:23]
  wire [3:0] _GEN_91 = 4'h7 == state ? io_outAxi_wr_bits_id : _GEN_61; // @[playground/src/noop/crossbar.scala 40:18 98:23]
  wire [1:0] _GEN_92 = 4'h7 == state ? io_outAxi_wr_bits_resp : _GEN_62; // @[playground/src/noop/crossbar.scala 40:18 98:23]
  wire  _GEN_93 = 4'h7 == state ? io_outAxi_wd_ready : _GEN_63; // @[playground/src/noop/crossbar.scala 40:18 98:23]
  wire  _GEN_94 = 4'h7 == state ? io_mmioAxi_wd_valid : _GEN_64; // @[playground/src/noop/crossbar.scala 40:18 98:23]
  wire [63:0] _GEN_95 = 4'h7 == state ? io_mmioAxi_wd_bits_data : _GEN_65; // @[playground/src/noop/crossbar.scala 40:18 98:23]
  wire [7:0] _GEN_96 = 4'h7 == state ? io_mmioAxi_wd_bits_strb : _GEN_66; // @[playground/src/noop/crossbar.scala 40:18 98:23]
  wire  _GEN_97 = 4'h7 == state ? io_mmioAxi_wd_bits_last : _GEN_67; // @[playground/src/noop/crossbar.scala 40:18 98:23]
  wire  _GEN_98 = 4'h7 == state ? io_outAxi_wa_ready : _GEN_68; // @[playground/src/noop/crossbar.scala 40:18 98:23]
  wire  _GEN_99 = 4'h7 == state ? io_mmioAxi_wa_valid : _GEN_69; // @[playground/src/noop/crossbar.scala 40:18 98:23]
  wire [3:0] _GEN_100 = 4'h7 == state ? io_mmioAxi_wa_bits_id : _GEN_70; // @[playground/src/noop/crossbar.scala 40:18 98:23]
  wire [31:0] _GEN_101 = 4'h7 == state ? io_mmioAxi_wa_bits_addr : _GEN_71; // @[playground/src/noop/crossbar.scala 40:18 98:23]
  wire [7:0] _GEN_102 = 4'h7 == state ? io_mmioAxi_wa_bits_len : _GEN_72; // @[playground/src/noop/crossbar.scala 40:18 98:23]
  wire [2:0] _GEN_103 = 4'h7 == state ? io_mmioAxi_wa_bits_size : _GEN_73; // @[playground/src/noop/crossbar.scala 40:18 98:23]
  wire [1:0] _GEN_104 = 4'h7 == state ? io_mmioAxi_wa_bits_burst : _GEN_74; // @[playground/src/noop/crossbar.scala 40:18 98:23]
  wire [3:0] _GEN_105 = 4'h7 == state ? _GEN_44 : _GEN_75; // @[playground/src/noop/crossbar.scala 40:18]
  wire  _GEN_106 = 4'h6 == state ? io_flashAxi_rd_ready : _GEN_76; // @[playground/src/noop/crossbar.scala 40:18 92:23]
  wire  _GEN_107 = 4'h6 == state & io_outAxi_rd_valid; // @[playground/src/axi/axi.scala 105:18 playground/src/noop/crossbar.scala 40:18 92:23]
  wire [3:0] _GEN_108 = 4'h6 == state ? io_outAxi_rd_bits_id : 4'h0; // @[playground/src/noop/crossbar.scala 40:18 playground/src/axi/axi.scala 68:23 playground/src/noop/crossbar.scala 92:23]
  wire [63:0] _GEN_109 = 4'h6 == state ? io_outAxi_rd_bits_data : 64'h0; // @[playground/src/noop/crossbar.scala 40:18 playground/src/axi/axi.scala 68:23 playground/src/noop/crossbar.scala 92:23]
  wire [1:0] _GEN_110 = 4'h6 == state ? io_outAxi_rd_bits_resp : 2'h0; // @[playground/src/noop/crossbar.scala 40:18 playground/src/axi/axi.scala 68:23 playground/src/noop/crossbar.scala 92:23]
  wire  _GEN_111 = 4'h6 == state & io_outAxi_rd_bits_last; // @[playground/src/noop/crossbar.scala 40:18 playground/src/axi/axi.scala 68:23 playground/src/noop/crossbar.scala 92:23]
  wire  _GEN_112 = 4'h6 == state & io_outAxi_ra_ready; // @[playground/src/axi/axi.scala 104:18 playground/src/noop/crossbar.scala 40:18 92:23]
  wire  _GEN_113 = 4'h6 == state ? io_flashAxi_ra_valid : _GEN_83; // @[playground/src/noop/crossbar.scala 40:18 92:23]
  wire [3:0] _GEN_114 = 4'h6 == state ? io_flashAxi_ra_bits_id : _GEN_84; // @[playground/src/noop/crossbar.scala 40:18 92:23]
  wire [31:0] _GEN_115 = 4'h6 == state ? io_flashAxi_ra_bits_addr : _GEN_85; // @[playground/src/noop/crossbar.scala 40:18 92:23]
  wire [7:0] _GEN_116 = 4'h6 == state ? io_flashAxi_ra_bits_len : _GEN_86; // @[playground/src/noop/crossbar.scala 40:18 92:23]
  wire [2:0] _GEN_117 = 4'h6 == state ? io_flashAxi_ra_bits_size : _GEN_87; // @[playground/src/noop/crossbar.scala 40:18 92:23]
  wire [1:0] _GEN_118 = 4'h6 == state ? io_flashAxi_ra_bits_burst : _GEN_88; // @[playground/src/noop/crossbar.scala 40:18 92:23]
  wire  _GEN_119 = 4'h6 == state ? io_flashAxi_wr_ready : _GEN_89; // @[playground/src/noop/crossbar.scala 40:18 92:23]
  wire  _GEN_120 = 4'h6 == state & io_outAxi_wr_valid; // @[playground/src/axi/axi.scala 103:18 playground/src/noop/crossbar.scala 40:18 92:23]
  wire [3:0] _GEN_121 = 4'h6 == state ? io_outAxi_wr_bits_id : 4'h0; // @[playground/src/noop/crossbar.scala 40:18 playground/src/axi/axi.scala 58:23 playground/src/noop/crossbar.scala 92:23]
  wire [1:0] _GEN_122 = 4'h6 == state ? io_outAxi_wr_bits_resp : 2'h0; // @[playground/src/noop/crossbar.scala 40:18 playground/src/axi/axi.scala 58:23 playground/src/noop/crossbar.scala 92:23]
  wire  _GEN_123 = 4'h6 == state & io_outAxi_wd_ready; // @[playground/src/axi/axi.scala 102:18 playground/src/noop/crossbar.scala 40:18 92:23]
  wire  _GEN_124 = 4'h6 == state ? io_flashAxi_wd_valid : _GEN_94; // @[playground/src/noop/crossbar.scala 40:18 92:23]
  wire [63:0] _GEN_125 = 4'h6 == state ? io_flashAxi_wd_bits_data : _GEN_95; // @[playground/src/noop/crossbar.scala 40:18 92:23]
  wire [7:0] _GEN_126 = 4'h6 == state ? io_flashAxi_wd_bits_strb : _GEN_96; // @[playground/src/noop/crossbar.scala 40:18 92:23]
  wire  _GEN_127 = 4'h6 == state ? io_flashAxi_wd_bits_last : _GEN_97; // @[playground/src/noop/crossbar.scala 40:18 92:23]
  wire  _GEN_128 = 4'h6 == state & io_outAxi_wa_ready; // @[playground/src/axi/axi.scala 101:18 playground/src/noop/crossbar.scala 40:18 92:23]
  wire  _GEN_129 = 4'h6 == state ? io_flashAxi_wa_valid : _GEN_99; // @[playground/src/noop/crossbar.scala 40:18 92:23]
  wire [3:0] _GEN_130 = 4'h6 == state ? io_flashAxi_wa_bits_id : _GEN_100; // @[playground/src/noop/crossbar.scala 40:18 92:23]
  wire [31:0] _GEN_131 = 4'h6 == state ? io_flashAxi_wa_bits_addr : _GEN_101; // @[playground/src/noop/crossbar.scala 40:18 92:23]
  wire [7:0] _GEN_132 = 4'h6 == state ? io_flashAxi_wa_bits_len : _GEN_102; // @[playground/src/noop/crossbar.scala 40:18 92:23]
  wire [2:0] _GEN_133 = 4'h6 == state ? io_flashAxi_wa_bits_size : _GEN_103; // @[playground/src/noop/crossbar.scala 40:18 92:23]
  wire [1:0] _GEN_134 = 4'h6 == state ? io_flashAxi_wa_bits_burst : _GEN_104; // @[playground/src/noop/crossbar.scala 40:18 92:23]
  wire [3:0] _GEN_135 = 4'h6 == state ? _GEN_43 : _GEN_105; // @[playground/src/noop/crossbar.scala 40:18]
  wire  _GEN_136 = 4'h6 == state ? 1'h0 : _GEN_77; // @[playground/src/axi/axi.scala 105:18 playground/src/noop/crossbar.scala 40:18]
  wire [3:0] _GEN_137 = 4'h6 == state ? 4'h0 : _GEN_78; // @[playground/src/noop/crossbar.scala 40:18 playground/src/axi/axi.scala 68:23]
  wire [63:0] _GEN_138 = 4'h6 == state ? 64'h0 : _GEN_79; // @[playground/src/noop/crossbar.scala 40:18 playground/src/axi/axi.scala 68:23]
  wire [1:0] _GEN_139 = 4'h6 == state ? 2'h0 : _GEN_80; // @[playground/src/noop/crossbar.scala 40:18 playground/src/axi/axi.scala 68:23]
  wire  _GEN_140 = 4'h6 == state ? 1'h0 : _GEN_81; // @[playground/src/noop/crossbar.scala 40:18 playground/src/axi/axi.scala 68:23]
  wire  _GEN_141 = 4'h6 == state ? 1'h0 : _GEN_82; // @[playground/src/axi/axi.scala 104:18 playground/src/noop/crossbar.scala 40:18]
  wire  _GEN_142 = 4'h6 == state ? 1'h0 : _GEN_90; // @[playground/src/axi/axi.scala 103:18 playground/src/noop/crossbar.scala 40:18]
  wire [3:0] _GEN_143 = 4'h6 == state ? 4'h0 : _GEN_91; // @[playground/src/noop/crossbar.scala 40:18 playground/src/axi/axi.scala 58:23]
  wire [1:0] _GEN_144 = 4'h6 == state ? 2'h0 : _GEN_92; // @[playground/src/noop/crossbar.scala 40:18 playground/src/axi/axi.scala 58:23]
  wire  _GEN_145 = 4'h6 == state ? 1'h0 : _GEN_93; // @[playground/src/axi/axi.scala 102:18 playground/src/noop/crossbar.scala 40:18]
  wire  _GEN_146 = 4'h6 == state ? 1'h0 : _GEN_98; // @[playground/src/axi/axi.scala 101:18 playground/src/noop/crossbar.scala 40:18]
  wire  _GEN_147 = 4'h5 == state ? io_flashAxi_rd_ready : _GEN_106; // @[playground/src/noop/crossbar.scala 40:18 86:23]
  wire  _GEN_148 = 4'h5 == state ? io_outAxi_rd_valid : _GEN_107; // @[playground/src/noop/crossbar.scala 40:18 86:23]
  wire [3:0] _GEN_149 = 4'h5 == state ? io_outAxi_rd_bits_id : _GEN_108; // @[playground/src/noop/crossbar.scala 40:18 86:23]
  wire [63:0] _GEN_150 = 4'h5 == state ? io_outAxi_rd_bits_data : _GEN_109; // @[playground/src/noop/crossbar.scala 40:18 86:23]
  wire [1:0] _GEN_151 = 4'h5 == state ? io_outAxi_rd_bits_resp : _GEN_110; // @[playground/src/noop/crossbar.scala 40:18 86:23]
  wire  _GEN_152 = 4'h5 == state ? io_outAxi_rd_bits_last : _GEN_111; // @[playground/src/noop/crossbar.scala 40:18 86:23]
  wire  _GEN_153 = 4'h5 == state ? io_outAxi_ra_ready : _GEN_112; // @[playground/src/noop/crossbar.scala 40:18 86:23]
  wire  _GEN_154 = 4'h5 == state ? io_flashAxi_ra_valid : _GEN_113; // @[playground/src/noop/crossbar.scala 40:18 86:23]
  wire [3:0] _GEN_155 = 4'h5 == state ? io_flashAxi_ra_bits_id : _GEN_114; // @[playground/src/noop/crossbar.scala 40:18 86:23]
  wire [31:0] _GEN_156 = 4'h5 == state ? io_flashAxi_ra_bits_addr : _GEN_115; // @[playground/src/noop/crossbar.scala 40:18 86:23]
  wire [7:0] _GEN_157 = 4'h5 == state ? io_flashAxi_ra_bits_len : _GEN_116; // @[playground/src/noop/crossbar.scala 40:18 86:23]
  wire [2:0] _GEN_158 = 4'h5 == state ? io_flashAxi_ra_bits_size : _GEN_117; // @[playground/src/noop/crossbar.scala 40:18 86:23]
  wire [1:0] _GEN_159 = 4'h5 == state ? io_flashAxi_ra_bits_burst : _GEN_118; // @[playground/src/noop/crossbar.scala 40:18 86:23]
  wire  _GEN_160 = 4'h5 == state ? io_flashAxi_wr_ready : _GEN_119; // @[playground/src/noop/crossbar.scala 40:18 86:23]
  wire  _GEN_161 = 4'h5 == state ? io_outAxi_wr_valid : _GEN_120; // @[playground/src/noop/crossbar.scala 40:18 86:23]
  wire [3:0] _GEN_162 = 4'h5 == state ? io_outAxi_wr_bits_id : _GEN_121; // @[playground/src/noop/crossbar.scala 40:18 86:23]
  wire [1:0] _GEN_163 = 4'h5 == state ? io_outAxi_wr_bits_resp : _GEN_122; // @[playground/src/noop/crossbar.scala 40:18 86:23]
  wire  _GEN_164 = 4'h5 == state ? io_outAxi_wd_ready : _GEN_123; // @[playground/src/noop/crossbar.scala 40:18 86:23]
  wire  _GEN_165 = 4'h5 == state ? io_flashAxi_wd_valid : _GEN_124; // @[playground/src/noop/crossbar.scala 40:18 86:23]
  wire [63:0] _GEN_166 = 4'h5 == state ? io_flashAxi_wd_bits_data : _GEN_125; // @[playground/src/noop/crossbar.scala 40:18 86:23]
  wire [7:0] _GEN_167 = 4'h5 == state ? io_flashAxi_wd_bits_strb : _GEN_126; // @[playground/src/noop/crossbar.scala 40:18 86:23]
  wire  _GEN_168 = 4'h5 == state ? io_flashAxi_wd_bits_last : _GEN_127; // @[playground/src/noop/crossbar.scala 40:18 86:23]
  wire  _GEN_169 = 4'h5 == state ? io_outAxi_wa_ready : _GEN_128; // @[playground/src/noop/crossbar.scala 40:18 86:23]
  wire  _GEN_170 = 4'h5 == state ? io_flashAxi_wa_valid : _GEN_129; // @[playground/src/noop/crossbar.scala 40:18 86:23]
  wire [3:0] _GEN_171 = 4'h5 == state ? io_flashAxi_wa_bits_id : _GEN_130; // @[playground/src/noop/crossbar.scala 40:18 86:23]
  wire [31:0] _GEN_172 = 4'h5 == state ? io_flashAxi_wa_bits_addr : _GEN_131; // @[playground/src/noop/crossbar.scala 40:18 86:23]
  wire [7:0] _GEN_173 = 4'h5 == state ? io_flashAxi_wa_bits_len : _GEN_132; // @[playground/src/noop/crossbar.scala 40:18 86:23]
  wire [2:0] _GEN_174 = 4'h5 == state ? io_flashAxi_wa_bits_size : _GEN_133; // @[playground/src/noop/crossbar.scala 40:18 86:23]
  wire [1:0] _GEN_175 = 4'h5 == state ? io_flashAxi_wa_bits_burst : _GEN_134; // @[playground/src/noop/crossbar.scala 40:18 86:23]
  wire [3:0] _GEN_176 = 4'h5 == state ? _GEN_42 : _GEN_135; // @[playground/src/noop/crossbar.scala 40:18]
  wire  _GEN_177 = 4'h5 == state ? 1'h0 : _GEN_136; // @[playground/src/axi/axi.scala 105:18 playground/src/noop/crossbar.scala 40:18]
  wire [3:0] _GEN_178 = 4'h5 == state ? 4'h0 : _GEN_137; // @[playground/src/noop/crossbar.scala 40:18 playground/src/axi/axi.scala 68:23]
  wire [63:0] _GEN_179 = 4'h5 == state ? 64'h0 : _GEN_138; // @[playground/src/noop/crossbar.scala 40:18 playground/src/axi/axi.scala 68:23]
  wire [1:0] _GEN_180 = 4'h5 == state ? 2'h0 : _GEN_139; // @[playground/src/noop/crossbar.scala 40:18 playground/src/axi/axi.scala 68:23]
  wire  _GEN_181 = 4'h5 == state ? 1'h0 : _GEN_140; // @[playground/src/noop/crossbar.scala 40:18 playground/src/axi/axi.scala 68:23]
  wire  _GEN_182 = 4'h5 == state ? 1'h0 : _GEN_141; // @[playground/src/axi/axi.scala 104:18 playground/src/noop/crossbar.scala 40:18]
  wire  _GEN_183 = 4'h5 == state ? 1'h0 : _GEN_142; // @[playground/src/axi/axi.scala 103:18 playground/src/noop/crossbar.scala 40:18]
  wire [3:0] _GEN_184 = 4'h5 == state ? 4'h0 : _GEN_143; // @[playground/src/noop/crossbar.scala 40:18 playground/src/axi/axi.scala 58:23]
  wire [1:0] _GEN_185 = 4'h5 == state ? 2'h0 : _GEN_144; // @[playground/src/noop/crossbar.scala 40:18 playground/src/axi/axi.scala 58:23]
  wire  _GEN_186 = 4'h5 == state ? 1'h0 : _GEN_145; // @[playground/src/axi/axi.scala 102:18 playground/src/noop/crossbar.scala 40:18]
  wire  _GEN_187 = 4'h5 == state ? 1'h0 : _GEN_146; // @[playground/src/axi/axi.scala 101:18 playground/src/noop/crossbar.scala 40:18]
  wire  _GEN_188 = 4'h4 == state | _GEN_147; // @[playground/src/noop/crossbar.scala 40:18 80:23]
  wire  _GEN_189 = 4'h4 == state & io_outAxi_rd_valid; // @[playground/src/axi/axi.scala 105:18 playground/src/noop/crossbar.scala 40:18 80:23]
  wire [63:0] _GEN_191 = 4'h4 == state ? io_outAxi_rd_bits_data : 64'h0; // @[playground/src/noop/crossbar.scala 40:18 playground/src/axi/axi.scala 68:23 playground/src/noop/crossbar.scala 80:23]
  wire  _GEN_193 = 4'h4 == state & io_outAxi_rd_bits_last; // @[playground/src/noop/crossbar.scala 40:18 playground/src/axi/axi.scala 68:23 playground/src/noop/crossbar.scala 80:23]
  wire  _GEN_194 = 4'h4 == state & io_outAxi_ra_ready; // @[playground/src/axi/axi.scala 104:18 playground/src/noop/crossbar.scala 40:18 80:23]
  wire  _GEN_195 = 4'h4 == state ? io_icAxi_ra_valid : _GEN_154; // @[playground/src/noop/crossbar.scala 40:18 80:23]
  wire [3:0] _GEN_196 = 4'h4 == state ? 4'h0 : _GEN_155; // @[playground/src/noop/crossbar.scala 40:18 80:23]
  wire [31:0] _GEN_197 = 4'h4 == state ? io_icAxi_ra_bits_addr : _GEN_156; // @[playground/src/noop/crossbar.scala 40:18 80:23]
  wire [7:0] _GEN_198 = 4'h4 == state ? 8'h7 : _GEN_157; // @[playground/src/noop/crossbar.scala 40:18 80:23]
  wire [2:0] _GEN_199 = 4'h4 == state ? 3'h3 : _GEN_158; // @[playground/src/noop/crossbar.scala 40:18 80:23]
  wire [1:0] _GEN_200 = 4'h4 == state ? 2'h1 : _GEN_159; // @[playground/src/noop/crossbar.scala 40:18 80:23]
  wire  _GEN_201 = 4'h4 == state | _GEN_160; // @[playground/src/noop/crossbar.scala 40:18 80:23]
  wire  _GEN_206 = 4'h4 == state ? 1'h0 : _GEN_165; // @[playground/src/noop/crossbar.scala 40:18 80:23]
  wire [63:0] _GEN_207 = 4'h4 == state ? 64'h0 : _GEN_166; // @[playground/src/noop/crossbar.scala 40:18 80:23]
  wire [7:0] _GEN_208 = 4'h4 == state ? 8'h0 : _GEN_167; // @[playground/src/noop/crossbar.scala 40:18 80:23]
  wire  _GEN_209 = 4'h4 == state ? 1'h0 : _GEN_168; // @[playground/src/noop/crossbar.scala 40:18 80:23]
  wire  _GEN_211 = 4'h4 == state ? 1'h0 : _GEN_170; // @[playground/src/noop/crossbar.scala 40:18 80:23]
  wire [3:0] _GEN_212 = 4'h4 == state ? 4'h0 : _GEN_171; // @[playground/src/noop/crossbar.scala 40:18 80:23]
  wire [31:0] _GEN_213 = 4'h4 == state ? 32'h0 : _GEN_172; // @[playground/src/noop/crossbar.scala 40:18 80:23]
  wire [7:0] _GEN_214 = 4'h4 == state ? 8'h0 : _GEN_173; // @[playground/src/noop/crossbar.scala 40:18 80:23]
  wire [2:0] _GEN_215 = 4'h4 == state ? 3'h0 : _GEN_174; // @[playground/src/noop/crossbar.scala 40:18 80:23]
  wire [1:0] _GEN_216 = 4'h4 == state ? 2'h0 : _GEN_175; // @[playground/src/noop/crossbar.scala 40:18 80:23]
  wire [3:0] _GEN_217 = 4'h4 == state ? _GEN_41 : _GEN_176; // @[playground/src/noop/crossbar.scala 40:18]
  wire  _GEN_218 = 4'h4 == state ? 1'h0 : _GEN_148; // @[playground/src/axi/axi.scala 105:18 playground/src/noop/crossbar.scala 40:18]
  wire [3:0] _GEN_219 = 4'h4 == state ? 4'h0 : _GEN_149; // @[playground/src/noop/crossbar.scala 40:18 playground/src/axi/axi.scala 68:23]
  wire [63:0] _GEN_220 = 4'h4 == state ? 64'h0 : _GEN_150; // @[playground/src/noop/crossbar.scala 40:18 playground/src/axi/axi.scala 68:23]
  wire [1:0] _GEN_221 = 4'h4 == state ? 2'h0 : _GEN_151; // @[playground/src/noop/crossbar.scala 40:18 playground/src/axi/axi.scala 68:23]
  wire  _GEN_222 = 4'h4 == state ? 1'h0 : _GEN_152; // @[playground/src/noop/crossbar.scala 40:18 playground/src/axi/axi.scala 68:23]
  wire  _GEN_223 = 4'h4 == state ? 1'h0 : _GEN_153; // @[playground/src/axi/axi.scala 104:18 playground/src/noop/crossbar.scala 40:18]
  wire  _GEN_224 = 4'h4 == state ? 1'h0 : _GEN_161; // @[playground/src/axi/axi.scala 103:18 playground/src/noop/crossbar.scala 40:18]
  wire [3:0] _GEN_225 = 4'h4 == state ? 4'h0 : _GEN_162; // @[playground/src/noop/crossbar.scala 40:18 playground/src/axi/axi.scala 58:23]
  wire [1:0] _GEN_226 = 4'h4 == state ? 2'h0 : _GEN_163; // @[playground/src/noop/crossbar.scala 40:18 playground/src/axi/axi.scala 58:23]
  wire  _GEN_227 = 4'h4 == state ? 1'h0 : _GEN_164; // @[playground/src/axi/axi.scala 102:18 playground/src/noop/crossbar.scala 40:18]
  wire  _GEN_228 = 4'h4 == state ? 1'h0 : _GEN_169; // @[playground/src/axi/axi.scala 101:18 playground/src/noop/crossbar.scala 40:18]
  wire  _GEN_229 = 4'h4 == state ? 1'h0 : _GEN_177; // @[playground/src/axi/axi.scala 105:18 playground/src/noop/crossbar.scala 40:18]
  wire [3:0] _GEN_230 = 4'h4 == state ? 4'h0 : _GEN_178; // @[playground/src/noop/crossbar.scala 40:18 playground/src/axi/axi.scala 68:23]
  wire [63:0] _GEN_231 = 4'h4 == state ? 64'h0 : _GEN_179; // @[playground/src/noop/crossbar.scala 40:18 playground/src/axi/axi.scala 68:23]
  wire [1:0] _GEN_232 = 4'h4 == state ? 2'h0 : _GEN_180; // @[playground/src/noop/crossbar.scala 40:18 playground/src/axi/axi.scala 68:23]
  wire  _GEN_233 = 4'h4 == state ? 1'h0 : _GEN_181; // @[playground/src/noop/crossbar.scala 40:18 playground/src/axi/axi.scala 68:23]
  wire  _GEN_234 = 4'h4 == state ? 1'h0 : _GEN_182; // @[playground/src/axi/axi.scala 104:18 playground/src/noop/crossbar.scala 40:18]
  wire  _GEN_235 = 4'h4 == state ? 1'h0 : _GEN_183; // @[playground/src/axi/axi.scala 103:18 playground/src/noop/crossbar.scala 40:18]
  wire [3:0] _GEN_236 = 4'h4 == state ? 4'h0 : _GEN_184; // @[playground/src/noop/crossbar.scala 40:18 playground/src/axi/axi.scala 58:23]
  wire [1:0] _GEN_237 = 4'h4 == state ? 2'h0 : _GEN_185; // @[playground/src/noop/crossbar.scala 40:18 playground/src/axi/axi.scala 58:23]
  wire  _GEN_238 = 4'h4 == state ? 1'h0 : _GEN_186; // @[playground/src/axi/axi.scala 102:18 playground/src/noop/crossbar.scala 40:18]
  wire  _GEN_239 = 4'h4 == state ? 1'h0 : _GEN_187; // @[playground/src/axi/axi.scala 101:18 playground/src/noop/crossbar.scala 40:18]
  wire  _GEN_240 = 4'h2 == state | _GEN_188; // @[playground/src/noop/crossbar.scala 40:18 74:23]
  wire  _GEN_241 = 4'h2 == state ? io_outAxi_rd_valid : _GEN_189; // @[playground/src/noop/crossbar.scala 40:18 74:23]
  wire [63:0] _GEN_243 = 4'h2 == state ? io_outAxi_rd_bits_data : _GEN_191; // @[playground/src/noop/crossbar.scala 40:18 74:23]
  wire  _GEN_245 = 4'h2 == state ? io_outAxi_rd_bits_last : _GEN_193; // @[playground/src/noop/crossbar.scala 40:18 74:23]
  wire  _GEN_246 = 4'h2 == state ? io_outAxi_ra_ready : _GEN_194; // @[playground/src/noop/crossbar.scala 40:18 74:23]
  wire  _GEN_247 = 4'h2 == state ? io_icAxi_ra_valid : _GEN_195; // @[playground/src/noop/crossbar.scala 40:18 74:23]
  wire [3:0] _GEN_248 = 4'h2 == state ? 4'h0 : _GEN_196; // @[playground/src/noop/crossbar.scala 40:18 74:23]
  wire [31:0] _GEN_249 = 4'h2 == state ? io_icAxi_ra_bits_addr : _GEN_197; // @[playground/src/noop/crossbar.scala 40:18 74:23]
  wire [7:0] _GEN_250 = 4'h2 == state ? 8'h7 : _GEN_198; // @[playground/src/noop/crossbar.scala 40:18 74:23]
  wire [2:0] _GEN_251 = 4'h2 == state ? 3'h3 : _GEN_199; // @[playground/src/noop/crossbar.scala 40:18 74:23]
  wire [1:0] _GEN_252 = 4'h2 == state ? 2'h1 : _GEN_200; // @[playground/src/noop/crossbar.scala 40:18 74:23]
  wire  _GEN_253 = 4'h2 == state | _GEN_201; // @[playground/src/noop/crossbar.scala 40:18 74:23]
  wire  _GEN_258 = 4'h2 == state ? 1'h0 : _GEN_206; // @[playground/src/noop/crossbar.scala 40:18 74:23]
  wire [63:0] _GEN_259 = 4'h2 == state ? 64'h0 : _GEN_207; // @[playground/src/noop/crossbar.scala 40:18 74:23]
  wire [7:0] _GEN_260 = 4'h2 == state ? 8'h0 : _GEN_208; // @[playground/src/noop/crossbar.scala 40:18 74:23]
  wire  _GEN_261 = 4'h2 == state ? 1'h0 : _GEN_209; // @[playground/src/noop/crossbar.scala 40:18 74:23]
  wire  _GEN_263 = 4'h2 == state ? 1'h0 : _GEN_211; // @[playground/src/noop/crossbar.scala 40:18 74:23]
  wire [3:0] _GEN_264 = 4'h2 == state ? 4'h0 : _GEN_212; // @[playground/src/noop/crossbar.scala 40:18 74:23]
  wire [31:0] _GEN_265 = 4'h2 == state ? 32'h0 : _GEN_213; // @[playground/src/noop/crossbar.scala 40:18 74:23]
  wire [7:0] _GEN_266 = 4'h2 == state ? 8'h0 : _GEN_214; // @[playground/src/noop/crossbar.scala 40:18 74:23]
  wire [2:0] _GEN_267 = 4'h2 == state ? 3'h0 : _GEN_215; // @[playground/src/noop/crossbar.scala 40:18 74:23]
  wire [1:0] _GEN_268 = 4'h2 == state ? 2'h0 : _GEN_216; // @[playground/src/noop/crossbar.scala 40:18 74:23]
  wire [3:0] _GEN_269 = 4'h2 == state ? _GEN_40 : _GEN_217; // @[playground/src/noop/crossbar.scala 40:18]
  wire  _GEN_270 = 4'h2 == state ? 1'h0 : _GEN_218; // @[playground/src/axi/axi.scala 105:18 playground/src/noop/crossbar.scala 40:18]
  wire [3:0] _GEN_271 = 4'h2 == state ? 4'h0 : _GEN_219; // @[playground/src/noop/crossbar.scala 40:18 playground/src/axi/axi.scala 68:23]
  wire [63:0] _GEN_272 = 4'h2 == state ? 64'h0 : _GEN_220; // @[playground/src/noop/crossbar.scala 40:18 playground/src/axi/axi.scala 68:23]
  wire [1:0] _GEN_273 = 4'h2 == state ? 2'h0 : _GEN_221; // @[playground/src/noop/crossbar.scala 40:18 playground/src/axi/axi.scala 68:23]
  wire  _GEN_274 = 4'h2 == state ? 1'h0 : _GEN_222; // @[playground/src/noop/crossbar.scala 40:18 playground/src/axi/axi.scala 68:23]
  wire  _GEN_275 = 4'h2 == state ? 1'h0 : _GEN_223; // @[playground/src/axi/axi.scala 104:18 playground/src/noop/crossbar.scala 40:18]
  wire  _GEN_276 = 4'h2 == state ? 1'h0 : _GEN_224; // @[playground/src/axi/axi.scala 103:18 playground/src/noop/crossbar.scala 40:18]
  wire [3:0] _GEN_277 = 4'h2 == state ? 4'h0 : _GEN_225; // @[playground/src/noop/crossbar.scala 40:18 playground/src/axi/axi.scala 58:23]
  wire [1:0] _GEN_278 = 4'h2 == state ? 2'h0 : _GEN_226; // @[playground/src/noop/crossbar.scala 40:18 playground/src/axi/axi.scala 58:23]
  wire  _GEN_279 = 4'h2 == state ? 1'h0 : _GEN_227; // @[playground/src/axi/axi.scala 102:18 playground/src/noop/crossbar.scala 40:18]
  wire  _GEN_280 = 4'h2 == state ? 1'h0 : _GEN_228; // @[playground/src/axi/axi.scala 101:18 playground/src/noop/crossbar.scala 40:18]
  wire  _GEN_281 = 4'h2 == state ? 1'h0 : _GEN_229; // @[playground/src/axi/axi.scala 105:18 playground/src/noop/crossbar.scala 40:18]
  wire [3:0] _GEN_282 = 4'h2 == state ? 4'h0 : _GEN_230; // @[playground/src/noop/crossbar.scala 40:18 playground/src/axi/axi.scala 68:23]
  wire [63:0] _GEN_283 = 4'h2 == state ? 64'h0 : _GEN_231; // @[playground/src/noop/crossbar.scala 40:18 playground/src/axi/axi.scala 68:23]
  wire [1:0] _GEN_284 = 4'h2 == state ? 2'h0 : _GEN_232; // @[playground/src/noop/crossbar.scala 40:18 playground/src/axi/axi.scala 68:23]
  wire  _GEN_285 = 4'h2 == state ? 1'h0 : _GEN_233; // @[playground/src/noop/crossbar.scala 40:18 playground/src/axi/axi.scala 68:23]
  wire  _GEN_286 = 4'h2 == state ? 1'h0 : _GEN_234; // @[playground/src/axi/axi.scala 104:18 playground/src/noop/crossbar.scala 40:18]
  wire  _GEN_287 = 4'h2 == state ? 1'h0 : _GEN_235; // @[playground/src/axi/axi.scala 103:18 playground/src/noop/crossbar.scala 40:18]
  wire [3:0] _GEN_288 = 4'h2 == state ? 4'h0 : _GEN_236; // @[playground/src/noop/crossbar.scala 40:18 playground/src/axi/axi.scala 58:23]
  wire [1:0] _GEN_289 = 4'h2 == state ? 2'h0 : _GEN_237; // @[playground/src/noop/crossbar.scala 40:18 playground/src/axi/axi.scala 58:23]
  wire  _GEN_290 = 4'h2 == state ? 1'h0 : _GEN_238; // @[playground/src/axi/axi.scala 102:18 playground/src/noop/crossbar.scala 40:18]
  wire  _GEN_291 = 4'h2 == state ? 1'h0 : _GEN_239; // @[playground/src/axi/axi.scala 101:18 playground/src/noop/crossbar.scala 40:18]
  wire  _GEN_292 = 4'h3 == state | _GEN_240; // @[playground/src/noop/crossbar.scala 40:18 67:23]
  wire  _GEN_293 = 4'h3 == state & io_outAxi_rd_valid; // @[playground/src/axi/axi.scala 105:18 playground/src/noop/crossbar.scala 40:18 67:23]
  wire [63:0] _GEN_295 = 4'h3 == state ? io_outAxi_rd_bits_data : 64'h0; // @[playground/src/noop/crossbar.scala 40:18 67:23 playground/src/axi/axi.scala 68:23]
  wire  _GEN_297 = 4'h3 == state & io_outAxi_rd_bits_last; // @[playground/src/noop/crossbar.scala 40:18 67:23 playground/src/axi/axi.scala 68:23]
  wire  _GEN_298 = 4'h3 == state & io_outAxi_ra_ready; // @[playground/src/axi/axi.scala 104:18 playground/src/noop/crossbar.scala 40:18 67:23]
  wire  _GEN_299 = 4'h3 == state ? io_memAxi_ra_valid : _GEN_247; // @[playground/src/noop/crossbar.scala 40:18 67:23]
  wire [3:0] _GEN_300 = 4'h3 == state ? 4'h0 : _GEN_248; // @[playground/src/noop/crossbar.scala 40:18 67:23]
  wire [31:0] _GEN_301 = 4'h3 == state ? io_memAxi_ra_bits_addr : _GEN_249; // @[playground/src/noop/crossbar.scala 40:18 67:23]
  wire [7:0] _GEN_302 = 4'h3 == state ? 8'h7 : _GEN_250; // @[playground/src/noop/crossbar.scala 40:18 67:23]
  wire [2:0] _GEN_303 = 4'h3 == state ? 3'h3 : _GEN_251; // @[playground/src/noop/crossbar.scala 40:18 67:23]
  wire [1:0] _GEN_304 = 4'h3 == state ? 2'h1 : _GEN_252; // @[playground/src/noop/crossbar.scala 40:18 67:23]
  wire  _GEN_305 = 4'h3 == state | _GEN_253; // @[playground/src/noop/crossbar.scala 40:18 67:23]
  wire  _GEN_309 = 4'h3 == state & io_outAxi_wd_ready; // @[playground/src/axi/axi.scala 102:18 playground/src/noop/crossbar.scala 40:18 67:23]
  wire  _GEN_310 = 4'h3 == state ? io_memAxi_wd_valid : _GEN_258; // @[playground/src/noop/crossbar.scala 40:18 67:23]
  wire [63:0] _GEN_311 = 4'h3 == state ? io_memAxi_wd_bits_data : _GEN_259; // @[playground/src/noop/crossbar.scala 40:18 67:23]
  wire [7:0] _GEN_312 = 4'h3 == state ? 8'hff : _GEN_260; // @[playground/src/noop/crossbar.scala 40:18 67:23]
  wire  _GEN_313 = 4'h3 == state ? io_memAxi_wd_bits_last : _GEN_261; // @[playground/src/noop/crossbar.scala 40:18 67:23]
  wire  _GEN_314 = 4'h3 == state & io_outAxi_wa_ready; // @[playground/src/axi/axi.scala 101:18 playground/src/noop/crossbar.scala 40:18 67:23]
  wire  _GEN_315 = 4'h3 == state ? io_memAxi_wa_valid : _GEN_263; // @[playground/src/noop/crossbar.scala 40:18 67:23]
  wire [3:0] _GEN_316 = 4'h3 == state ? 4'h0 : _GEN_264; // @[playground/src/noop/crossbar.scala 40:18 67:23]
  wire [31:0] _GEN_317 = 4'h3 == state ? io_memAxi_wa_bits_addr : _GEN_265; // @[playground/src/noop/crossbar.scala 40:18 67:23]
  wire [7:0] _GEN_318 = 4'h3 == state ? 8'h7 : _GEN_266; // @[playground/src/noop/crossbar.scala 40:18 67:23]
  wire [2:0] _GEN_319 = 4'h3 == state ? 3'h3 : _GEN_267; // @[playground/src/noop/crossbar.scala 40:18 67:23]
  wire [1:0] _GEN_320 = 4'h3 == state ? 2'h1 : _GEN_268; // @[playground/src/noop/crossbar.scala 40:18 67:23]
  wire  _GEN_323 = 4'h3 == state ? 1'h0 : _GEN_241; // @[playground/src/axi/axi.scala 105:18 playground/src/noop/crossbar.scala 40:18]
  wire [63:0] _GEN_325 = 4'h3 == state ? 64'h0 : _GEN_243; // @[playground/src/noop/crossbar.scala 40:18 playground/src/axi/axi.scala 68:23]
  wire  _GEN_327 = 4'h3 == state ? 1'h0 : _GEN_245; // @[playground/src/noop/crossbar.scala 40:18 playground/src/axi/axi.scala 68:23]
  wire  _GEN_328 = 4'h3 == state ? 1'h0 : _GEN_246; // @[playground/src/axi/axi.scala 104:18 playground/src/noop/crossbar.scala 40:18]
  wire  _GEN_334 = 4'h3 == state ? 1'h0 : _GEN_270; // @[playground/src/axi/axi.scala 105:18 playground/src/noop/crossbar.scala 40:18]
  wire [3:0] _GEN_335 = 4'h3 == state ? 4'h0 : _GEN_271; // @[playground/src/noop/crossbar.scala 40:18 playground/src/axi/axi.scala 68:23]
  wire [63:0] _GEN_336 = 4'h3 == state ? 64'h0 : _GEN_272; // @[playground/src/noop/crossbar.scala 40:18 playground/src/axi/axi.scala 68:23]
  wire [1:0] _GEN_337 = 4'h3 == state ? 2'h0 : _GEN_273; // @[playground/src/noop/crossbar.scala 40:18 playground/src/axi/axi.scala 68:23]
  wire  _GEN_338 = 4'h3 == state ? 1'h0 : _GEN_274; // @[playground/src/noop/crossbar.scala 40:18 playground/src/axi/axi.scala 68:23]
  wire  _GEN_339 = 4'h3 == state ? 1'h0 : _GEN_275; // @[playground/src/axi/axi.scala 104:18 playground/src/noop/crossbar.scala 40:18]
  wire  _GEN_340 = 4'h3 == state ? 1'h0 : _GEN_276; // @[playground/src/axi/axi.scala 103:18 playground/src/noop/crossbar.scala 40:18]
  wire [3:0] _GEN_341 = 4'h3 == state ? 4'h0 : _GEN_277; // @[playground/src/noop/crossbar.scala 40:18 playground/src/axi/axi.scala 58:23]
  wire [1:0] _GEN_342 = 4'h3 == state ? 2'h0 : _GEN_278; // @[playground/src/noop/crossbar.scala 40:18 playground/src/axi/axi.scala 58:23]
  wire  _GEN_343 = 4'h3 == state ? 1'h0 : _GEN_279; // @[playground/src/axi/axi.scala 102:18 playground/src/noop/crossbar.scala 40:18]
  wire  _GEN_344 = 4'h3 == state ? 1'h0 : _GEN_280; // @[playground/src/axi/axi.scala 101:18 playground/src/noop/crossbar.scala 40:18]
  wire  _GEN_345 = 4'h3 == state ? 1'h0 : _GEN_281; // @[playground/src/axi/axi.scala 105:18 playground/src/noop/crossbar.scala 40:18]
  wire [3:0] _GEN_346 = 4'h3 == state ? 4'h0 : _GEN_282; // @[playground/src/noop/crossbar.scala 40:18 playground/src/axi/axi.scala 68:23]
  wire [63:0] _GEN_347 = 4'h3 == state ? 64'h0 : _GEN_283; // @[playground/src/noop/crossbar.scala 40:18 playground/src/axi/axi.scala 68:23]
  wire [1:0] _GEN_348 = 4'h3 == state ? 2'h0 : _GEN_284; // @[playground/src/noop/crossbar.scala 40:18 playground/src/axi/axi.scala 68:23]
  wire  _GEN_349 = 4'h3 == state ? 1'h0 : _GEN_285; // @[playground/src/noop/crossbar.scala 40:18 playground/src/axi/axi.scala 68:23]
  wire  _GEN_350 = 4'h3 == state ? 1'h0 : _GEN_286; // @[playground/src/axi/axi.scala 104:18 playground/src/noop/crossbar.scala 40:18]
  wire  _GEN_351 = 4'h3 == state ? 1'h0 : _GEN_287; // @[playground/src/axi/axi.scala 103:18 playground/src/noop/crossbar.scala 40:18]
  wire [3:0] _GEN_352 = 4'h3 == state ? 4'h0 : _GEN_288; // @[playground/src/noop/crossbar.scala 40:18 playground/src/axi/axi.scala 58:23]
  wire [1:0] _GEN_353 = 4'h3 == state ? 2'h0 : _GEN_289; // @[playground/src/noop/crossbar.scala 40:18 playground/src/axi/axi.scala 58:23]
  wire  _GEN_354 = 4'h3 == state ? 1'h0 : _GEN_290; // @[playground/src/axi/axi.scala 102:18 playground/src/noop/crossbar.scala 40:18]
  wire  _GEN_355 = 4'h3 == state ? 1'h0 : _GEN_291; // @[playground/src/axi/axi.scala 101:18 playground/src/noop/crossbar.scala 40:18]
  wire  _GEN_358 = 4'h1 == state ? _GEN_9 : _GEN_292; // @[playground/src/noop/crossbar.scala 40:18]
  wire  _GEN_359 = 4'h1 == state ? _GEN_10 : _GEN_293; // @[playground/src/noop/crossbar.scala 40:18]
  wire [63:0] _GEN_361 = 4'h1 == state ? _GEN_12 : _GEN_295; // @[playground/src/noop/crossbar.scala 40:18]
  wire  _GEN_363 = 4'h1 == state ? _GEN_14 : _GEN_297; // @[playground/src/noop/crossbar.scala 40:18]
  wire  _GEN_364 = 4'h1 == state ? _GEN_15 : _GEN_298; // @[playground/src/noop/crossbar.scala 40:18]
  wire  _GEN_365 = 4'h1 == state ? _GEN_16 : _GEN_299; // @[playground/src/noop/crossbar.scala 40:18]
  wire [3:0] _GEN_366 = 4'h1 == state ? 4'h0 : _GEN_300; // @[playground/src/noop/crossbar.scala 40:18]
  wire [31:0] _GEN_367 = 4'h1 == state ? _GEN_18 : _GEN_301; // @[playground/src/noop/crossbar.scala 40:18]
  wire [7:0] _GEN_368 = 4'h1 == state ? _GEN_19 : _GEN_302; // @[playground/src/noop/crossbar.scala 40:18]
  wire [2:0] _GEN_369 = 4'h1 == state ? _GEN_20 : _GEN_303; // @[playground/src/noop/crossbar.scala 40:18]
  wire [1:0] _GEN_370 = 4'h1 == state ? _GEN_21 : _GEN_304; // @[playground/src/noop/crossbar.scala 40:18]
  wire  _GEN_375 = 4'h1 == state ? _GEN_26 : _GEN_309; // @[playground/src/noop/crossbar.scala 40:18]
  wire  _GEN_376 = 4'h1 == state ? _GEN_27 : _GEN_310; // @[playground/src/noop/crossbar.scala 40:18]
  wire [63:0] _GEN_377 = 4'h1 == state ? _GEN_28 : _GEN_311; // @[playground/src/noop/crossbar.scala 40:18]
  wire [7:0] _GEN_378 = 4'h1 == state ? _GEN_29 : _GEN_312; // @[playground/src/noop/crossbar.scala 40:18]
  wire  _GEN_379 = 4'h1 == state ? _GEN_30 : _GEN_313; // @[playground/src/noop/crossbar.scala 40:18]
  wire  _GEN_380 = 4'h1 == state ? _GEN_31 : _GEN_314; // @[playground/src/noop/crossbar.scala 40:18]
  wire  _GEN_381 = 4'h1 == state ? _GEN_32 : _GEN_315; // @[playground/src/noop/crossbar.scala 40:18]
  wire [3:0] _GEN_382 = 4'h1 == state ? 4'h0 : _GEN_316; // @[playground/src/noop/crossbar.scala 40:18]
  wire [31:0] _GEN_383 = 4'h1 == state ? _GEN_34 : _GEN_317; // @[playground/src/noop/crossbar.scala 40:18]
  wire [7:0] _GEN_384 = 4'h1 == state ? _GEN_19 : _GEN_318; // @[playground/src/noop/crossbar.scala 40:18]
  wire [2:0] _GEN_385 = 4'h1 == state ? _GEN_20 : _GEN_319; // @[playground/src/noop/crossbar.scala 40:18]
  wire [1:0] _GEN_386 = 4'h1 == state ? _GEN_21 : _GEN_320; // @[playground/src/noop/crossbar.scala 40:18]
  wire  _GEN_387 = 4'h1 == state ? 1'h0 : _GEN_323; // @[playground/src/axi/axi.scala 105:18 playground/src/noop/crossbar.scala 40:18]
  wire [63:0] _GEN_389 = 4'h1 == state ? 64'h0 : _GEN_325; // @[playground/src/noop/crossbar.scala 40:18 playground/src/axi/axi.scala 68:23]
  wire  _GEN_391 = 4'h1 == state ? 1'h0 : _GEN_327; // @[playground/src/noop/crossbar.scala 40:18 playground/src/axi/axi.scala 68:23]
  wire  _GEN_392 = 4'h1 == state ? 1'h0 : _GEN_328; // @[playground/src/axi/axi.scala 104:18 playground/src/noop/crossbar.scala 40:18]
  wire  _GEN_398 = 4'h1 == state ? 1'h0 : _GEN_334; // @[playground/src/axi/axi.scala 105:18 playground/src/noop/crossbar.scala 40:18]
  wire [3:0] _GEN_399 = 4'h1 == state ? 4'h0 : _GEN_335; // @[playground/src/noop/crossbar.scala 40:18 playground/src/axi/axi.scala 68:23]
  wire [63:0] _GEN_400 = 4'h1 == state ? 64'h0 : _GEN_336; // @[playground/src/noop/crossbar.scala 40:18 playground/src/axi/axi.scala 68:23]
  wire [1:0] _GEN_401 = 4'h1 == state ? 2'h0 : _GEN_337; // @[playground/src/noop/crossbar.scala 40:18 playground/src/axi/axi.scala 68:23]
  wire  _GEN_402 = 4'h1 == state ? 1'h0 : _GEN_338; // @[playground/src/noop/crossbar.scala 40:18 playground/src/axi/axi.scala 68:23]
  wire  _GEN_403 = 4'h1 == state ? 1'h0 : _GEN_339; // @[playground/src/axi/axi.scala 104:18 playground/src/noop/crossbar.scala 40:18]
  wire  _GEN_404 = 4'h1 == state ? 1'h0 : _GEN_340; // @[playground/src/axi/axi.scala 103:18 playground/src/noop/crossbar.scala 40:18]
  wire [3:0] _GEN_405 = 4'h1 == state ? 4'h0 : _GEN_341; // @[playground/src/noop/crossbar.scala 40:18 playground/src/axi/axi.scala 58:23]
  wire [1:0] _GEN_406 = 4'h1 == state ? 2'h0 : _GEN_342; // @[playground/src/noop/crossbar.scala 40:18 playground/src/axi/axi.scala 58:23]
  wire  _GEN_407 = 4'h1 == state ? 1'h0 : _GEN_343; // @[playground/src/axi/axi.scala 102:18 playground/src/noop/crossbar.scala 40:18]
  wire  _GEN_408 = 4'h1 == state ? 1'h0 : _GEN_344; // @[playground/src/axi/axi.scala 101:18 playground/src/noop/crossbar.scala 40:18]
  wire  _GEN_409 = 4'h1 == state ? 1'h0 : _GEN_345; // @[playground/src/axi/axi.scala 105:18 playground/src/noop/crossbar.scala 40:18]
  wire [3:0] _GEN_410 = 4'h1 == state ? 4'h0 : _GEN_346; // @[playground/src/noop/crossbar.scala 40:18 playground/src/axi/axi.scala 68:23]
  wire [63:0] _GEN_411 = 4'h1 == state ? 64'h0 : _GEN_347; // @[playground/src/noop/crossbar.scala 40:18 playground/src/axi/axi.scala 68:23]
  wire [1:0] _GEN_412 = 4'h1 == state ? 2'h0 : _GEN_348; // @[playground/src/noop/crossbar.scala 40:18 playground/src/axi/axi.scala 68:23]
  wire  _GEN_413 = 4'h1 == state ? 1'h0 : _GEN_349; // @[playground/src/noop/crossbar.scala 40:18 playground/src/axi/axi.scala 68:23]
  wire  _GEN_414 = 4'h1 == state ? 1'h0 : _GEN_350; // @[playground/src/axi/axi.scala 104:18 playground/src/noop/crossbar.scala 40:18]
  wire  _GEN_415 = 4'h1 == state ? 1'h0 : _GEN_351; // @[playground/src/axi/axi.scala 103:18 playground/src/noop/crossbar.scala 40:18]
  wire [3:0] _GEN_416 = 4'h1 == state ? 4'h0 : _GEN_352; // @[playground/src/noop/crossbar.scala 40:18 playground/src/axi/axi.scala 58:23]
  wire [1:0] _GEN_417 = 4'h1 == state ? 2'h0 : _GEN_353; // @[playground/src/noop/crossbar.scala 40:18 playground/src/axi/axi.scala 58:23]
  wire  _GEN_418 = 4'h1 == state ? 1'h0 : _GEN_354; // @[playground/src/axi/axi.scala 102:18 playground/src/noop/crossbar.scala 40:18]
  wire  _GEN_419 = 4'h1 == state ? 1'h0 : _GEN_355; // @[playground/src/axi/axi.scala 101:18 playground/src/noop/crossbar.scala 40:18]
  assign io_icAxi_ra_ready = 4'h0 == state ? 1'h0 : _GEN_392; // @[playground/src/axi/axi.scala 104:18 playground/src/noop/crossbar.scala 40:18]
  assign io_icAxi_rd_valid = 4'h0 == state ? 1'h0 : _GEN_387; // @[playground/src/axi/axi.scala 105:18 playground/src/noop/crossbar.scala 40:18]
  assign io_icAxi_rd_bits_data = 4'h0 == state ? 64'h0 : _GEN_389; // @[playground/src/noop/crossbar.scala 40:18 playground/src/axi/axi.scala 68:23]
  assign io_icAxi_rd_bits_last = 4'h0 == state ? 1'h0 : _GEN_391; // @[playground/src/noop/crossbar.scala 40:18 playground/src/axi/axi.scala 68:23]
  assign io_flashAxi_wa_ready = 4'h0 == state ? 1'h0 : _GEN_408; // @[playground/src/axi/axi.scala 101:18 playground/src/noop/crossbar.scala 40:18]
  assign io_flashAxi_wd_ready = 4'h0 == state ? 1'h0 : _GEN_407; // @[playground/src/axi/axi.scala 102:18 playground/src/noop/crossbar.scala 40:18]
  assign io_flashAxi_wr_valid = 4'h0 == state ? 1'h0 : _GEN_404; // @[playground/src/axi/axi.scala 103:18 playground/src/noop/crossbar.scala 40:18]
  assign io_flashAxi_wr_bits_id = 4'h0 == state ? 4'h0 : _GEN_405; // @[playground/src/noop/crossbar.scala 40:18 playground/src/axi/axi.scala 58:23]
  assign io_flashAxi_wr_bits_resp = 4'h0 == state ? 2'h0 : _GEN_406; // @[playground/src/noop/crossbar.scala 40:18 playground/src/axi/axi.scala 58:23]
  assign io_flashAxi_ra_ready = 4'h0 == state ? 1'h0 : _GEN_403; // @[playground/src/axi/axi.scala 104:18 playground/src/noop/crossbar.scala 40:18]
  assign io_flashAxi_rd_valid = 4'h0 == state ? 1'h0 : _GEN_398; // @[playground/src/axi/axi.scala 105:18 playground/src/noop/crossbar.scala 40:18]
  assign io_flashAxi_rd_bits_id = 4'h0 == state ? 4'h0 : _GEN_399; // @[playground/src/noop/crossbar.scala 40:18 playground/src/axi/axi.scala 68:23]
  assign io_flashAxi_rd_bits_data = 4'h0 == state ? 64'h0 : _GEN_400; // @[playground/src/noop/crossbar.scala 40:18 playground/src/axi/axi.scala 68:23]
  assign io_flashAxi_rd_bits_resp = 4'h0 == state ? 2'h0 : _GEN_401; // @[playground/src/noop/crossbar.scala 40:18 playground/src/axi/axi.scala 68:23]
  assign io_flashAxi_rd_bits_last = 4'h0 == state ? 1'h0 : _GEN_402; // @[playground/src/noop/crossbar.scala 40:18 playground/src/axi/axi.scala 68:23]
  assign io_memAxi_wa_ready = 4'h0 == state ? 1'h0 : _GEN_380; // @[playground/src/axi/axi.scala 101:18 playground/src/noop/crossbar.scala 40:18]
  assign io_memAxi_wd_ready = 4'h0 == state ? 1'h0 : _GEN_375; // @[playground/src/axi/axi.scala 102:18 playground/src/noop/crossbar.scala 40:18]
  assign io_memAxi_ra_ready = 4'h0 == state ? 1'h0 : _GEN_364; // @[playground/src/axi/axi.scala 104:18 playground/src/noop/crossbar.scala 40:18]
  assign io_memAxi_rd_valid = 4'h0 == state ? 1'h0 : _GEN_359; // @[playground/src/axi/axi.scala 105:18 playground/src/noop/crossbar.scala 40:18]
  assign io_memAxi_rd_bits_data = 4'h0 == state ? 64'h0 : _GEN_361; // @[playground/src/noop/crossbar.scala 40:18 playground/src/axi/axi.scala 68:23]
  assign io_memAxi_rd_bits_last = 4'h0 == state ? 1'h0 : _GEN_363; // @[playground/src/noop/crossbar.scala 40:18 playground/src/axi/axi.scala 68:23]
  assign io_mmioAxi_wa_ready = 4'h0 == state ? 1'h0 : _GEN_419; // @[playground/src/axi/axi.scala 101:18 playground/src/noop/crossbar.scala 40:18]
  assign io_mmioAxi_wd_ready = 4'h0 == state ? 1'h0 : _GEN_418; // @[playground/src/axi/axi.scala 102:18 playground/src/noop/crossbar.scala 40:18]
  assign io_mmioAxi_wr_valid = 4'h0 == state ? 1'h0 : _GEN_415; // @[playground/src/axi/axi.scala 103:18 playground/src/noop/crossbar.scala 40:18]
  assign io_mmioAxi_wr_bits_id = 4'h0 == state ? 4'h0 : _GEN_416; // @[playground/src/noop/crossbar.scala 40:18 playground/src/axi/axi.scala 58:23]
  assign io_mmioAxi_wr_bits_resp = 4'h0 == state ? 2'h0 : _GEN_417; // @[playground/src/noop/crossbar.scala 40:18 playground/src/axi/axi.scala 58:23]
  assign io_mmioAxi_ra_ready = 4'h0 == state ? 1'h0 : _GEN_414; // @[playground/src/axi/axi.scala 104:18 playground/src/noop/crossbar.scala 40:18]
  assign io_mmioAxi_rd_valid = 4'h0 == state ? 1'h0 : _GEN_409; // @[playground/src/axi/axi.scala 105:18 playground/src/noop/crossbar.scala 40:18]
  assign io_mmioAxi_rd_bits_id = 4'h0 == state ? 4'h0 : _GEN_410; // @[playground/src/noop/crossbar.scala 40:18 playground/src/axi/axi.scala 68:23]
  assign io_mmioAxi_rd_bits_data = 4'h0 == state ? 64'h0 : _GEN_411; // @[playground/src/noop/crossbar.scala 40:18 playground/src/axi/axi.scala 68:23]
  assign io_mmioAxi_rd_bits_resp = 4'h0 == state ? 2'h0 : _GEN_412; // @[playground/src/noop/crossbar.scala 40:18 playground/src/axi/axi.scala 68:23]
  assign io_mmioAxi_rd_bits_last = 4'h0 == state ? 1'h0 : _GEN_413; // @[playground/src/noop/crossbar.scala 40:18 playground/src/axi/axi.scala 68:23]
  assign io_outAxi_wa_valid = 4'h0 == state ? 1'h0 : _GEN_381; // @[playground/src/noop/crossbar.scala 40:18 playground/src/axi/axi.scala 83:18]
  assign io_outAxi_wa_bits_id = 4'h0 == state ? 4'h0 : _GEN_382; // @[playground/src/noop/crossbar.scala 40:18 playground/src/axi/axi.scala 41:23]
  assign io_outAxi_wa_bits_addr = 4'h0 == state ? 32'h0 : _GEN_383; // @[playground/src/noop/crossbar.scala 40:18 playground/src/axi/axi.scala 41:23]
  assign io_outAxi_wa_bits_len = 4'h0 == state ? 8'h0 : _GEN_384; // @[playground/src/noop/crossbar.scala 40:18 playground/src/axi/axi.scala 41:23]
  assign io_outAxi_wa_bits_size = 4'h0 == state ? 3'h0 : _GEN_385; // @[playground/src/noop/crossbar.scala 40:18 playground/src/axi/axi.scala 41:23]
  assign io_outAxi_wa_bits_burst = 4'h0 == state ? 2'h0 : _GEN_386; // @[playground/src/noop/crossbar.scala 40:18 playground/src/axi/axi.scala 41:23]
  assign io_outAxi_wd_valid = 4'h0 == state ? 1'h0 : _GEN_376; // @[playground/src/noop/crossbar.scala 40:18 playground/src/axi/axi.scala 84:18]
  assign io_outAxi_wd_bits_data = 4'h0 == state ? 64'h0 : _GEN_377; // @[playground/src/noop/crossbar.scala 40:18 playground/src/axi/axi.scala 50:23]
  assign io_outAxi_wd_bits_strb = 4'h0 == state ? 8'h0 : _GEN_378; // @[playground/src/noop/crossbar.scala 40:18 playground/src/axi/axi.scala 50:23]
  assign io_outAxi_wd_bits_last = 4'h0 == state ? 1'h0 : _GEN_379; // @[playground/src/noop/crossbar.scala 40:18 playground/src/axi/axi.scala 50:23]
  assign io_outAxi_wr_ready = 4'h0 == state | (4'h1 == state | _GEN_305); // @[playground/src/noop/crossbar.scala 40:18 29:24]
  assign io_outAxi_ra_valid = 4'h0 == state ? 1'h0 : _GEN_365; // @[playground/src/noop/crossbar.scala 40:18 playground/src/axi/axi.scala 86:18]
  assign io_outAxi_ra_bits_id = 4'h0 == state ? 4'h0 : _GEN_366; // @[playground/src/noop/crossbar.scala 40:18 playground/src/axi/axi.scala 41:23]
  assign io_outAxi_ra_bits_addr = 4'h0 == state ? 32'h0 : _GEN_367; // @[playground/src/noop/crossbar.scala 40:18 playground/src/axi/axi.scala 41:23]
  assign io_outAxi_ra_bits_len = 4'h0 == state ? 8'h0 : _GEN_368; // @[playground/src/noop/crossbar.scala 40:18 playground/src/axi/axi.scala 41:23]
  assign io_outAxi_ra_bits_size = 4'h0 == state ? 3'h0 : _GEN_369; // @[playground/src/noop/crossbar.scala 40:18 playground/src/axi/axi.scala 41:23]
  assign io_outAxi_ra_bits_burst = 4'h0 == state ? 2'h0 : _GEN_370; // @[playground/src/noop/crossbar.scala 40:18 playground/src/axi/axi.scala 41:23]
  assign io_outAxi_rd_ready = 4'h0 == state ? 1'h0 : _GEN_358; // @[playground/src/noop/crossbar.scala 40:18 playground/src/axi/axi.scala 87:18]
  always @(posedge clock) begin
    if (reset) begin // @[playground/src/noop/crossbar.scala 20:24]
      state <= 4'h0; // @[playground/src/noop/crossbar.scala 20:24]
    end else if (4'h0 == state) begin // @[playground/src/noop/crossbar.scala 40:18]
      if (io_selectMem) begin // @[playground/src/noop/crossbar.scala 42:31]
        state <= 4'h1; // @[playground/src/noop/crossbar.scala 43:23]
      end else if (io_memAxi_ra_valid | io_memAxi_wa_valid) begin // @[playground/src/noop/crossbar.scala 45:65]
        state <= 4'h1; // @[playground/src/noop/crossbar.scala 46:23]
      end else begin
        state <= _GEN_2;
      end
    end else if (4'h1 == state) begin // @[playground/src/noop/crossbar.scala 40:18]
      if (selectMem_r & ~io_selectMem) begin // @[playground/src/noop/crossbar.scala 56:47]
        state <= 4'h0; // @[playground/src/noop/crossbar.scala 57:23]
      end else begin
        state <= _GEN_6;
      end
    end else if (4'h3 == state) begin // @[playground/src/noop/crossbar.scala 40:18]
      state <= _GEN_38;
    end else begin
      state <= _GEN_269;
    end
    if (reset) begin // @[playground/src/noop/crossbar.scala 22:30]
      selectMem_r <= 1'h0; // @[playground/src/noop/crossbar.scala 22:30]
    end else if (4'h0 == state) begin // @[playground/src/noop/crossbar.scala 40:18]
      selectMem_r <= _GEN_5;
    end else if (4'h1 == state) begin // @[playground/src/noop/crossbar.scala 40:18]
      if (selectMem_r & ~io_selectMem) begin // @[playground/src/noop/crossbar.scala 56:47]
        selectMem_r <= 1'h0; // @[playground/src/noop/crossbar.scala 58:29]
      end
    end else if (4'h3 == state) begin // @[playground/src/noop/crossbar.scala 40:18]
      selectMem_r <= _GEN_39;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[3:0];
  _RAND_1 = {1{`RANDOM}};
  selectMem_r = _RAND_1[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module FetchCrossBar(
  input         clock,
  input         reset,
  input  [31:0] io_instIO_addr, // @[playground/src/noop/fetch.scala 13:16]
  output [63:0] io_instIO_inst, // @[playground/src/noop/fetch.scala 13:16]
  input         io_instIO_arvalid, // @[playground/src/noop/fetch.scala 13:16]
  output        io_instIO_rvalid, // @[playground/src/noop/fetch.scala 13:16]
  output [31:0] io_icRead_addr, // @[playground/src/noop/fetch.scala 13:16]
  input  [63:0] io_icRead_inst, // @[playground/src/noop/fetch.scala 13:16]
  output        io_icRead_arvalid, // @[playground/src/noop/fetch.scala 13:16]
  input         io_icRead_rvalid, // @[playground/src/noop/fetch.scala 13:16]
  output [31:0] io_flashRead_addr, // @[playground/src/noop/fetch.scala 13:16]
  input  [63:0] io_flashRead_rdata, // @[playground/src/noop/fetch.scala 13:16]
  input         io_flashRead_rvalid, // @[playground/src/noop/fetch.scala 13:16]
  output [4:0]  io_flashRead_dc_mode // @[playground/src/noop/fetch.scala 13:16]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  reg  pre_mem; // @[playground/src/noop/fetch.scala 18:26]
  wire  inp_mem = io_instIO_addr[31]; // @[playground/src/noop/fetch.scala 19:33]
  wire [4:0] _GEN_2 = inp_mem ? 5'h0 : 5'h7; // @[playground/src/noop/fetch.scala 28:22 22:26 32:34]
  assign io_instIO_inst = pre_mem ? io_icRead_inst : io_flashRead_rdata; // @[playground/src/noop/fetch.scala 38:18 39:25 42:25]
  assign io_instIO_rvalid = pre_mem ? io_icRead_rvalid : io_flashRead_rvalid; // @[playground/src/noop/fetch.scala 38:18 40:26 43:26]
  assign io_icRead_addr = io_instIO_addr; // @[playground/src/noop/fetch.scala 23:25]
  assign io_icRead_arvalid = io_instIO_arvalid & inp_mem; // @[playground/src/noop/fetch.scala 24:25 26:28]
  assign io_flashRead_addr = io_instIO_addr; // @[playground/src/noop/fetch.scala 20:25]
  assign io_flashRead_dc_mode = io_instIO_arvalid ? _GEN_2 : 5'h0; // @[playground/src/noop/fetch.scala 22:26 26:28]
  always @(posedge clock) begin
    if (reset) begin // @[playground/src/noop/fetch.scala 18:26]
      pre_mem <= 1'h0; // @[playground/src/noop/fetch.scala 18:26]
    end else if (io_instIO_arvalid) begin // @[playground/src/noop/fetch.scala 26:28]
      pre_mem <= inp_mem; // @[playground/src/noop/fetch.scala 27:17]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  pre_mem = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Splite64to32(
  input         clock,
  input         reset,
  input  [31:0] io_data_in_addr, // @[playground/src/axi/toaxi.scala 12:16]
  output [63:0] io_data_in_rdata, // @[playground/src/axi/toaxi.scala 12:16]
  output        io_data_in_rvalid, // @[playground/src/axi/toaxi.scala 12:16]
  input  [4:0]  io_data_in_dc_mode, // @[playground/src/axi/toaxi.scala 12:16]
  output [31:0] io_data_out_addr, // @[playground/src/axi/toaxi.scala 12:16]
  input  [63:0] io_data_out_rdata, // @[playground/src/axi/toaxi.scala 12:16]
  input         io_data_out_rvalid, // @[playground/src/axi/toaxi.scala 12:16]
  output [4:0]  io_data_out_dc_mode, // @[playground/src/axi/toaxi.scala 12:16]
  input         io_data_out_ready // @[playground/src/axi/toaxi.scala 12:16]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] data_buf; // @[playground/src/axi/toaxi.scala 16:27]
  reg [31:0] addr_r; // @[playground/src/axi/toaxi.scala 18:25]
  reg  is_64; // @[playground/src/axi/toaxi.scala 19:24]
  reg  busy; // @[playground/src/axi/toaxi.scala 20:23]
  reg  state; // @[playground/src/axi/toaxi.scala 21:24]
  wire  hs_out = io_data_out_dc_mode != 5'h0 & io_data_out_ready; // @[playground/src/axi/toaxi.scala 22:53]
  wire [63:0] _io_data_in_rdata_T_1 = {io_data_out_rdata[31:0],data_buf}; // @[playground/src/axi/toaxi.scala 25:39]
  wire [31:0] _io_data_out_addr_T_1 = {io_data_in_addr[31:3],3'h0}; // @[playground/src/axi/toaxi.scala 30:44]
  wire  _GEN_0 = hs_out ? 1'h0 : is_64; // @[playground/src/axi/toaxi.scala 19:24 37:39 38:31]
  wire  _GEN_1 = hs_out & io_data_out_dc_mode != 5'h7 | state; // @[playground/src/axi/toaxi.scala 21:24 33:68 34:31]
  wire  _GEN_3 = hs_out & io_data_out_dc_mode != 5'h7 | _GEN_0; // @[playground/src/axi/toaxi.scala 33:68 36:31]
  wire  _GEN_4 = io_data_in_rvalid ? 1'h0 : busy; // @[playground/src/axi/toaxi.scala 20:23 40:46 41:26]
  wire  _GEN_5 = io_data_in_dc_mode != 5'h0 | _GEN_4; // @[playground/src/axi/toaxi.scala 28:54 29:26]
  wire [31:0] _GEN_6 = io_data_in_dc_mode != 5'h0 ? _io_data_out_addr_T_1 : 32'h0; // @[playground/src/axi/toaxi.scala 23:108 28:54 30:38]
  wire [4:0] _GEN_7 = io_data_in_dc_mode != 5'h0 ? 5'h16 : 5'h0; // @[playground/src/axi/toaxi.scala 28:54 31:41 23:77]
  wire  _GEN_12 = busy & io_data_out_rvalid; // @[playground/src/axi/toaxi.scala 43:27 44:39 24:52]
  wire [63:0] _GEN_13 = io_data_out_rvalid ? io_data_out_rdata : {{32'd0}, data_buf}; // @[playground/src/axi/toaxi.scala 48:37 49:26 16:27]
  wire [31:0] _io_data_out_addr_T_3 = addr_r + 32'h4; // @[playground/src/axi/toaxi.scala 51:40]
  wire [63:0] _GEN_15 = state ? _GEN_13 : {{32'd0}, data_buf}; // @[playground/src/axi/toaxi.scala 26:18 16:27]
  wire [31:0] _GEN_16 = state ? _io_data_out_addr_T_3 : 32'h0; // @[playground/src/axi/toaxi.scala 23:108 26:18 51:30]
  wire [4:0] _GEN_17 = state ? 5'h16 : 5'h0; // @[playground/src/axi/toaxi.scala 26:18 52:33 23:77]
  wire [63:0] _GEN_27 = ~state ? {{32'd0}, data_buf} : _GEN_15; // @[playground/src/axi/toaxi.scala 26:18 16:27]
  wire [63:0] _GEN_8 = reset ? 64'h0 : _GEN_27; // @[playground/src/axi/toaxi.scala 16:{27,27}]
  assign io_data_in_rdata = is_64 ? _io_data_in_rdata_T_1 : io_data_out_rdata; // @[playground/src/axi/toaxi.scala 25:28]
  assign io_data_in_rvalid = ~state & _GEN_12; // @[playground/src/axi/toaxi.scala 26:18 24:52]
  assign io_data_out_addr = ~state ? _GEN_6 : _GEN_16; // @[playground/src/axi/toaxi.scala 26:18]
  assign io_data_out_dc_mode = ~state ? _GEN_7 : _GEN_17; // @[playground/src/axi/toaxi.scala 26:18]
  always @(posedge clock) begin
    data_buf <= _GEN_8[31:0]; // @[playground/src/axi/toaxi.scala 16:{27,27}]
    if (reset) begin // @[playground/src/axi/toaxi.scala 18:25]
      addr_r <= 32'h0; // @[playground/src/axi/toaxi.scala 18:25]
    end else if (~state) begin // @[playground/src/axi/toaxi.scala 26:18]
      if (io_data_in_dc_mode != 5'h0) begin // @[playground/src/axi/toaxi.scala 28:54]
        if (hs_out & io_data_out_dc_mode != 5'h7) begin // @[playground/src/axi/toaxi.scala 33:68]
          addr_r <= _io_data_out_addr_T_1; // @[playground/src/axi/toaxi.scala 35:32]
        end
      end
    end
    if (reset) begin // @[playground/src/axi/toaxi.scala 19:24]
      is_64 <= 1'h0; // @[playground/src/axi/toaxi.scala 19:24]
    end else if (~state) begin // @[playground/src/axi/toaxi.scala 26:18]
      if (io_data_in_dc_mode != 5'h0) begin // @[playground/src/axi/toaxi.scala 28:54]
        is_64 <= _GEN_3;
      end
    end
    if (reset) begin // @[playground/src/axi/toaxi.scala 20:23]
      busy <= 1'h0; // @[playground/src/axi/toaxi.scala 20:23]
    end else if (~state) begin // @[playground/src/axi/toaxi.scala 26:18]
      busy <= _GEN_5;
    end
    if (reset) begin // @[playground/src/axi/toaxi.scala 21:24]
      state <= 1'h0; // @[playground/src/axi/toaxi.scala 21:24]
    end else if (~state) begin // @[playground/src/axi/toaxi.scala 26:18]
      if (io_data_in_dc_mode != 5'h0) begin // @[playground/src/axi/toaxi.scala 28:54]
        state <= _GEN_1;
      end
    end else if (state) begin // @[playground/src/axi/toaxi.scala 26:18]
      if (hs_out) begin // @[playground/src/axi/toaxi.scala 53:25]
        state <= 1'h0; // @[playground/src/axi/toaxi.scala 54:23]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  data_buf = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  addr_r = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  is_64 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  busy = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  state = _RAND_4[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module MemCrossBar(
  input         clock,
  input         reset,
  input  [31:0] io_dataRW_addr, // @[playground/src/noop/memory.scala 16:16]
  output [63:0] io_dataRW_rdata, // @[playground/src/noop/memory.scala 16:16]
  output        io_dataRW_rvalid, // @[playground/src/noop/memory.scala 16:16]
  input  [63:0] io_dataRW_wdata, // @[playground/src/noop/memory.scala 16:16]
  input  [4:0]  io_dataRW_dc_mode, // @[playground/src/noop/memory.scala 16:16]
  input  [4:0]  io_dataRW_amo, // @[playground/src/noop/memory.scala 16:16]
  output        io_dataRW_ready, // @[playground/src/noop/memory.scala 16:16]
  output [31:0] io_mmio_addr, // @[playground/src/noop/memory.scala 16:16]
  input  [63:0] io_mmio_rdata, // @[playground/src/noop/memory.scala 16:16]
  input         io_mmio_rvalid, // @[playground/src/noop/memory.scala 16:16]
  output [63:0] io_mmio_wdata, // @[playground/src/noop/memory.scala 16:16]
  output [4:0]  io_mmio_dc_mode, // @[playground/src/noop/memory.scala 16:16]
  input         io_mmio_ready, // @[playground/src/noop/memory.scala 16:16]
  output [31:0] io_dcRW_addr, // @[playground/src/noop/memory.scala 16:16]
  input  [63:0] io_dcRW_rdata, // @[playground/src/noop/memory.scala 16:16]
  input         io_dcRW_rvalid, // @[playground/src/noop/memory.scala 16:16]
  output [63:0] io_dcRW_wdata, // @[playground/src/noop/memory.scala 16:16]
  output [4:0]  io_dcRW_dc_mode, // @[playground/src/noop/memory.scala 16:16]
  output [4:0]  io_dcRW_amo, // @[playground/src/noop/memory.scala 16:16]
  input         io_dcRW_ready, // @[playground/src/noop/memory.scala 16:16]
  output [31:0] io_clintIO_addr, // @[playground/src/noop/memory.scala 16:16]
  input  [63:0] io_clintIO_rdata, // @[playground/src/noop/memory.scala 16:16]
  output [63:0] io_clintIO_wdata, // @[playground/src/noop/memory.scala 16:16]
  output        io_clintIO_wvalid, // @[playground/src/noop/memory.scala 16:16]
  output [31:0] io_plicIO_addr, // @[playground/src/noop/memory.scala 16:16]
  input  [63:0] io_plicIO_rdata, // @[playground/src/noop/memory.scala 16:16]
  output [63:0] io_plicIO_wdata, // @[playground/src/noop/memory.scala 16:16]
  output        io_plicIO_wvalid, // @[playground/src/noop/memory.scala 16:16]
  output        io_plicIO_arvalid // @[playground/src/noop/memory.scala 16:16]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg [1:0] pre_type; // @[playground/src/noop/memory.scala 23:30]
  reg [63:0] data_r; // @[playground/src/noop/memory.scala 24:30]
  reg  data_valid; // @[playground/src/noop/memory.scala 25:30]
  wire  is_clint = io_dataRW_addr == 32'h200bff8 | io_dataRW_addr == 32'h2004000 | io_dataRW_addr == 32'h2000000; // @[playground/src/noop/memory.scala 27:79]
  wire  is_plic = io_dataRW_addr >= 32'hc000000 & io_dataRW_addr <= 32'hfffffff; // @[playground/src/noop/memory.scala 28:51]
  wire  inp_mem = io_dataRW_addr >= 32'h80000000 & io_dataRW_addr < 32'h90000000; // @[playground/src/noop/memory.scala 29:55]
  wire [4:0] _GEN_1 = inp_mem ? io_dataRW_dc_mode : 5'h0; // @[playground/src/noop/memory.scala 37:21 58:28 60:29]
  wire  _GEN_2 = inp_mem ? io_dcRW_ready : io_mmio_ready; // @[playground/src/noop/memory.scala 58:28 61:29 65:29]
  wire [4:0] _GEN_3 = inp_mem ? 5'h0 : io_dataRW_dc_mode; // @[playground/src/noop/memory.scala 38:21 58:28 64:29]
  wire  _GEN_5 = is_plic & io_dataRW_dc_mode[2]; // @[playground/src/noop/memory.scala 45:23 52:28 54:33]
  wire  _GEN_6 = is_plic & io_dataRW_dc_mode[3]; // @[playground/src/noop/memory.scala 44:23 52:28 55:33]
  wire  _GEN_8 = is_plic | data_valid; // @[playground/src/noop/memory.scala 52:28 25:30 57:33]
  wire [4:0] _GEN_9 = is_plic ? 5'h0 : _GEN_1; // @[playground/src/noop/memory.scala 37:21 52:28]
  wire  _GEN_10 = is_plic ? 1'h0 : _GEN_2; // @[playground/src/noop/memory.scala 42:21 52:28]
  wire [4:0] _GEN_11 = is_plic ? 5'h0 : _GEN_3; // @[playground/src/noop/memory.scala 38:21 52:28]
  wire  _GEN_13 = is_clint & io_dataRW_dc_mode[3]; // @[playground/src/noop/memory.scala 43:23 47:23 49:33]
  wire  _GEN_15 = is_clint | _GEN_8; // @[playground/src/noop/memory.scala 47:23 51:33]
  wire  _GEN_16 = is_clint ? 1'h0 : _GEN_5; // @[playground/src/noop/memory.scala 45:23 47:23]
  wire  _GEN_17 = is_clint ? 1'h0 : _GEN_6; // @[playground/src/noop/memory.scala 44:23 47:23]
  wire [4:0] _GEN_18 = is_clint ? 5'h0 : _GEN_9; // @[playground/src/noop/memory.scala 37:21 47:23]
  wire  _GEN_19 = is_clint ? 1'h0 : _GEN_10; // @[playground/src/noop/memory.scala 42:21 47:23]
  wire [4:0] _GEN_20 = is_clint ? 5'h0 : _GEN_11; // @[playground/src/noop/memory.scala 38:21 47:23]
  wire [63:0] _GEN_30 = pre_type == 2'h0 ? io_mmio_rdata : 64'h0; // @[playground/src/noop/memory.scala 75:33 76:29 79:29]
  wire  _GEN_31 = pre_type == 2'h0 & io_mmio_rvalid; // @[playground/src/noop/memory.scala 75:33 77:29 80:29]
  wire [63:0] _GEN_32 = pre_type == 2'h1 ? io_dcRW_rdata : _GEN_30; // @[playground/src/noop/memory.scala 72:33 73:29]
  wire  _GEN_33 = pre_type == 2'h1 ? io_dcRW_rvalid : _GEN_31; // @[playground/src/noop/memory.scala 72:33 74:29]
  assign io_dataRW_rdata = (pre_type == 2'h2 | pre_type == 2'h3) & data_valid ? data_r : _GEN_32; // @[playground/src/noop/memory.scala 68:63 69:29]
  assign io_dataRW_rvalid = (pre_type == 2'h2 | pre_type == 2'h3) & data_valid | _GEN_33; // @[playground/src/noop/memory.scala 68:63 70:29]
  assign io_dataRW_ready = io_dataRW_dc_mode != 5'h0 & _GEN_19; // @[playground/src/noop/memory.scala 42:21 46:41]
  assign io_mmio_addr = io_dataRW_addr; // @[playground/src/noop/memory.scala 30:21]
  assign io_mmio_wdata = io_dataRW_wdata; // @[playground/src/noop/memory.scala 31:21]
  assign io_mmio_dc_mode = io_dataRW_dc_mode != 5'h0 ? _GEN_20 : 5'h0; // @[playground/src/noop/memory.scala 38:21 46:41]
  assign io_dcRW_addr = io_dataRW_addr; // @[playground/src/noop/memory.scala 32:21]
  assign io_dcRW_wdata = io_dataRW_wdata; // @[playground/src/noop/memory.scala 33:21]
  assign io_dcRW_dc_mode = io_dataRW_dc_mode != 5'h0 ? _GEN_18 : 5'h0; // @[playground/src/noop/memory.scala 37:21 46:41]
  assign io_dcRW_amo = io_dataRW_amo; // @[playground/src/noop/memory.scala 34:21]
  assign io_clintIO_addr = io_dataRW_addr; // @[playground/src/noop/memory.scala 35:24]
  assign io_clintIO_wdata = io_dataRW_wdata; // @[playground/src/noop/memory.scala 36:24]
  assign io_clintIO_wvalid = io_dataRW_dc_mode != 5'h0 & _GEN_13; // @[playground/src/noop/memory.scala 43:23 46:41]
  assign io_plicIO_addr = io_dataRW_addr; // @[playground/src/noop/memory.scala 40:21]
  assign io_plicIO_wdata = io_dataRW_wdata; // @[playground/src/noop/memory.scala 41:21]
  assign io_plicIO_wvalid = io_dataRW_dc_mode != 5'h0 & _GEN_17; // @[playground/src/noop/memory.scala 44:23 46:41]
  assign io_plicIO_arvalid = io_dataRW_dc_mode != 5'h0 & _GEN_16; // @[playground/src/noop/memory.scala 45:23 46:41]
  always @(posedge clock) begin
    if (reset) begin // @[playground/src/noop/memory.scala 23:30]
      pre_type <= 2'h0; // @[playground/src/noop/memory.scala 23:30]
    end else if (io_dataRW_dc_mode != 5'h0) begin // @[playground/src/noop/memory.scala 46:41]
      if (is_clint) begin // @[playground/src/noop/memory.scala 47:23]
        pre_type <= 2'h2; // @[playground/src/noop/memory.scala 48:33]
      end else if (is_plic) begin // @[playground/src/noop/memory.scala 52:28]
        pre_type <= 2'h3; // @[playground/src/noop/memory.scala 53:33]
      end else begin
        pre_type <= {{1'd0}, inp_mem};
      end
    end
    if (reset) begin // @[playground/src/noop/memory.scala 24:30]
      data_r <= 64'h0; // @[playground/src/noop/memory.scala 24:30]
    end else if (io_dataRW_dc_mode != 5'h0) begin // @[playground/src/noop/memory.scala 46:41]
      if (is_clint) begin // @[playground/src/noop/memory.scala 47:23]
        data_r <= io_clintIO_rdata; // @[playground/src/noop/memory.scala 50:33]
      end else if (is_plic) begin // @[playground/src/noop/memory.scala 52:28]
        data_r <= io_plicIO_rdata; // @[playground/src/noop/memory.scala 56:33]
      end
    end
    if (reset) begin // @[playground/src/noop/memory.scala 25:30]
      data_valid <= 1'h0; // @[playground/src/noop/memory.scala 25:30]
    end else if ((pre_type == 2'h2 | pre_type == 2'h3) & data_valid) begin // @[playground/src/noop/memory.scala 68:63]
      data_valid <= 1'h0; // @[playground/src/noop/memory.scala 71:29]
    end else if (io_dataRW_dc_mode != 5'h0) begin // @[playground/src/noop/memory.scala 46:41]
      data_valid <= _GEN_15;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  pre_type = _RAND_0[1:0];
  _RAND_1 = {2{`RANDOM}};
  data_r = _RAND_1[63:0];
  _RAND_2 = {1{`RANDOM}};
  data_valid = _RAND_2[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module MaxPeriodFibonacciLFSR_2(
  input   clock,
  input   reset,
  output  io_out_0, // @[src/main/scala/chisel3/util/random/PRNG.scala 42:22]
  output  io_out_1, // @[src/main/scala/chisel3/util/random/PRNG.scala 42:22]
  output  io_out_2, // @[src/main/scala/chisel3/util/random/PRNG.scala 42:22]
  output  io_out_3 // @[src/main/scala/chisel3/util/random/PRNG.scala 42:22]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  reg  state_0; // @[src/main/scala/chisel3/util/random/PRNG.scala 55:49]
  reg  state_1; // @[src/main/scala/chisel3/util/random/PRNG.scala 55:49]
  reg  state_2; // @[src/main/scala/chisel3/util/random/PRNG.scala 55:49]
  reg  state_3; // @[src/main/scala/chisel3/util/random/PRNG.scala 55:49]
  wire  _T = state_3 ^ state_2; // @[src/main/scala/chisel3/util/random/LFSR.scala 15:41]
  assign io_out_0 = state_0; // @[src/main/scala/chisel3/util/random/PRNG.scala 78:10]
  assign io_out_1 = state_1; // @[src/main/scala/chisel3/util/random/PRNG.scala 78:10]
  assign io_out_2 = state_2; // @[src/main/scala/chisel3/util/random/PRNG.scala 78:10]
  assign io_out_3 = state_3; // @[src/main/scala/chisel3/util/random/PRNG.scala 78:10]
  always @(posedge clock) begin
    state_0 <= reset | _T; // @[src/main/scala/chisel3/util/random/PRNG.scala 55:{49,49}]
    if (reset) begin // @[src/main/scala/chisel3/util/random/PRNG.scala 55:49]
      state_1 <= 1'h0; // @[src/main/scala/chisel3/util/random/PRNG.scala 55:49]
    end else begin
      state_1 <= state_0;
    end
    if (reset) begin // @[src/main/scala/chisel3/util/random/PRNG.scala 55:49]
      state_2 <= 1'h0; // @[src/main/scala/chisel3/util/random/PRNG.scala 55:49]
    end else begin
      state_2 <= state_1;
    end
    if (reset) begin // @[src/main/scala/chisel3/util/random/PRNG.scala 55:49]
      state_3 <= 1'h0; // @[src/main/scala/chisel3/util/random/PRNG.scala 55:49]
    end else begin
      state_3 <= state_2;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state_0 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  state_1 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  state_2 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  state_3 = _RAND_3[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TLB(
  input         clock,
  input         reset,
  input  [63:0] io_va2pa_vaddr, // @[playground/src/noop/tlb.scala 33:16]
  input         io_va2pa_vvalid, // @[playground/src/noop/tlb.scala 33:16]
  output        io_va2pa_ready, // @[playground/src/noop/tlb.scala 33:16]
  output [31:0] io_va2pa_paddr, // @[playground/src/noop/tlb.scala 33:16]
  output        io_va2pa_pvalid, // @[playground/src/noop/tlb.scala 33:16]
  output [63:0] io_va2pa_tlb_excep_cause, // @[playground/src/noop/tlb.scala 33:16]
  output [63:0] io_va2pa_tlb_excep_tval, // @[playground/src/noop/tlb.scala 33:16]
  output        io_va2pa_tlb_excep_en, // @[playground/src/noop/tlb.scala 33:16]
  input  [1:0]  io_mmuState_priv, // @[playground/src/noop/tlb.scala 33:16]
  input  [63:0] io_mmuState_mstatus, // @[playground/src/noop/tlb.scala 33:16]
  input  [63:0] io_mmuState_satp, // @[playground/src/noop/tlb.scala 33:16]
  input         io_flush, // @[playground/src/noop/tlb.scala 33:16]
  output [31:0] io_dcacheRW_addr, // @[playground/src/noop/tlb.scala 33:16]
  input  [63:0] io_dcacheRW_rdata, // @[playground/src/noop/tlb.scala 33:16]
  input         io_dcacheRW_rvalid, // @[playground/src/noop/tlb.scala 33:16]
  output [63:0] io_dcacheRW_wdata, // @[playground/src/noop/tlb.scala 33:16]
  output [4:0]  io_dcacheRW_dc_mode, // @[playground/src/noop/tlb.scala 33:16]
  input         io_dcacheRW_ready // @[playground/src/noop/tlb.scala 33:16]
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [63:0] _RAND_12;
  reg [63:0] _RAND_13;
  reg [63:0] _RAND_14;
  reg [63:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [63:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [63:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [63:0] _RAND_102;
  reg [63:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
`endif // RANDOMIZE_REG_INIT
  wire  select_prng_clock; // @[src/main/scala/chisel3/util/random/PRNG.scala 91:22]
  wire  select_prng_reset; // @[src/main/scala/chisel3/util/random/PRNG.scala 91:22]
  wire  select_prng_io_out_0; // @[src/main/scala/chisel3/util/random/PRNG.scala 91:22]
  wire  select_prng_io_out_1; // @[src/main/scala/chisel3/util/random/PRNG.scala 91:22]
  wire  select_prng_io_out_2; // @[src/main/scala/chisel3/util/random/PRNG.scala 91:22]
  wire  select_prng_io_out_3; // @[src/main/scala/chisel3/util/random/PRNG.scala 91:22]
  reg [51:0] tag_0; // @[playground/src/noop/tlb.scala 39:26]
  reg [51:0] tag_1; // @[playground/src/noop/tlb.scala 39:26]
  reg [51:0] tag_2; // @[playground/src/noop/tlb.scala 39:26]
  reg [51:0] tag_3; // @[playground/src/noop/tlb.scala 39:26]
  reg [51:0] tag_4; // @[playground/src/noop/tlb.scala 39:26]
  reg [51:0] tag_5; // @[playground/src/noop/tlb.scala 39:26]
  reg [51:0] tag_6; // @[playground/src/noop/tlb.scala 39:26]
  reg [51:0] tag_7; // @[playground/src/noop/tlb.scala 39:26]
  reg [51:0] tag_8; // @[playground/src/noop/tlb.scala 39:26]
  reg [51:0] tag_9; // @[playground/src/noop/tlb.scala 39:26]
  reg [51:0] tag_10; // @[playground/src/noop/tlb.scala 39:26]
  reg [51:0] tag_11; // @[playground/src/noop/tlb.scala 39:26]
  reg [51:0] tag_12; // @[playground/src/noop/tlb.scala 39:26]
  reg [51:0] tag_13; // @[playground/src/noop/tlb.scala 39:26]
  reg [51:0] tag_14; // @[playground/src/noop/tlb.scala 39:26]
  reg [51:0] tag_15; // @[playground/src/noop/tlb.scala 39:26]
  reg [19:0] paddr_0; // @[playground/src/noop/tlb.scala 40:26]
  reg [19:0] paddr_1; // @[playground/src/noop/tlb.scala 40:26]
  reg [19:0] paddr_2; // @[playground/src/noop/tlb.scala 40:26]
  reg [19:0] paddr_3; // @[playground/src/noop/tlb.scala 40:26]
  reg [19:0] paddr_4; // @[playground/src/noop/tlb.scala 40:26]
  reg [19:0] paddr_5; // @[playground/src/noop/tlb.scala 40:26]
  reg [19:0] paddr_6; // @[playground/src/noop/tlb.scala 40:26]
  reg [19:0] paddr_7; // @[playground/src/noop/tlb.scala 40:26]
  reg [19:0] paddr_8; // @[playground/src/noop/tlb.scala 40:26]
  reg [19:0] paddr_9; // @[playground/src/noop/tlb.scala 40:26]
  reg [19:0] paddr_10; // @[playground/src/noop/tlb.scala 40:26]
  reg [19:0] paddr_11; // @[playground/src/noop/tlb.scala 40:26]
  reg [19:0] paddr_12; // @[playground/src/noop/tlb.scala 40:26]
  reg [19:0] paddr_13; // @[playground/src/noop/tlb.scala 40:26]
  reg [19:0] paddr_14; // @[playground/src/noop/tlb.scala 40:26]
  reg [19:0] paddr_15; // @[playground/src/noop/tlb.scala 40:26]
  reg [9:0] info_0; // @[playground/src/noop/tlb.scala 41:26]
  reg [9:0] info_1; // @[playground/src/noop/tlb.scala 41:26]
  reg [9:0] info_2; // @[playground/src/noop/tlb.scala 41:26]
  reg [9:0] info_3; // @[playground/src/noop/tlb.scala 41:26]
  reg [9:0] info_4; // @[playground/src/noop/tlb.scala 41:26]
  reg [9:0] info_5; // @[playground/src/noop/tlb.scala 41:26]
  reg [9:0] info_6; // @[playground/src/noop/tlb.scala 41:26]
  reg [9:0] info_7; // @[playground/src/noop/tlb.scala 41:26]
  reg [9:0] info_8; // @[playground/src/noop/tlb.scala 41:26]
  reg [9:0] info_9; // @[playground/src/noop/tlb.scala 41:26]
  reg [9:0] info_10; // @[playground/src/noop/tlb.scala 41:26]
  reg [9:0] info_11; // @[playground/src/noop/tlb.scala 41:26]
  reg [9:0] info_12; // @[playground/src/noop/tlb.scala 41:26]
  reg [9:0] info_13; // @[playground/src/noop/tlb.scala 41:26]
  reg [9:0] info_14; // @[playground/src/noop/tlb.scala 41:26]
  reg [9:0] info_15; // @[playground/src/noop/tlb.scala 41:26]
  reg [31:0] pte_addr_0; // @[playground/src/noop/tlb.scala 42:30]
  reg [31:0] pte_addr_1; // @[playground/src/noop/tlb.scala 42:30]
  reg [31:0] pte_addr_2; // @[playground/src/noop/tlb.scala 42:30]
  reg [31:0] pte_addr_3; // @[playground/src/noop/tlb.scala 42:30]
  reg [31:0] pte_addr_4; // @[playground/src/noop/tlb.scala 42:30]
  reg [31:0] pte_addr_5; // @[playground/src/noop/tlb.scala 42:30]
  reg [31:0] pte_addr_6; // @[playground/src/noop/tlb.scala 42:30]
  reg [31:0] pte_addr_7; // @[playground/src/noop/tlb.scala 42:30]
  reg [31:0] pte_addr_8; // @[playground/src/noop/tlb.scala 42:30]
  reg [31:0] pte_addr_9; // @[playground/src/noop/tlb.scala 42:30]
  reg [31:0] pte_addr_10; // @[playground/src/noop/tlb.scala 42:30]
  reg [31:0] pte_addr_11; // @[playground/src/noop/tlb.scala 42:30]
  reg [31:0] pte_addr_12; // @[playground/src/noop/tlb.scala 42:30]
  reg [31:0] pte_addr_13; // @[playground/src/noop/tlb.scala 42:30]
  reg [31:0] pte_addr_14; // @[playground/src/noop/tlb.scala 42:30]
  reg [31:0] pte_addr_15; // @[playground/src/noop/tlb.scala 42:30]
  reg [1:0] pte_level_0; // @[playground/src/noop/tlb.scala 43:30]
  reg [1:0] pte_level_1; // @[playground/src/noop/tlb.scala 43:30]
  reg [1:0] pte_level_2; // @[playground/src/noop/tlb.scala 43:30]
  reg [1:0] pte_level_3; // @[playground/src/noop/tlb.scala 43:30]
  reg [1:0] pte_level_4; // @[playground/src/noop/tlb.scala 43:30]
  reg [1:0] pte_level_5; // @[playground/src/noop/tlb.scala 43:30]
  reg [1:0] pte_level_6; // @[playground/src/noop/tlb.scala 43:30]
  reg [1:0] pte_level_7; // @[playground/src/noop/tlb.scala 43:30]
  reg [1:0] pte_level_8; // @[playground/src/noop/tlb.scala 43:30]
  reg [1:0] pte_level_9; // @[playground/src/noop/tlb.scala 43:30]
  reg [1:0] pte_level_10; // @[playground/src/noop/tlb.scala 43:30]
  reg [1:0] pte_level_11; // @[playground/src/noop/tlb.scala 43:30]
  reg [1:0] pte_level_12; // @[playground/src/noop/tlb.scala 43:30]
  reg [1:0] pte_level_13; // @[playground/src/noop/tlb.scala 43:30]
  reg [1:0] pte_level_14; // @[playground/src/noop/tlb.scala 43:30]
  reg [1:0] pte_level_15; // @[playground/src/noop/tlb.scala 43:30]
  reg  valid_0; // @[playground/src/noop/tlb.scala 44:26]
  reg  valid_1; // @[playground/src/noop/tlb.scala 44:26]
  reg  valid_2; // @[playground/src/noop/tlb.scala 44:26]
  reg  valid_3; // @[playground/src/noop/tlb.scala 44:26]
  reg  valid_4; // @[playground/src/noop/tlb.scala 44:26]
  reg  valid_5; // @[playground/src/noop/tlb.scala 44:26]
  reg  valid_6; // @[playground/src/noop/tlb.scala 44:26]
  reg  valid_7; // @[playground/src/noop/tlb.scala 44:26]
  reg  valid_8; // @[playground/src/noop/tlb.scala 44:26]
  reg  valid_9; // @[playground/src/noop/tlb.scala 44:26]
  reg  valid_10; // @[playground/src/noop/tlb.scala 44:26]
  reg  valid_11; // @[playground/src/noop/tlb.scala 44:26]
  reg  valid_12; // @[playground/src/noop/tlb.scala 44:26]
  reg  valid_13; // @[playground/src/noop/tlb.scala 44:26]
  reg  valid_14; // @[playground/src/noop/tlb.scala 44:26]
  reg  valid_15; // @[playground/src/noop/tlb.scala 44:26]
  reg [63:0] pre_addr; // @[playground/src/noop/tlb.scala 46:30]
  reg [31:0] pte_addr_r; // @[playground/src/noop/tlb.scala 47:30]
  reg [63:0] wpte_data_r; // @[playground/src/noop/tlb.scala 48:30]
  reg [4:0] dc_mode_r; // @[playground/src/noop/tlb.scala 49:30]
  reg  out_valid_r; // @[playground/src/noop/tlb.scala 51:30]
  reg [31:0] out_paddr_r; // @[playground/src/noop/tlb.scala 52:30]
  reg [63:0] out_excep_r_cause; // @[playground/src/noop/tlb.scala 53:30]
  reg [63:0] out_excep_r_tval; // @[playground/src/noop/tlb.scala 53:30]
  reg  out_excep_r_en; // @[playground/src/noop/tlb.scala 53:30]
  wire [51:0] inp_tag = io_va2pa_vaddr[63:12]; // @[playground/src/noop/tlb.scala 58:33]
  wire [3:0] mmuMode = io_mmuState_priv == 2'h3 ? 4'h0 : io_mmuState_satp[63:60]; // @[playground/src/noop/tlb.scala 65:22]
  wire  is_Sv39 = mmuMode == 4'h8; // @[playground/src/noop/tlb.scala 66:27]
  wire [51:0] _tlb_tag_mask_T_4 = 2'h0 == pte_level_0 ? 52'hfffffffffffff : 52'h0; // @[src/main/scala/chisel3/util/Mux.scala 81:58]
  wire [51:0] _tlb_tag_mask_T_6 = 2'h1 == pte_level_0 ? 52'hffffffffffe00 : _tlb_tag_mask_T_4; // @[src/main/scala/chisel3/util/Mux.scala 81:58]
  wire [51:0] tlb_tag_mask = 2'h2 == pte_level_0 ? 52'hffffffffc0000 : _tlb_tag_mask_T_6; // @[src/main/scala/chisel3/util/Mux.scala 81:58]
  wire [51:0] _T_1 = inp_tag & tlb_tag_mask; // @[playground/src/noop/tlb.scala 73:24]
  wire [19:0] _GEN_2 = _T_1 == tag_0 & valid_0 ? paddr_0 : 20'h0; // @[playground/src/noop/tlb.scala 73:64 75:28 68:40]
  wire [9:0] _GEN_4 = _T_1 == tag_0 & valid_0 ? info_0 : 10'h0; // @[playground/src/noop/tlb.scala 73:64 77:28 68:86]
  wire [31:0] _GEN_5 = _T_1 == tag_0 & valid_0 ? pte_addr_0 : 32'h0; // @[playground/src/noop/tlb.scala 69:23 73:64 78:31]
  wire [1:0] _GEN_7 = _T_1 == tag_0 & valid_0 ? pte_level_0 : 2'h0; // @[playground/src/noop/tlb.scala 73:64 80:31 69:69]
  wire [51:0] _tlb_tag_mask_T_12 = 2'h0 == pte_level_1 ? 52'hfffffffffffff : 52'h0; // @[src/main/scala/chisel3/util/Mux.scala 81:58]
  wire [51:0] _tlb_tag_mask_T_14 = 2'h1 == pte_level_1 ? 52'hffffffffffe00 : _tlb_tag_mask_T_12; // @[src/main/scala/chisel3/util/Mux.scala 81:58]
  wire [51:0] tlb_tag_mask_1 = 2'h2 == pte_level_1 ? 52'hffffffffc0000 : _tlb_tag_mask_T_14; // @[src/main/scala/chisel3/util/Mux.scala 81:58]
  wire [51:0] _T_4 = inp_tag & tlb_tag_mask_1; // @[playground/src/noop/tlb.scala 73:24]
  wire  _T_6 = _T_4 == tag_1 & valid_1; // @[playground/src/noop/tlb.scala 73:52]
  wire [19:0] _GEN_9 = _T_4 == tag_1 & valid_1 ? paddr_1 : _GEN_2; // @[playground/src/noop/tlb.scala 73:64 75:28]
  wire [9:0] _GEN_11 = _T_4 == tag_1 & valid_1 ? info_1 : _GEN_4; // @[playground/src/noop/tlb.scala 73:64 77:28]
  wire [31:0] _GEN_12 = _T_4 == tag_1 & valid_1 ? pte_addr_1 : _GEN_5; // @[playground/src/noop/tlb.scala 73:64 78:31]
  wire [1:0] _GEN_14 = _T_4 == tag_1 & valid_1 ? pte_level_1 : _GEN_7; // @[playground/src/noop/tlb.scala 73:64 80:31]
  wire [51:0] _tlb_tag_mask_T_20 = 2'h0 == pte_level_2 ? 52'hfffffffffffff : 52'h0; // @[src/main/scala/chisel3/util/Mux.scala 81:58]
  wire [51:0] _tlb_tag_mask_T_22 = 2'h1 == pte_level_2 ? 52'hffffffffffe00 : _tlb_tag_mask_T_20; // @[src/main/scala/chisel3/util/Mux.scala 81:58]
  wire [51:0] tlb_tag_mask_2 = 2'h2 == pte_level_2 ? 52'hffffffffc0000 : _tlb_tag_mask_T_22; // @[src/main/scala/chisel3/util/Mux.scala 81:58]
  wire [51:0] _T_7 = inp_tag & tlb_tag_mask_2; // @[playground/src/noop/tlb.scala 73:24]
  wire [19:0] _GEN_16 = _T_7 == tag_2 & valid_2 ? paddr_2 : _GEN_9; // @[playground/src/noop/tlb.scala 73:64 75:28]
  wire [9:0] _GEN_18 = _T_7 == tag_2 & valid_2 ? info_2 : _GEN_11; // @[playground/src/noop/tlb.scala 73:64 77:28]
  wire [31:0] _GEN_19 = _T_7 == tag_2 & valid_2 ? pte_addr_2 : _GEN_12; // @[playground/src/noop/tlb.scala 73:64 78:31]
  wire [1:0] _GEN_20 = _T_7 == tag_2 & valid_2 ? 2'h2 : {{1'd0}, _T_6}; // @[playground/src/noop/tlb.scala 73:64 79:28]
  wire [1:0] _GEN_21 = _T_7 == tag_2 & valid_2 ? pte_level_2 : _GEN_14; // @[playground/src/noop/tlb.scala 73:64 80:31]
  wire [51:0] _tlb_tag_mask_T_28 = 2'h0 == pte_level_3 ? 52'hfffffffffffff : 52'h0; // @[src/main/scala/chisel3/util/Mux.scala 81:58]
  wire [51:0] _tlb_tag_mask_T_30 = 2'h1 == pte_level_3 ? 52'hffffffffffe00 : _tlb_tag_mask_T_28; // @[src/main/scala/chisel3/util/Mux.scala 81:58]
  wire [51:0] tlb_tag_mask_3 = 2'h2 == pte_level_3 ? 52'hffffffffc0000 : _tlb_tag_mask_T_30; // @[src/main/scala/chisel3/util/Mux.scala 81:58]
  wire [51:0] _T_10 = inp_tag & tlb_tag_mask_3; // @[playground/src/noop/tlb.scala 73:24]
  wire [19:0] _GEN_23 = _T_10 == tag_3 & valid_3 ? paddr_3 : _GEN_16; // @[playground/src/noop/tlb.scala 73:64 75:28]
  wire [9:0] _GEN_25 = _T_10 == tag_3 & valid_3 ? info_3 : _GEN_18; // @[playground/src/noop/tlb.scala 73:64 77:28]
  wire [31:0] _GEN_26 = _T_10 == tag_3 & valid_3 ? pte_addr_3 : _GEN_19; // @[playground/src/noop/tlb.scala 73:64 78:31]
  wire [1:0] _GEN_27 = _T_10 == tag_3 & valid_3 ? 2'h3 : _GEN_20; // @[playground/src/noop/tlb.scala 73:64 79:28]
  wire [1:0] _GEN_28 = _T_10 == tag_3 & valid_3 ? pte_level_3 : _GEN_21; // @[playground/src/noop/tlb.scala 73:64 80:31]
  wire [51:0] _tlb_tag_mask_T_36 = 2'h0 == pte_level_4 ? 52'hfffffffffffff : 52'h0; // @[src/main/scala/chisel3/util/Mux.scala 81:58]
  wire [51:0] _tlb_tag_mask_T_38 = 2'h1 == pte_level_4 ? 52'hffffffffffe00 : _tlb_tag_mask_T_36; // @[src/main/scala/chisel3/util/Mux.scala 81:58]
  wire [51:0] tlb_tag_mask_4 = 2'h2 == pte_level_4 ? 52'hffffffffc0000 : _tlb_tag_mask_T_38; // @[src/main/scala/chisel3/util/Mux.scala 81:58]
  wire [51:0] _T_13 = inp_tag & tlb_tag_mask_4; // @[playground/src/noop/tlb.scala 73:24]
  wire [19:0] _GEN_30 = _T_13 == tag_4 & valid_4 ? paddr_4 : _GEN_23; // @[playground/src/noop/tlb.scala 73:64 75:28]
  wire [9:0] _GEN_32 = _T_13 == tag_4 & valid_4 ? info_4 : _GEN_25; // @[playground/src/noop/tlb.scala 73:64 77:28]
  wire [31:0] _GEN_33 = _T_13 == tag_4 & valid_4 ? pte_addr_4 : _GEN_26; // @[playground/src/noop/tlb.scala 73:64 78:31]
  wire [2:0] _GEN_34 = _T_13 == tag_4 & valid_4 ? 3'h4 : {{1'd0}, _GEN_27}; // @[playground/src/noop/tlb.scala 73:64 79:28]
  wire [1:0] _GEN_35 = _T_13 == tag_4 & valid_4 ? pte_level_4 : _GEN_28; // @[playground/src/noop/tlb.scala 73:64 80:31]
  wire [51:0] _tlb_tag_mask_T_44 = 2'h0 == pte_level_5 ? 52'hfffffffffffff : 52'h0; // @[src/main/scala/chisel3/util/Mux.scala 81:58]
  wire [51:0] _tlb_tag_mask_T_46 = 2'h1 == pte_level_5 ? 52'hffffffffffe00 : _tlb_tag_mask_T_44; // @[src/main/scala/chisel3/util/Mux.scala 81:58]
  wire [51:0] tlb_tag_mask_5 = 2'h2 == pte_level_5 ? 52'hffffffffc0000 : _tlb_tag_mask_T_46; // @[src/main/scala/chisel3/util/Mux.scala 81:58]
  wire [51:0] _T_16 = inp_tag & tlb_tag_mask_5; // @[playground/src/noop/tlb.scala 73:24]
  wire [19:0] _GEN_37 = _T_16 == tag_5 & valid_5 ? paddr_5 : _GEN_30; // @[playground/src/noop/tlb.scala 73:64 75:28]
  wire [9:0] _GEN_39 = _T_16 == tag_5 & valid_5 ? info_5 : _GEN_32; // @[playground/src/noop/tlb.scala 73:64 77:28]
  wire [31:0] _GEN_40 = _T_16 == tag_5 & valid_5 ? pte_addr_5 : _GEN_33; // @[playground/src/noop/tlb.scala 73:64 78:31]
  wire [2:0] _GEN_41 = _T_16 == tag_5 & valid_5 ? 3'h5 : _GEN_34; // @[playground/src/noop/tlb.scala 73:64 79:28]
  wire [1:0] _GEN_42 = _T_16 == tag_5 & valid_5 ? pte_level_5 : _GEN_35; // @[playground/src/noop/tlb.scala 73:64 80:31]
  wire [51:0] _tlb_tag_mask_T_52 = 2'h0 == pte_level_6 ? 52'hfffffffffffff : 52'h0; // @[src/main/scala/chisel3/util/Mux.scala 81:58]
  wire [51:0] _tlb_tag_mask_T_54 = 2'h1 == pte_level_6 ? 52'hffffffffffe00 : _tlb_tag_mask_T_52; // @[src/main/scala/chisel3/util/Mux.scala 81:58]
  wire [51:0] tlb_tag_mask_6 = 2'h2 == pte_level_6 ? 52'hffffffffc0000 : _tlb_tag_mask_T_54; // @[src/main/scala/chisel3/util/Mux.scala 81:58]
  wire [51:0] _T_19 = inp_tag & tlb_tag_mask_6; // @[playground/src/noop/tlb.scala 73:24]
  wire [19:0] _GEN_44 = _T_19 == tag_6 & valid_6 ? paddr_6 : _GEN_37; // @[playground/src/noop/tlb.scala 73:64 75:28]
  wire [9:0] _GEN_46 = _T_19 == tag_6 & valid_6 ? info_6 : _GEN_39; // @[playground/src/noop/tlb.scala 73:64 77:28]
  wire [31:0] _GEN_47 = _T_19 == tag_6 & valid_6 ? pte_addr_6 : _GEN_40; // @[playground/src/noop/tlb.scala 73:64 78:31]
  wire [2:0] _GEN_48 = _T_19 == tag_6 & valid_6 ? 3'h6 : _GEN_41; // @[playground/src/noop/tlb.scala 73:64 79:28]
  wire [1:0] _GEN_49 = _T_19 == tag_6 & valid_6 ? pte_level_6 : _GEN_42; // @[playground/src/noop/tlb.scala 73:64 80:31]
  wire [51:0] _tlb_tag_mask_T_60 = 2'h0 == pte_level_7 ? 52'hfffffffffffff : 52'h0; // @[src/main/scala/chisel3/util/Mux.scala 81:58]
  wire [51:0] _tlb_tag_mask_T_62 = 2'h1 == pte_level_7 ? 52'hffffffffffe00 : _tlb_tag_mask_T_60; // @[src/main/scala/chisel3/util/Mux.scala 81:58]
  wire [51:0] tlb_tag_mask_7 = 2'h2 == pte_level_7 ? 52'hffffffffc0000 : _tlb_tag_mask_T_62; // @[src/main/scala/chisel3/util/Mux.scala 81:58]
  wire [51:0] _T_22 = inp_tag & tlb_tag_mask_7; // @[playground/src/noop/tlb.scala 73:24]
  wire [19:0] _GEN_51 = _T_22 == tag_7 & valid_7 ? paddr_7 : _GEN_44; // @[playground/src/noop/tlb.scala 73:64 75:28]
  wire [9:0] _GEN_53 = _T_22 == tag_7 & valid_7 ? info_7 : _GEN_46; // @[playground/src/noop/tlb.scala 73:64 77:28]
  wire [31:0] _GEN_54 = _T_22 == tag_7 & valid_7 ? pte_addr_7 : _GEN_47; // @[playground/src/noop/tlb.scala 73:64 78:31]
  wire [2:0] _GEN_55 = _T_22 == tag_7 & valid_7 ? 3'h7 : _GEN_48; // @[playground/src/noop/tlb.scala 73:64 79:28]
  wire [1:0] _GEN_56 = _T_22 == tag_7 & valid_7 ? pte_level_7 : _GEN_49; // @[playground/src/noop/tlb.scala 73:64 80:31]
  wire [51:0] _tlb_tag_mask_T_68 = 2'h0 == pte_level_8 ? 52'hfffffffffffff : 52'h0; // @[src/main/scala/chisel3/util/Mux.scala 81:58]
  wire [51:0] _tlb_tag_mask_T_70 = 2'h1 == pte_level_8 ? 52'hffffffffffe00 : _tlb_tag_mask_T_68; // @[src/main/scala/chisel3/util/Mux.scala 81:58]
  wire [51:0] tlb_tag_mask_8 = 2'h2 == pte_level_8 ? 52'hffffffffc0000 : _tlb_tag_mask_T_70; // @[src/main/scala/chisel3/util/Mux.scala 81:58]
  wire [51:0] _T_25 = inp_tag & tlb_tag_mask_8; // @[playground/src/noop/tlb.scala 73:24]
  wire [19:0] _GEN_58 = _T_25 == tag_8 & valid_8 ? paddr_8 : _GEN_51; // @[playground/src/noop/tlb.scala 73:64 75:28]
  wire [9:0] _GEN_60 = _T_25 == tag_8 & valid_8 ? info_8 : _GEN_53; // @[playground/src/noop/tlb.scala 73:64 77:28]
  wire [31:0] _GEN_61 = _T_25 == tag_8 & valid_8 ? pte_addr_8 : _GEN_54; // @[playground/src/noop/tlb.scala 73:64 78:31]
  wire [3:0] _GEN_62 = _T_25 == tag_8 & valid_8 ? 4'h8 : {{1'd0}, _GEN_55}; // @[playground/src/noop/tlb.scala 73:64 79:28]
  wire [1:0] _GEN_63 = _T_25 == tag_8 & valid_8 ? pte_level_8 : _GEN_56; // @[playground/src/noop/tlb.scala 73:64 80:31]
  wire [51:0] _tlb_tag_mask_T_76 = 2'h0 == pte_level_9 ? 52'hfffffffffffff : 52'h0; // @[src/main/scala/chisel3/util/Mux.scala 81:58]
  wire [51:0] _tlb_tag_mask_T_78 = 2'h1 == pte_level_9 ? 52'hffffffffffe00 : _tlb_tag_mask_T_76; // @[src/main/scala/chisel3/util/Mux.scala 81:58]
  wire [51:0] tlb_tag_mask_9 = 2'h2 == pte_level_9 ? 52'hffffffffc0000 : _tlb_tag_mask_T_78; // @[src/main/scala/chisel3/util/Mux.scala 81:58]
  wire [51:0] _T_28 = inp_tag & tlb_tag_mask_9; // @[playground/src/noop/tlb.scala 73:24]
  wire  _GEN_64 = _T_28 == tag_9 & valid_9 | (_T_25 == tag_8 & valid_8 | (_T_22 == tag_7 & valid_7 | (_T_19 == tag_6 &
    valid_6 | (_T_16 == tag_5 & valid_5 | (_T_13 == tag_4 & valid_4 | (_T_10 == tag_3 & valid_3 | (_T_7 == tag_2 &
    valid_2 | (_T_4 == tag_1 & valid_1 | _T_1 == tag_0 & valid_0)))))))); // @[playground/src/noop/tlb.scala 73:64 74:28]
  wire [19:0] _GEN_65 = _T_28 == tag_9 & valid_9 ? paddr_9 : _GEN_58; // @[playground/src/noop/tlb.scala 73:64 75:28]
  wire [9:0] _GEN_67 = _T_28 == tag_9 & valid_9 ? info_9 : _GEN_60; // @[playground/src/noop/tlb.scala 73:64 77:28]
  wire [31:0] _GEN_68 = _T_28 == tag_9 & valid_9 ? pte_addr_9 : _GEN_61; // @[playground/src/noop/tlb.scala 73:64 78:31]
  wire [3:0] _GEN_69 = _T_28 == tag_9 & valid_9 ? 4'h9 : _GEN_62; // @[playground/src/noop/tlb.scala 73:64 79:28]
  wire [1:0] _GEN_70 = _T_28 == tag_9 & valid_9 ? pte_level_9 : _GEN_63; // @[playground/src/noop/tlb.scala 73:64 80:31]
  wire [51:0] _tlb_tag_mask_T_84 = 2'h0 == pte_level_10 ? 52'hfffffffffffff : 52'h0; // @[src/main/scala/chisel3/util/Mux.scala 81:58]
  wire [51:0] _tlb_tag_mask_T_86 = 2'h1 == pte_level_10 ? 52'hffffffffffe00 : _tlb_tag_mask_T_84; // @[src/main/scala/chisel3/util/Mux.scala 81:58]
  wire [51:0] tlb_tag_mask_10 = 2'h2 == pte_level_10 ? 52'hffffffffc0000 : _tlb_tag_mask_T_86; // @[src/main/scala/chisel3/util/Mux.scala 81:58]
  wire [51:0] _T_31 = inp_tag & tlb_tag_mask_10; // @[playground/src/noop/tlb.scala 73:24]
  wire [19:0] _GEN_72 = _T_31 == tag_10 & valid_10 ? paddr_10 : _GEN_65; // @[playground/src/noop/tlb.scala 73:64 75:28]
  wire [9:0] _GEN_74 = _T_31 == tag_10 & valid_10 ? info_10 : _GEN_67; // @[playground/src/noop/tlb.scala 73:64 77:28]
  wire [31:0] _GEN_75 = _T_31 == tag_10 & valid_10 ? pte_addr_10 : _GEN_68; // @[playground/src/noop/tlb.scala 73:64 78:31]
  wire [3:0] _GEN_76 = _T_31 == tag_10 & valid_10 ? 4'ha : _GEN_69; // @[playground/src/noop/tlb.scala 73:64 79:28]
  wire [1:0] _GEN_77 = _T_31 == tag_10 & valid_10 ? pte_level_10 : _GEN_70; // @[playground/src/noop/tlb.scala 73:64 80:31]
  wire [51:0] _tlb_tag_mask_T_92 = 2'h0 == pte_level_11 ? 52'hfffffffffffff : 52'h0; // @[src/main/scala/chisel3/util/Mux.scala 81:58]
  wire [51:0] _tlb_tag_mask_T_94 = 2'h1 == pte_level_11 ? 52'hffffffffffe00 : _tlb_tag_mask_T_92; // @[src/main/scala/chisel3/util/Mux.scala 81:58]
  wire [51:0] tlb_tag_mask_11 = 2'h2 == pte_level_11 ? 52'hffffffffc0000 : _tlb_tag_mask_T_94; // @[src/main/scala/chisel3/util/Mux.scala 81:58]
  wire [51:0] _T_34 = inp_tag & tlb_tag_mask_11; // @[playground/src/noop/tlb.scala 73:24]
  wire [19:0] _GEN_79 = _T_34 == tag_11 & valid_11 ? paddr_11 : _GEN_72; // @[playground/src/noop/tlb.scala 73:64 75:28]
  wire [9:0] _GEN_81 = _T_34 == tag_11 & valid_11 ? info_11 : _GEN_74; // @[playground/src/noop/tlb.scala 73:64 77:28]
  wire [31:0] _GEN_82 = _T_34 == tag_11 & valid_11 ? pte_addr_11 : _GEN_75; // @[playground/src/noop/tlb.scala 73:64 78:31]
  wire [3:0] _GEN_83 = _T_34 == tag_11 & valid_11 ? 4'hb : _GEN_76; // @[playground/src/noop/tlb.scala 73:64 79:28]
  wire [1:0] _GEN_84 = _T_34 == tag_11 & valid_11 ? pte_level_11 : _GEN_77; // @[playground/src/noop/tlb.scala 73:64 80:31]
  wire [51:0] _tlb_tag_mask_T_100 = 2'h0 == pte_level_12 ? 52'hfffffffffffff : 52'h0; // @[src/main/scala/chisel3/util/Mux.scala 81:58]
  wire [51:0] _tlb_tag_mask_T_102 = 2'h1 == pte_level_12 ? 52'hffffffffffe00 : _tlb_tag_mask_T_100; // @[src/main/scala/chisel3/util/Mux.scala 81:58]
  wire [51:0] tlb_tag_mask_12 = 2'h2 == pte_level_12 ? 52'hffffffffc0000 : _tlb_tag_mask_T_102; // @[src/main/scala/chisel3/util/Mux.scala 81:58]
  wire [51:0] _T_37 = inp_tag & tlb_tag_mask_12; // @[playground/src/noop/tlb.scala 73:24]
  wire [19:0] _GEN_86 = _T_37 == tag_12 & valid_12 ? paddr_12 : _GEN_79; // @[playground/src/noop/tlb.scala 73:64 75:28]
  wire [9:0] _GEN_88 = _T_37 == tag_12 & valid_12 ? info_12 : _GEN_81; // @[playground/src/noop/tlb.scala 73:64 77:28]
  wire [31:0] _GEN_89 = _T_37 == tag_12 & valid_12 ? pte_addr_12 : _GEN_82; // @[playground/src/noop/tlb.scala 73:64 78:31]
  wire [3:0] _GEN_90 = _T_37 == tag_12 & valid_12 ? 4'hc : _GEN_83; // @[playground/src/noop/tlb.scala 73:64 79:28]
  wire [1:0] _GEN_91 = _T_37 == tag_12 & valid_12 ? pte_level_12 : _GEN_84; // @[playground/src/noop/tlb.scala 73:64 80:31]
  wire [51:0] _tlb_tag_mask_T_108 = 2'h0 == pte_level_13 ? 52'hfffffffffffff : 52'h0; // @[src/main/scala/chisel3/util/Mux.scala 81:58]
  wire [51:0] _tlb_tag_mask_T_110 = 2'h1 == pte_level_13 ? 52'hffffffffffe00 : _tlb_tag_mask_T_108; // @[src/main/scala/chisel3/util/Mux.scala 81:58]
  wire [51:0] tlb_tag_mask_13 = 2'h2 == pte_level_13 ? 52'hffffffffc0000 : _tlb_tag_mask_T_110; // @[src/main/scala/chisel3/util/Mux.scala 81:58]
  wire [51:0] _T_40 = inp_tag & tlb_tag_mask_13; // @[playground/src/noop/tlb.scala 73:24]
  wire [19:0] _GEN_93 = _T_40 == tag_13 & valid_13 ? paddr_13 : _GEN_86; // @[playground/src/noop/tlb.scala 73:64 75:28]
  wire [9:0] _GEN_95 = _T_40 == tag_13 & valid_13 ? info_13 : _GEN_88; // @[playground/src/noop/tlb.scala 73:64 77:28]
  wire [31:0] _GEN_96 = _T_40 == tag_13 & valid_13 ? pte_addr_13 : _GEN_89; // @[playground/src/noop/tlb.scala 73:64 78:31]
  wire [3:0] _GEN_97 = _T_40 == tag_13 & valid_13 ? 4'hd : _GEN_90; // @[playground/src/noop/tlb.scala 73:64 79:28]
  wire [1:0] _GEN_98 = _T_40 == tag_13 & valid_13 ? pte_level_13 : _GEN_91; // @[playground/src/noop/tlb.scala 73:64 80:31]
  wire [51:0] _tlb_tag_mask_T_116 = 2'h0 == pte_level_14 ? 52'hfffffffffffff : 52'h0; // @[src/main/scala/chisel3/util/Mux.scala 81:58]
  wire [51:0] _tlb_tag_mask_T_118 = 2'h1 == pte_level_14 ? 52'hffffffffffe00 : _tlb_tag_mask_T_116; // @[src/main/scala/chisel3/util/Mux.scala 81:58]
  wire [51:0] tlb_tag_mask_14 = 2'h2 == pte_level_14 ? 52'hffffffffc0000 : _tlb_tag_mask_T_118; // @[src/main/scala/chisel3/util/Mux.scala 81:58]
  wire [51:0] _T_43 = inp_tag & tlb_tag_mask_14; // @[playground/src/noop/tlb.scala 73:24]
  wire [19:0] _GEN_100 = _T_43 == tag_14 & valid_14 ? paddr_14 : _GEN_93; // @[playground/src/noop/tlb.scala 73:64 75:28]
  wire [9:0] _GEN_102 = _T_43 == tag_14 & valid_14 ? info_14 : _GEN_95; // @[playground/src/noop/tlb.scala 73:64 77:28]
  wire [31:0] _GEN_103 = _T_43 == tag_14 & valid_14 ? pte_addr_14 : _GEN_96; // @[playground/src/noop/tlb.scala 73:64 78:31]
  wire [3:0] _GEN_104 = _T_43 == tag_14 & valid_14 ? 4'he : _GEN_97; // @[playground/src/noop/tlb.scala 73:64 79:28]
  wire [1:0] _GEN_105 = _T_43 == tag_14 & valid_14 ? pte_level_14 : _GEN_98; // @[playground/src/noop/tlb.scala 73:64 80:31]
  wire [51:0] _tlb_tag_mask_T_124 = 2'h0 == pte_level_15 ? 52'hfffffffffffff : 52'h0; // @[src/main/scala/chisel3/util/Mux.scala 81:58]
  wire [51:0] _tlb_tag_mask_T_126 = 2'h1 == pte_level_15 ? 52'hffffffffffe00 : _tlb_tag_mask_T_124; // @[src/main/scala/chisel3/util/Mux.scala 81:58]
  wire [51:0] tlb_tag_mask_15 = 2'h2 == pte_level_15 ? 52'hffffffffc0000 : _tlb_tag_mask_T_126; // @[src/main/scala/chisel3/util/Mux.scala 81:58]
  wire [51:0] _T_46 = inp_tag & tlb_tag_mask_15; // @[playground/src/noop/tlb.scala 73:24]
  wire  tlbMsg_tlbHit = _T_46 == tag_15 & valid_15 | (_T_43 == tag_14 & valid_14 | (_T_40 == tag_13 & valid_13 | (_T_37
     == tag_12 & valid_12 | (_T_34 == tag_11 & valid_11 | (_T_31 == tag_10 & valid_10 | _GEN_64))))); // @[playground/src/noop/tlb.scala 73:64 74:28]
  wire [19:0] tlbMsg_tlbPa = _T_46 == tag_15 & valid_15 ? paddr_15 : _GEN_100; // @[playground/src/noop/tlb.scala 73:64 75:28]
  wire [9:0] tlbMsg_tlbInfo = _T_46 == tag_15 & valid_15 ? info_15 : _GEN_102; // @[playground/src/noop/tlb.scala 73:64 77:28]
  wire [31:0] tlbMsg_tlbPteAddr = _T_46 == tag_15 & valid_15 ? pte_addr_15 : _GEN_103; // @[playground/src/noop/tlb.scala 73:64 78:31]
  wire [3:0] tlbMsg_tlbIdx = _T_46 == tag_15 & valid_15 ? 4'hf : _GEN_104; // @[playground/src/noop/tlb.scala 73:64 79:28]
  wire [1:0] tlbMsg_tlbLevel = _T_46 == tag_15 & valid_15 ? pte_level_15 : _GEN_105; // @[playground/src/noop/tlb.scala 73:64 80:31]
  reg [1:0] state; // @[playground/src/noop/tlb.scala 84:24]
  reg  flush_r; // @[playground/src/noop/tlb.scala 85:26]
  wire  _T_50 = state == 2'h0; // @[playground/src/noop/tlb.scala 87:20]
  wire  _GEN_113 = state == 2'h0 ? 1'h0 : valid_0; // @[playground/src/noop/tlb.scala 87:30 88:19 44:26]
  wire  _GEN_114 = state == 2'h0 ? 1'h0 : valid_1; // @[playground/src/noop/tlb.scala 87:30 88:19 44:26]
  wire  _GEN_115 = state == 2'h0 ? 1'h0 : valid_2; // @[playground/src/noop/tlb.scala 87:30 88:19 44:26]
  wire  _GEN_116 = state == 2'h0 ? 1'h0 : valid_3; // @[playground/src/noop/tlb.scala 87:30 88:19 44:26]
  wire  _GEN_117 = state == 2'h0 ? 1'h0 : valid_4; // @[playground/src/noop/tlb.scala 87:30 88:19 44:26]
  wire  _GEN_118 = state == 2'h0 ? 1'h0 : valid_5; // @[playground/src/noop/tlb.scala 87:30 88:19 44:26]
  wire  _GEN_119 = state == 2'h0 ? 1'h0 : valid_6; // @[playground/src/noop/tlb.scala 87:30 88:19 44:26]
  wire  _GEN_120 = state == 2'h0 ? 1'h0 : valid_7; // @[playground/src/noop/tlb.scala 87:30 88:19 44:26]
  wire  _GEN_121 = state == 2'h0 ? 1'h0 : valid_8; // @[playground/src/noop/tlb.scala 87:30 88:19 44:26]
  wire  _GEN_122 = state == 2'h0 ? 1'h0 : valid_9; // @[playground/src/noop/tlb.scala 87:30 88:19 44:26]
  wire  _GEN_123 = state == 2'h0 ? 1'h0 : valid_10; // @[playground/src/noop/tlb.scala 87:30 88:19 44:26]
  wire  _GEN_124 = state == 2'h0 ? 1'h0 : valid_11; // @[playground/src/noop/tlb.scala 87:30 88:19 44:26]
  wire  _GEN_125 = state == 2'h0 ? 1'h0 : valid_12; // @[playground/src/noop/tlb.scala 87:30 88:19 44:26]
  wire  _GEN_126 = state == 2'h0 ? 1'h0 : valid_13; // @[playground/src/noop/tlb.scala 87:30 88:19 44:26]
  wire  _GEN_127 = state == 2'h0 ? 1'h0 : valid_14; // @[playground/src/noop/tlb.scala 87:30 88:19 44:26]
  wire  _GEN_128 = state == 2'h0 ? 1'h0 : valid_15; // @[playground/src/noop/tlb.scala 87:30 88:19 44:26]
  wire  _GEN_130 = io_flush | flush_r ? _GEN_113 : valid_0; // @[playground/src/noop/tlb.scala 44:26 86:30]
  wire  _GEN_131 = io_flush | flush_r ? _GEN_114 : valid_1; // @[playground/src/noop/tlb.scala 44:26 86:30]
  wire  _GEN_132 = io_flush | flush_r ? _GEN_115 : valid_2; // @[playground/src/noop/tlb.scala 44:26 86:30]
  wire  _GEN_133 = io_flush | flush_r ? _GEN_116 : valid_3; // @[playground/src/noop/tlb.scala 44:26 86:30]
  wire  _GEN_134 = io_flush | flush_r ? _GEN_117 : valid_4; // @[playground/src/noop/tlb.scala 44:26 86:30]
  wire  _GEN_135 = io_flush | flush_r ? _GEN_118 : valid_5; // @[playground/src/noop/tlb.scala 44:26 86:30]
  wire  _GEN_136 = io_flush | flush_r ? _GEN_119 : valid_6; // @[playground/src/noop/tlb.scala 44:26 86:30]
  wire  _GEN_137 = io_flush | flush_r ? _GEN_120 : valid_7; // @[playground/src/noop/tlb.scala 44:26 86:30]
  wire  _GEN_138 = io_flush | flush_r ? _GEN_121 : valid_8; // @[playground/src/noop/tlb.scala 44:26 86:30]
  wire  _GEN_139 = io_flush | flush_r ? _GEN_122 : valid_9; // @[playground/src/noop/tlb.scala 44:26 86:30]
  wire  _GEN_140 = io_flush | flush_r ? _GEN_123 : valid_10; // @[playground/src/noop/tlb.scala 44:26 86:30]
  wire  _GEN_141 = io_flush | flush_r ? _GEN_124 : valid_11; // @[playground/src/noop/tlb.scala 44:26 86:30]
  wire  _GEN_142 = io_flush | flush_r ? _GEN_125 : valid_12; // @[playground/src/noop/tlb.scala 44:26 86:30]
  wire  _GEN_143 = io_flush | flush_r ? _GEN_126 : valid_13; // @[playground/src/noop/tlb.scala 44:26 86:30]
  wire  _GEN_144 = io_flush | flush_r ? _GEN_127 : valid_14; // @[playground/src/noop/tlb.scala 44:26 86:30]
  wire  _GEN_145 = io_flush | flush_r ? _GEN_128 : valid_15; // @[playground/src/noop/tlb.scala 44:26 86:30]
  wire  handshake = io_va2pa_vvalid & io_va2pa_ready; // @[playground/src/noop/tlb.scala 94:37]
  reg [1:0] m_type_r; // @[playground/src/noop/tlb.scala 95:27]
  wire [1:0] cur_m_type = handshake ? 2'h1 : m_type_r; // @[playground/src/noop/tlb.scala 96:25]
  wire  _ad_T = cur_m_type == 2'h3; // @[playground/src/noop/common.scala 243:20]
  wire [9:0] ad = cur_m_type == 2'h3 ? 10'hc0 : 10'h40; // @[playground/src/noop/common.scala 243:12]
  wire  _GEN_150 = io_va2pa_pvalid | io_va2pa_tlb_excep_en ? 1'h0 : out_valid_r; // @[playground/src/noop/tlb.scala 108:51 109:21 51:30]
  wire  _GEN_151 = io_va2pa_pvalid | io_va2pa_tlb_excep_en ? 1'h0 : out_excep_r_en; // @[playground/src/noop/tlb.scala 108:51 110:24 53:30]
  wire  dc_hand = io_dcacheRW_ready & io_dcacheRW_dc_mode != 5'h0; // @[playground/src/noop/tlb.scala 122:37]
  wire [24:0] _tlb_high_legal_T_2 = io_va2pa_vaddr[38] ? 25'h1ffffff : 25'h0; // @[playground/src/noop/tlb.scala 125:30]
  wire  tlb_high_legal = _tlb_high_legal_T_2 == io_va2pa_vaddr[63:39]; // @[playground/src/noop/tlb.scala 125:55]
  wire  _tlb_access_illegal_T_11 = cur_m_type == 2'h2 & ~(tlbMsg_tlbInfo[1] | io_mmuState_mstatus[19] & tlbMsg_tlbInfo[3
    ]); // @[playground/src/noop/tlb.scala 127:60]
  wire  _tlb_access_illegal_T_12 = cur_m_type == 2'h1 & ~tlbMsg_tlbInfo[3] | _tlb_access_illegal_T_11; // @[playground/src/noop/tlb.scala 126:89]
  wire  _tlb_access_illegal_T_16 = _ad_T & ~tlbMsg_tlbInfo[2]; // @[playground/src/noop/tlb.scala 128:57]
  wire  tlb_access_illegal = _tlb_access_illegal_T_12 | _tlb_access_illegal_T_16; // @[playground/src/noop/tlb.scala 127:152]
  wire [3:0] select = {select_prng_io_out_3,select_prng_io_out_2,select_prng_io_out_1,select_prng_io_out_0}; // @[src/main/scala/chisel3/util/random/PRNG.scala 95:17]
  reg [3:0] select_r; // @[playground/src/noop/tlb.scala 130:27]
  reg [7:0] offset; // @[playground/src/noop/tlb.scala 131:26]
  reg [1:0] level; // @[playground/src/noop/tlb.scala 132:26]
  reg  wpte_hs_r; // @[playground/src/noop/tlb.scala 134:28]
  wire [51:0] _paddr_mask_T_4 = 2'h0 == tlbMsg_tlbLevel ? 52'hfffffffffffff : 52'h0; // @[src/main/scala/chisel3/util/Mux.scala 81:58]
  wire [51:0] _paddr_mask_T_6 = 2'h1 == tlbMsg_tlbLevel ? 52'hffffffffffe00 : _paddr_mask_T_4; // @[src/main/scala/chisel3/util/Mux.scala 81:58]
  wire [51:0] _paddr_mask_T_8 = 2'h2 == tlbMsg_tlbLevel ? 52'hffffffffc0000 : _paddr_mask_T_6; // @[src/main/scala/chisel3/util/Mux.scala 81:58]
  wire [63:0] paddr_mask = {_paddr_mask_T_8,12'h0}; // @[playground/src/noop/tlb.scala 147:41]
  wire [31:0] _out_paddr_r_T = {tlbMsg_tlbPa, 12'h0}; // @[playground/src/noop/tlb.scala 148:93]
  wire [63:0] _out_paddr_r_T_1 = ~paddr_mask; // @[playground/src/noop/common.scala 201:19]
  wire [63:0] _out_paddr_r_T_2 = io_va2pa_vaddr & _out_paddr_r_T_1; // @[playground/src/noop/common.scala 201:17]
  wire [63:0] _GEN_3 = {{32'd0}, _out_paddr_r_T}; // @[playground/src/noop/common.scala 201:36]
  wire [63:0] _out_paddr_r_T_3 = _GEN_3 & paddr_mask; // @[playground/src/noop/common.scala 201:36]
  wire [63:0] _out_paddr_r_T_4 = _out_paddr_r_T_2 | _out_paddr_r_T_3; // @[playground/src/noop/common.scala 201:26]
  wire [9:0] _T_59 = ad & tlbMsg_tlbInfo; // @[playground/src/noop/tlb.scala 149:30]
  wire [9:0] _wpte_data_r_T = tlbMsg_tlbInfo | ad; // @[playground/src/noop/tlb.scala 153:84]
  wire [63:0] _wpte_data_r_T_1 = {34'h0,tlbMsg_tlbPa,_wpte_data_r_T}; // @[playground/src/noop/tlb.scala 153:43]
  wire [9:0] _GEN_152 = 4'h0 == tlbMsg_tlbIdx ? _wpte_data_r_T : info_0; // @[playground/src/noop/tlb.scala 154:{45,45} 41:26]
  wire [9:0] _GEN_153 = 4'h1 == tlbMsg_tlbIdx ? _wpte_data_r_T : info_1; // @[playground/src/noop/tlb.scala 154:{45,45} 41:26]
  wire [9:0] _GEN_154 = 4'h2 == tlbMsg_tlbIdx ? _wpte_data_r_T : info_2; // @[playground/src/noop/tlb.scala 154:{45,45} 41:26]
  wire [9:0] _GEN_155 = 4'h3 == tlbMsg_tlbIdx ? _wpte_data_r_T : info_3; // @[playground/src/noop/tlb.scala 154:{45,45} 41:26]
  wire [9:0] _GEN_156 = 4'h4 == tlbMsg_tlbIdx ? _wpte_data_r_T : info_4; // @[playground/src/noop/tlb.scala 154:{45,45} 41:26]
  wire [9:0] _GEN_157 = 4'h5 == tlbMsg_tlbIdx ? _wpte_data_r_T : info_5; // @[playground/src/noop/tlb.scala 154:{45,45} 41:26]
  wire [9:0] _GEN_158 = 4'h6 == tlbMsg_tlbIdx ? _wpte_data_r_T : info_6; // @[playground/src/noop/tlb.scala 154:{45,45} 41:26]
  wire [9:0] _GEN_159 = 4'h7 == tlbMsg_tlbIdx ? _wpte_data_r_T : info_7; // @[playground/src/noop/tlb.scala 154:{45,45} 41:26]
  wire [9:0] _GEN_160 = 4'h8 == tlbMsg_tlbIdx ? _wpte_data_r_T : info_8; // @[playground/src/noop/tlb.scala 154:{45,45} 41:26]
  wire [9:0] _GEN_161 = 4'h9 == tlbMsg_tlbIdx ? _wpte_data_r_T : info_9; // @[playground/src/noop/tlb.scala 154:{45,45} 41:26]
  wire [9:0] _GEN_162 = 4'ha == tlbMsg_tlbIdx ? _wpte_data_r_T : info_10; // @[playground/src/noop/tlb.scala 154:{45,45} 41:26]
  wire [9:0] _GEN_163 = 4'hb == tlbMsg_tlbIdx ? _wpte_data_r_T : info_11; // @[playground/src/noop/tlb.scala 154:{45,45} 41:26]
  wire [9:0] _GEN_164 = 4'hc == tlbMsg_tlbIdx ? _wpte_data_r_T : info_12; // @[playground/src/noop/tlb.scala 154:{45,45} 41:26]
  wire [9:0] _GEN_165 = 4'hd == tlbMsg_tlbIdx ? _wpte_data_r_T : info_13; // @[playground/src/noop/tlb.scala 154:{45,45} 41:26]
  wire [9:0] _GEN_166 = 4'he == tlbMsg_tlbIdx ? _wpte_data_r_T : info_14; // @[playground/src/noop/tlb.scala 154:{45,45} 41:26]
  wire [9:0] _GEN_167 = 4'hf == tlbMsg_tlbIdx ? _wpte_data_r_T : info_15; // @[playground/src/noop/tlb.scala 154:{45,45} 41:26]
  wire [1:0] _GEN_168 = _T_59 != ad & is_Sv39 ? 2'h3 : state; // @[playground/src/noop/tlb.scala 149:66 150:31 84:24]
  wire  _GEN_169 = _T_59 != ad & is_Sv39 ? 1'h0 : wpte_hs_r; // @[playground/src/noop/tlb.scala 134:28 149:66 151:35]
  wire [31:0] _GEN_170 = _T_59 != ad & is_Sv39 ? tlbMsg_tlbPteAddr : pte_addr_r; // @[playground/src/noop/tlb.scala 149:66 152:37 47:30]
  wire [63:0] _GEN_171 = _T_59 != ad & is_Sv39 ? _wpte_data_r_T_1 : wpte_data_r; // @[playground/src/noop/tlb.scala 149:66 153:37 48:30]
  wire [9:0] _GEN_172 = _T_59 != ad & is_Sv39 ? _GEN_152 : info_0; // @[playground/src/noop/tlb.scala 149:66 41:26]
  wire [9:0] _GEN_173 = _T_59 != ad & is_Sv39 ? _GEN_153 : info_1; // @[playground/src/noop/tlb.scala 149:66 41:26]
  wire [9:0] _GEN_174 = _T_59 != ad & is_Sv39 ? _GEN_154 : info_2; // @[playground/src/noop/tlb.scala 149:66 41:26]
  wire [9:0] _GEN_175 = _T_59 != ad & is_Sv39 ? _GEN_155 : info_3; // @[playground/src/noop/tlb.scala 149:66 41:26]
  wire [9:0] _GEN_176 = _T_59 != ad & is_Sv39 ? _GEN_156 : info_4; // @[playground/src/noop/tlb.scala 149:66 41:26]
  wire [9:0] _GEN_177 = _T_59 != ad & is_Sv39 ? _GEN_157 : info_5; // @[playground/src/noop/tlb.scala 149:66 41:26]
  wire [9:0] _GEN_178 = _T_59 != ad & is_Sv39 ? _GEN_158 : info_6; // @[playground/src/noop/tlb.scala 149:66 41:26]
  wire [9:0] _GEN_179 = _T_59 != ad & is_Sv39 ? _GEN_159 : info_7; // @[playground/src/noop/tlb.scala 149:66 41:26]
  wire [9:0] _GEN_180 = _T_59 != ad & is_Sv39 ? _GEN_160 : info_8; // @[playground/src/noop/tlb.scala 149:66 41:26]
  wire [9:0] _GEN_181 = _T_59 != ad & is_Sv39 ? _GEN_161 : info_9; // @[playground/src/noop/tlb.scala 149:66 41:26]
  wire [9:0] _GEN_182 = _T_59 != ad & is_Sv39 ? _GEN_162 : info_10; // @[playground/src/noop/tlb.scala 149:66 41:26]
  wire [9:0] _GEN_183 = _T_59 != ad & is_Sv39 ? _GEN_163 : info_11; // @[playground/src/noop/tlb.scala 149:66 41:26]
  wire [9:0] _GEN_184 = _T_59 != ad & is_Sv39 ? _GEN_164 : info_12; // @[playground/src/noop/tlb.scala 149:66 41:26]
  wire [9:0] _GEN_185 = _T_59 != ad & is_Sv39 ? _GEN_165 : info_13; // @[playground/src/noop/tlb.scala 149:66 41:26]
  wire [9:0] _GEN_186 = _T_59 != ad & is_Sv39 ? _GEN_166 : info_14; // @[playground/src/noop/tlb.scala 149:66 41:26]
  wire [9:0] _GEN_187 = _T_59 != ad & is_Sv39 ? _GEN_167 : info_15; // @[playground/src/noop/tlb.scala 149:66 41:26]
  wire [63:0] _pte_addr_r_T_1 = {{30'd0}, io_va2pa_vaddr[63:30]}; // @[playground/src/noop/tlb.scala 166:83]
  wire [55:0] _pte_addr_r_T_3 = {io_mmuState_satp[43:0],_pte_addr_r_T_1[8:0],3'h0}; // @[playground/src/noop/tlb.scala 166:42]
  wire  _GEN_188 = io_va2pa_vaddr[63:39] != _tlb_high_legal_T_2 | _GEN_151; // @[playground/src/noop/tlb.scala 162:81 164:40]
  wire [55:0] _GEN_189 = io_va2pa_vaddr[63:39] != _tlb_high_legal_T_2 ? {{24'd0}, pte_addr_r} : _pte_addr_r_T_3; // @[playground/src/noop/tlb.scala 162:81 47:30 166:36]
  wire [4:0] _GEN_190 = io_va2pa_vaddr[63:39] != _tlb_high_legal_T_2 ? 5'h0 : 5'h7; // @[playground/src/noop/tlb.scala 138:27 162:81 167:36]
  wire [7:0] _GEN_191 = io_va2pa_vaddr[63:39] != _tlb_high_legal_T_2 ? offset : 8'h1e; // @[playground/src/noop/tlb.scala 131:26 162:81 168:33]
  wire [1:0] _GEN_192 = io_va2pa_vaddr[63:39] != _tlb_high_legal_T_2 ? level : 2'h3; // @[playground/src/noop/tlb.scala 132:26 162:81 169:33]
  wire [1:0] _GEN_194 = ~tlbMsg_tlbHit ? 2'h1 : state; // @[playground/src/noop/tlb.scala 156:43 84:24]
  wire [3:0] _GEN_195 = ~tlbMsg_tlbHit ? select : select_r; // @[playground/src/noop/tlb.scala 130:27 156:43 158:32]
  wire [1:0] _GEN_196 = ~tlbMsg_tlbHit ? 2'h1 : m_type_r; // @[playground/src/noop/tlb.scala 156:43 159:32 95:27]
  wire [63:0] _GEN_197 = ~tlbMsg_tlbHit ? 64'hc : out_excep_r_cause; // @[playground/src/noop/tlb.scala 156:43 160:39 53:30]
  wire [63:0] _GEN_198 = ~tlbMsg_tlbHit ? io_va2pa_vaddr : out_excep_r_tval; // @[playground/src/noop/tlb.scala 156:43 161:39 53:30]
  wire  _GEN_199 = ~tlbMsg_tlbHit ? _GEN_188 : _GEN_151; // @[playground/src/noop/tlb.scala 156:43]
  wire [55:0] _GEN_200 = ~tlbMsg_tlbHit ? _GEN_189 : {{24'd0}, pte_addr_r}; // @[playground/src/noop/tlb.scala 156:43 47:30]
  wire [4:0] _GEN_201 = ~tlbMsg_tlbHit ? _GEN_190 : 5'h0; // @[playground/src/noop/tlb.scala 138:27 156:43]
  wire [7:0] _GEN_202 = ~tlbMsg_tlbHit ? _GEN_191 : offset; // @[playground/src/noop/tlb.scala 131:26 156:43]
  wire [1:0] _GEN_203 = ~tlbMsg_tlbHit ? _GEN_192 : level; // @[playground/src/noop/tlb.scala 132:26 156:43]
  wire  _GEN_204 = tlbMsg_tlbHit | _GEN_150; // @[playground/src/noop/tlb.scala 144:42 145:33]
  wire [63:0] _GEN_205 = tlbMsg_tlbHit ? _out_paddr_r_T_4 : {{32'd0}, out_paddr_r}; // @[playground/src/noop/tlb.scala 144:42 148:33 52:30]
  wire [1:0] _GEN_206 = tlbMsg_tlbHit ? _GEN_168 : _GEN_194; // @[playground/src/noop/tlb.scala 144:42]
  wire  _GEN_207 = tlbMsg_tlbHit ? _GEN_169 : wpte_hs_r; // @[playground/src/noop/tlb.scala 134:28 144:42]
  wire [55:0] _GEN_208 = tlbMsg_tlbHit ? {{24'd0}, _GEN_170} : _GEN_200; // @[playground/src/noop/tlb.scala 144:42]
  wire [63:0] _GEN_209 = tlbMsg_tlbHit ? _GEN_171 : wpte_data_r; // @[playground/src/noop/tlb.scala 144:42 48:30]
  wire [9:0] _GEN_210 = tlbMsg_tlbHit ? _GEN_172 : info_0; // @[playground/src/noop/tlb.scala 144:42 41:26]
  wire [9:0] _GEN_211 = tlbMsg_tlbHit ? _GEN_173 : info_1; // @[playground/src/noop/tlb.scala 144:42 41:26]
  wire [9:0] _GEN_212 = tlbMsg_tlbHit ? _GEN_174 : info_2; // @[playground/src/noop/tlb.scala 144:42 41:26]
  wire [9:0] _GEN_213 = tlbMsg_tlbHit ? _GEN_175 : info_3; // @[playground/src/noop/tlb.scala 144:42 41:26]
  wire [9:0] _GEN_214 = tlbMsg_tlbHit ? _GEN_176 : info_4; // @[playground/src/noop/tlb.scala 144:42 41:26]
  wire [9:0] _GEN_215 = tlbMsg_tlbHit ? _GEN_177 : info_5; // @[playground/src/noop/tlb.scala 144:42 41:26]
  wire [9:0] _GEN_216 = tlbMsg_tlbHit ? _GEN_178 : info_6; // @[playground/src/noop/tlb.scala 144:42 41:26]
  wire [9:0] _GEN_217 = tlbMsg_tlbHit ? _GEN_179 : info_7; // @[playground/src/noop/tlb.scala 144:42 41:26]
  wire [9:0] _GEN_218 = tlbMsg_tlbHit ? _GEN_180 : info_8; // @[playground/src/noop/tlb.scala 144:42 41:26]
  wire [9:0] _GEN_219 = tlbMsg_tlbHit ? _GEN_181 : info_9; // @[playground/src/noop/tlb.scala 144:42 41:26]
  wire [9:0] _GEN_220 = tlbMsg_tlbHit ? _GEN_182 : info_10; // @[playground/src/noop/tlb.scala 144:42 41:26]
  wire [9:0] _GEN_221 = tlbMsg_tlbHit ? _GEN_183 : info_11; // @[playground/src/noop/tlb.scala 144:42 41:26]
  wire [9:0] _GEN_222 = tlbMsg_tlbHit ? _GEN_184 : info_12; // @[playground/src/noop/tlb.scala 144:42 41:26]
  wire [9:0] _GEN_223 = tlbMsg_tlbHit ? _GEN_185 : info_13; // @[playground/src/noop/tlb.scala 144:42 41:26]
  wire [9:0] _GEN_224 = tlbMsg_tlbHit ? _GEN_186 : info_14; // @[playground/src/noop/tlb.scala 144:42 41:26]
  wire [9:0] _GEN_225 = tlbMsg_tlbHit ? _GEN_187 : info_15; // @[playground/src/noop/tlb.scala 144:42 41:26]
  wire [3:0] _GEN_226 = tlbMsg_tlbHit ? select_r : _GEN_195; // @[playground/src/noop/tlb.scala 130:27 144:42]
  wire [1:0] _GEN_227 = tlbMsg_tlbHit ? m_type_r : _GEN_196; // @[playground/src/noop/tlb.scala 144:42 95:27]
  wire [63:0] _GEN_228 = tlbMsg_tlbHit ? out_excep_r_cause : _GEN_197; // @[playground/src/noop/tlb.scala 144:42 53:30]
  wire [63:0] _GEN_229 = tlbMsg_tlbHit ? out_excep_r_tval : _GEN_198; // @[playground/src/noop/tlb.scala 144:42 53:30]
  wire  _GEN_230 = tlbMsg_tlbHit ? _GEN_151 : _GEN_199; // @[playground/src/noop/tlb.scala 144:42]
  wire [4:0] _GEN_231 = tlbMsg_tlbHit ? 5'h0 : _GEN_201; // @[playground/src/noop/tlb.scala 138:27 144:42]
  wire [7:0] _GEN_232 = tlbMsg_tlbHit ? offset : _GEN_202; // @[playground/src/noop/tlb.scala 131:26 144:42]
  wire [1:0] _GEN_233 = tlbMsg_tlbHit ? level : _GEN_203; // @[playground/src/noop/tlb.scala 132:26 144:42]
  wire  _GEN_234 = ~tlb_high_legal | tlbMsg_tlbHit & tlb_access_illegal | _GEN_230; // @[playground/src/noop/tlb.scala 140:85 141:36]
  wire [63:0] _GEN_235 = ~tlb_high_legal | tlbMsg_tlbHit & tlb_access_illegal ? 64'hc : _GEN_228; // @[playground/src/noop/tlb.scala 140:85 142:39]
  wire [63:0] _GEN_236 = ~tlb_high_legal | tlbMsg_tlbHit & tlb_access_illegal ? io_va2pa_vaddr : _GEN_229; // @[playground/src/noop/tlb.scala 140:85 143:39]
  wire  _GEN_237 = ~tlb_high_legal | tlbMsg_tlbHit & tlb_access_illegal ? _GEN_150 : _GEN_204; // @[playground/src/noop/tlb.scala 140:85]
  wire [63:0] _GEN_238 = ~tlb_high_legal | tlbMsg_tlbHit & tlb_access_illegal ? {{32'd0}, out_paddr_r} : _GEN_205; // @[playground/src/noop/tlb.scala 140:85 52:30]
  wire [1:0] _GEN_239 = ~tlb_high_legal | tlbMsg_tlbHit & tlb_access_illegal ? state : _GEN_206; // @[playground/src/noop/tlb.scala 140:85 84:24]
  wire  _GEN_240 = ~tlb_high_legal | tlbMsg_tlbHit & tlb_access_illegal ? wpte_hs_r : _GEN_207; // @[playground/src/noop/tlb.scala 134:28 140:85]
  wire [55:0] _GEN_241 = ~tlb_high_legal | tlbMsg_tlbHit & tlb_access_illegal ? {{24'd0}, pte_addr_r} : _GEN_208; // @[playground/src/noop/tlb.scala 140:85 47:30]
  wire [63:0] _GEN_242 = ~tlb_high_legal | tlbMsg_tlbHit & tlb_access_illegal ? wpte_data_r : _GEN_209; // @[playground/src/noop/tlb.scala 140:85 48:30]
  wire [9:0] _GEN_243 = ~tlb_high_legal | tlbMsg_tlbHit & tlb_access_illegal ? info_0 : _GEN_210; // @[playground/src/noop/tlb.scala 140:85 41:26]
  wire [9:0] _GEN_244 = ~tlb_high_legal | tlbMsg_tlbHit & tlb_access_illegal ? info_1 : _GEN_211; // @[playground/src/noop/tlb.scala 140:85 41:26]
  wire [9:0] _GEN_245 = ~tlb_high_legal | tlbMsg_tlbHit & tlb_access_illegal ? info_2 : _GEN_212; // @[playground/src/noop/tlb.scala 140:85 41:26]
  wire [9:0] _GEN_246 = ~tlb_high_legal | tlbMsg_tlbHit & tlb_access_illegal ? info_3 : _GEN_213; // @[playground/src/noop/tlb.scala 140:85 41:26]
  wire [9:0] _GEN_247 = ~tlb_high_legal | tlbMsg_tlbHit & tlb_access_illegal ? info_4 : _GEN_214; // @[playground/src/noop/tlb.scala 140:85 41:26]
  wire [9:0] _GEN_248 = ~tlb_high_legal | tlbMsg_tlbHit & tlb_access_illegal ? info_5 : _GEN_215; // @[playground/src/noop/tlb.scala 140:85 41:26]
  wire [9:0] _GEN_249 = ~tlb_high_legal | tlbMsg_tlbHit & tlb_access_illegal ? info_6 : _GEN_216; // @[playground/src/noop/tlb.scala 140:85 41:26]
  wire [9:0] _GEN_250 = ~tlb_high_legal | tlbMsg_tlbHit & tlb_access_illegal ? info_7 : _GEN_217; // @[playground/src/noop/tlb.scala 140:85 41:26]
  wire [9:0] _GEN_251 = ~tlb_high_legal | tlbMsg_tlbHit & tlb_access_illegal ? info_8 : _GEN_218; // @[playground/src/noop/tlb.scala 140:85 41:26]
  wire [9:0] _GEN_252 = ~tlb_high_legal | tlbMsg_tlbHit & tlb_access_illegal ? info_9 : _GEN_219; // @[playground/src/noop/tlb.scala 140:85 41:26]
  wire [9:0] _GEN_253 = ~tlb_high_legal | tlbMsg_tlbHit & tlb_access_illegal ? info_10 : _GEN_220; // @[playground/src/noop/tlb.scala 140:85 41:26]
  wire [9:0] _GEN_254 = ~tlb_high_legal | tlbMsg_tlbHit & tlb_access_illegal ? info_11 : _GEN_221; // @[playground/src/noop/tlb.scala 140:85 41:26]
  wire [9:0] _GEN_255 = ~tlb_high_legal | tlbMsg_tlbHit & tlb_access_illegal ? info_12 : _GEN_222; // @[playground/src/noop/tlb.scala 140:85 41:26]
  wire [9:0] _GEN_256 = ~tlb_high_legal | tlbMsg_tlbHit & tlb_access_illegal ? info_13 : _GEN_223; // @[playground/src/noop/tlb.scala 140:85 41:26]
  wire [9:0] _GEN_257 = ~tlb_high_legal | tlbMsg_tlbHit & tlb_access_illegal ? info_14 : _GEN_224; // @[playground/src/noop/tlb.scala 140:85 41:26]
  wire [9:0] _GEN_258 = ~tlb_high_legal | tlbMsg_tlbHit & tlb_access_illegal ? info_15 : _GEN_225; // @[playground/src/noop/tlb.scala 140:85 41:26]
  wire [3:0] _GEN_259 = ~tlb_high_legal | tlbMsg_tlbHit & tlb_access_illegal ? select_r : _GEN_226; // @[playground/src/noop/tlb.scala 130:27 140:85]
  wire [1:0] _GEN_260 = ~tlb_high_legal | tlbMsg_tlbHit & tlb_access_illegal ? m_type_r : _GEN_227; // @[playground/src/noop/tlb.scala 140:85 95:27]
  wire [4:0] _GEN_261 = ~tlb_high_legal | tlbMsg_tlbHit & tlb_access_illegal ? 5'h0 : _GEN_231; // @[playground/src/noop/tlb.scala 138:27 140:85]
  wire [7:0] _GEN_262 = ~tlb_high_legal | tlbMsg_tlbHit & tlb_access_illegal ? offset : _GEN_232; // @[playground/src/noop/tlb.scala 131:26 140:85]
  wire [1:0] _GEN_263 = ~tlb_high_legal | tlbMsg_tlbHit & tlb_access_illegal ? level : _GEN_233; // @[playground/src/noop/tlb.scala 132:26 140:85]
  wire [63:0] _GEN_268 = ~handshake ? {{32'd0}, out_paddr_r} : _GEN_238; // @[playground/src/noop/tlb.scala 139:33 52:30]
  wire [55:0] _GEN_271 = ~handshake ? {{24'd0}, pte_addr_r} : _GEN_241; // @[playground/src/noop/tlb.scala 139:33 47:30]
  wire [4:0] _dc_mode_r_T = wpte_hs_r ? 5'h0 : 5'hb; // @[playground/src/noop/tlb.scala 175:33]
  wire [4:0] _GEN_294 = io_dcacheRW_ready ? 5'h0 : _dc_mode_r_T; // @[playground/src/noop/tlb.scala 175:27 176:40 177:31]
  wire  _GEN_295 = io_dcacheRW_ready | wpte_hs_r; // @[playground/src/noop/tlb.scala 134:28 176:40 178:31]
  wire [1:0] _GEN_296 = io_dcacheRW_rvalid ? 2'h0 : state; // @[playground/src/noop/tlb.scala 180:41 181:27 84:24]
  wire [7:0] _offset_T_1 = offset - 8'h9; // @[playground/src/noop/tlb.scala 187:39]
  wire [1:0] _level_T_1 = level - 2'h1; // @[playground/src/noop/tlb.scala 188:38]
  wire [4:0] _GEN_297 = dc_hand ? 5'h0 : dc_mode_r; // @[playground/src/noop/tlb.scala 185:30 186:31 49:30]
  wire [7:0] _GEN_298 = dc_hand ? _offset_T_1 : offset; // @[playground/src/noop/tlb.scala 131:26 185:30 187:29]
  wire [1:0] _GEN_299 = dc_hand ? _level_T_1 : level; // @[playground/src/noop/tlb.scala 132:26 185:30 188:29]
  wire [63:0] _T_73 = io_dcacheRW_rdata & 64'hf; // @[playground/src/noop/tlb.scala 191:31]
  wire [63:0] _T_77 = io_dcacheRW_rdata & 64'hd0; // @[playground/src/noop/tlb.scala 192:35]
  wire [63:0] _pte_addr_r_T_5 = pre_addr >> offset; // @[playground/src/noop/tlb.scala 196:69]
  wire [55:0] _pte_addr_r_T_7 = {io_dcacheRW_rdata[53:10],_pte_addr_r_T_5[8:0],3'h0}; // @[playground/src/noop/tlb.scala 196:46]
  wire [1:0] _GEN_300 = _T_77 != 64'h0 ? 2'h0 : state; // @[playground/src/noop/tlb.scala 192:70 193:35 84:24]
  wire  _GEN_301 = _T_77 != 64'h0 | _GEN_151; // @[playground/src/noop/tlb.scala 192:70 194:44]
  wire [55:0] _GEN_302 = _T_77 != 64'h0 ? {{24'd0}, pte_addr_r} : _pte_addr_r_T_7; // @[playground/src/noop/tlb.scala 192:70 47:30 196:40]
  wire [4:0] _GEN_303 = _T_77 != 64'h0 ? _GEN_297 : 5'h7; // @[playground/src/noop/tlb.scala 192:70 197:40]
  wire  _T_83 = out_excep_r_cause == 64'hc; // @[playground/src/noop/tlb.scala 199:133]
  wire  _T_87 = io_dcacheRW_rdata[4] ? io_mmuState_priv == 2'h1 & (~io_mmuState_mstatus[18] | out_excep_r_cause == 64'hc
    ) : io_mmuState_priv == 2'h0; // @[playground/src/noop/tlb.scala 199:35]
  wire  _T_106 = out_excep_r_cause == 64'hd & ~(io_dcacheRW_rdata[1] | io_mmuState_mstatus[19] & io_dcacheRW_rdata[3]); // @[playground/src/noop/tlb.scala 208:82]
  wire  _T_107 = _T_83 & ~io_dcacheRW_rdata[3] | _T_106; // @[playground/src/noop/tlb.scala 207:102]
  wire  _T_111 = out_excep_r_cause == 64'hf & ~io_dcacheRW_rdata[2]; // @[playground/src/noop/tlb.scala 209:79]
  wire  _T_112 = _T_107 | _T_111; // @[playground/src/noop/tlb.scala 208:152]
  wire [51:0] _ppn_mask_T_4 = 2'h0 == level ? 52'hfffffffffffff : 52'h0; // @[src/main/scala/chisel3/util/Mux.scala 81:58]
  wire [51:0] _ppn_mask_T_6 = 2'h1 == level ? 52'hffffffffffe00 : _ppn_mask_T_4; // @[src/main/scala/chisel3/util/Mux.scala 81:58]
  wire [51:0] ppn_mask = 2'h2 == level ? 52'hffffffffc0000 : _ppn_mask_T_6; // @[src/main/scala/chisel3/util/Mux.scala 81:58]
  wire [51:0] _tag_T_1 = pre_addr[63:12] & ppn_mask; // @[playground/src/noop/tlb.scala 220:78]
  wire [51:0] _GEN_304 = 4'h0 == select_r ? _tag_T_1 : tag_0; // @[playground/src/noop/tlb.scala 220:{39,39} 39:26]
  wire [51:0] _GEN_305 = 4'h1 == select_r ? _tag_T_1 : tag_1; // @[playground/src/noop/tlb.scala 220:{39,39} 39:26]
  wire [51:0] _GEN_306 = 4'h2 == select_r ? _tag_T_1 : tag_2; // @[playground/src/noop/tlb.scala 220:{39,39} 39:26]
  wire [51:0] _GEN_307 = 4'h3 == select_r ? _tag_T_1 : tag_3; // @[playground/src/noop/tlb.scala 220:{39,39} 39:26]
  wire [51:0] _GEN_308 = 4'h4 == select_r ? _tag_T_1 : tag_4; // @[playground/src/noop/tlb.scala 220:{39,39} 39:26]
  wire [51:0] _GEN_309 = 4'h5 == select_r ? _tag_T_1 : tag_5; // @[playground/src/noop/tlb.scala 220:{39,39} 39:26]
  wire [51:0] _GEN_310 = 4'h6 == select_r ? _tag_T_1 : tag_6; // @[playground/src/noop/tlb.scala 220:{39,39} 39:26]
  wire [51:0] _GEN_311 = 4'h7 == select_r ? _tag_T_1 : tag_7; // @[playground/src/noop/tlb.scala 220:{39,39} 39:26]
  wire [51:0] _GEN_312 = 4'h8 == select_r ? _tag_T_1 : tag_8; // @[playground/src/noop/tlb.scala 220:{39,39} 39:26]
  wire [51:0] _GEN_313 = 4'h9 == select_r ? _tag_T_1 : tag_9; // @[playground/src/noop/tlb.scala 220:{39,39} 39:26]
  wire [51:0] _GEN_314 = 4'ha == select_r ? _tag_T_1 : tag_10; // @[playground/src/noop/tlb.scala 220:{39,39} 39:26]
  wire [51:0] _GEN_315 = 4'hb == select_r ? _tag_T_1 : tag_11; // @[playground/src/noop/tlb.scala 220:{39,39} 39:26]
  wire [51:0] _GEN_316 = 4'hc == select_r ? _tag_T_1 : tag_12; // @[playground/src/noop/tlb.scala 220:{39,39} 39:26]
  wire [51:0] _GEN_317 = 4'hd == select_r ? _tag_T_1 : tag_13; // @[playground/src/noop/tlb.scala 220:{39,39} 39:26]
  wire [51:0] _GEN_318 = 4'he == select_r ? _tag_T_1 : tag_14; // @[playground/src/noop/tlb.scala 220:{39,39} 39:26]
  wire [51:0] _GEN_319 = 4'hf == select_r ? _tag_T_1 : tag_15; // @[playground/src/noop/tlb.scala 220:{39,39} 39:26]
  wire  _GEN_320 = 4'h0 == select_r | _GEN_130; // @[playground/src/noop/tlb.scala 221:{41,41}]
  wire  _GEN_321 = 4'h1 == select_r | _GEN_131; // @[playground/src/noop/tlb.scala 221:{41,41}]
  wire  _GEN_322 = 4'h2 == select_r | _GEN_132; // @[playground/src/noop/tlb.scala 221:{41,41}]
  wire  _GEN_323 = 4'h3 == select_r | _GEN_133; // @[playground/src/noop/tlb.scala 221:{41,41}]
  wire  _GEN_324 = 4'h4 == select_r | _GEN_134; // @[playground/src/noop/tlb.scala 221:{41,41}]
  wire  _GEN_325 = 4'h5 == select_r | _GEN_135; // @[playground/src/noop/tlb.scala 221:{41,41}]
  wire  _GEN_326 = 4'h6 == select_r | _GEN_136; // @[playground/src/noop/tlb.scala 221:{41,41}]
  wire  _GEN_327 = 4'h7 == select_r | _GEN_137; // @[playground/src/noop/tlb.scala 221:{41,41}]
  wire  _GEN_328 = 4'h8 == select_r | _GEN_138; // @[playground/src/noop/tlb.scala 221:{41,41}]
  wire  _GEN_329 = 4'h9 == select_r | _GEN_139; // @[playground/src/noop/tlb.scala 221:{41,41}]
  wire  _GEN_330 = 4'ha == select_r | _GEN_140; // @[playground/src/noop/tlb.scala 221:{41,41}]
  wire  _GEN_331 = 4'hb == select_r | _GEN_141; // @[playground/src/noop/tlb.scala 221:{41,41}]
  wire  _GEN_332 = 4'hc == select_r | _GEN_142; // @[playground/src/noop/tlb.scala 221:{41,41}]
  wire  _GEN_333 = 4'hd == select_r | _GEN_143; // @[playground/src/noop/tlb.scala 221:{41,41}]
  wire  _GEN_334 = 4'he == select_r | _GEN_144; // @[playground/src/noop/tlb.scala 221:{41,41}]
  wire  _GEN_335 = 4'hf == select_r | _GEN_145; // @[playground/src/noop/tlb.scala 221:{41,41}]
  wire [51:0] _GEN_1417 = {{32'd0}, io_dcacheRW_rdata[29:10]}; // @[playground/src/noop/tlb.scala 222:53]
  wire [51:0] update_pa = _GEN_1417 & ppn_mask; // @[playground/src/noop/tlb.scala 222:53]
  wire [19:0] _GEN_336 = 4'h0 == select_r ? update_pa[19:0] : paddr_0; // @[playground/src/noop/tlb.scala 223:{41,41} 40:26]
  wire [19:0] _GEN_337 = 4'h1 == select_r ? update_pa[19:0] : paddr_1; // @[playground/src/noop/tlb.scala 223:{41,41} 40:26]
  wire [19:0] _GEN_338 = 4'h2 == select_r ? update_pa[19:0] : paddr_2; // @[playground/src/noop/tlb.scala 223:{41,41} 40:26]
  wire [19:0] _GEN_339 = 4'h3 == select_r ? update_pa[19:0] : paddr_3; // @[playground/src/noop/tlb.scala 223:{41,41} 40:26]
  wire [19:0] _GEN_340 = 4'h4 == select_r ? update_pa[19:0] : paddr_4; // @[playground/src/noop/tlb.scala 223:{41,41} 40:26]
  wire [19:0] _GEN_341 = 4'h5 == select_r ? update_pa[19:0] : paddr_5; // @[playground/src/noop/tlb.scala 223:{41,41} 40:26]
  wire [19:0] _GEN_342 = 4'h6 == select_r ? update_pa[19:0] : paddr_6; // @[playground/src/noop/tlb.scala 223:{41,41} 40:26]
  wire [19:0] _GEN_343 = 4'h7 == select_r ? update_pa[19:0] : paddr_7; // @[playground/src/noop/tlb.scala 223:{41,41} 40:26]
  wire [19:0] _GEN_344 = 4'h8 == select_r ? update_pa[19:0] : paddr_8; // @[playground/src/noop/tlb.scala 223:{41,41} 40:26]
  wire [19:0] _GEN_345 = 4'h9 == select_r ? update_pa[19:0] : paddr_9; // @[playground/src/noop/tlb.scala 223:{41,41} 40:26]
  wire [19:0] _GEN_346 = 4'ha == select_r ? update_pa[19:0] : paddr_10; // @[playground/src/noop/tlb.scala 223:{41,41} 40:26]
  wire [19:0] _GEN_347 = 4'hb == select_r ? update_pa[19:0] : paddr_11; // @[playground/src/noop/tlb.scala 223:{41,41} 40:26]
  wire [19:0] _GEN_348 = 4'hc == select_r ? update_pa[19:0] : paddr_12; // @[playground/src/noop/tlb.scala 223:{41,41} 40:26]
  wire [19:0] _GEN_349 = 4'hd == select_r ? update_pa[19:0] : paddr_13; // @[playground/src/noop/tlb.scala 223:{41,41} 40:26]
  wire [19:0] _GEN_350 = 4'he == select_r ? update_pa[19:0] : paddr_14; // @[playground/src/noop/tlb.scala 223:{41,41} 40:26]
  wire [19:0] _GEN_351 = 4'hf == select_r ? update_pa[19:0] : paddr_15; // @[playground/src/noop/tlb.scala 223:{41,41} 40:26]
  wire [31:0] _GEN_352 = 4'h0 == select_r ? pte_addr_r : pte_addr_0; // @[playground/src/noop/tlb.scala 224:{44,44} 42:30]
  wire [31:0] _GEN_353 = 4'h1 == select_r ? pte_addr_r : pte_addr_1; // @[playground/src/noop/tlb.scala 224:{44,44} 42:30]
  wire [31:0] _GEN_354 = 4'h2 == select_r ? pte_addr_r : pte_addr_2; // @[playground/src/noop/tlb.scala 224:{44,44} 42:30]
  wire [31:0] _GEN_355 = 4'h3 == select_r ? pte_addr_r : pte_addr_3; // @[playground/src/noop/tlb.scala 224:{44,44} 42:30]
  wire [31:0] _GEN_356 = 4'h4 == select_r ? pte_addr_r : pte_addr_4; // @[playground/src/noop/tlb.scala 224:{44,44} 42:30]
  wire [31:0] _GEN_357 = 4'h5 == select_r ? pte_addr_r : pte_addr_5; // @[playground/src/noop/tlb.scala 224:{44,44} 42:30]
  wire [31:0] _GEN_358 = 4'h6 == select_r ? pte_addr_r : pte_addr_6; // @[playground/src/noop/tlb.scala 224:{44,44} 42:30]
  wire [31:0] _GEN_359 = 4'h7 == select_r ? pte_addr_r : pte_addr_7; // @[playground/src/noop/tlb.scala 224:{44,44} 42:30]
  wire [31:0] _GEN_360 = 4'h8 == select_r ? pte_addr_r : pte_addr_8; // @[playground/src/noop/tlb.scala 224:{44,44} 42:30]
  wire [31:0] _GEN_361 = 4'h9 == select_r ? pte_addr_r : pte_addr_9; // @[playground/src/noop/tlb.scala 224:{44,44} 42:30]
  wire [31:0] _GEN_362 = 4'ha == select_r ? pte_addr_r : pte_addr_10; // @[playground/src/noop/tlb.scala 224:{44,44} 42:30]
  wire [31:0] _GEN_363 = 4'hb == select_r ? pte_addr_r : pte_addr_11; // @[playground/src/noop/tlb.scala 224:{44,44} 42:30]
  wire [31:0] _GEN_364 = 4'hc == select_r ? pte_addr_r : pte_addr_12; // @[playground/src/noop/tlb.scala 224:{44,44} 42:30]
  wire [31:0] _GEN_365 = 4'hd == select_r ? pte_addr_r : pte_addr_13; // @[playground/src/noop/tlb.scala 224:{44,44} 42:30]
  wire [31:0] _GEN_366 = 4'he == select_r ? pte_addr_r : pte_addr_14; // @[playground/src/noop/tlb.scala 224:{44,44} 42:30]
  wire [31:0] _GEN_367 = 4'hf == select_r ? pte_addr_r : pte_addr_15; // @[playground/src/noop/tlb.scala 224:{44,44} 42:30]
  wire [1:0] _GEN_368 = 4'h0 == select_r ? level : pte_level_0; // @[playground/src/noop/tlb.scala 225:{45,45} 43:30]
  wire [1:0] _GEN_369 = 4'h1 == select_r ? level : pte_level_1; // @[playground/src/noop/tlb.scala 225:{45,45} 43:30]
  wire [1:0] _GEN_370 = 4'h2 == select_r ? level : pte_level_2; // @[playground/src/noop/tlb.scala 225:{45,45} 43:30]
  wire [1:0] _GEN_371 = 4'h3 == select_r ? level : pte_level_3; // @[playground/src/noop/tlb.scala 225:{45,45} 43:30]
  wire [1:0] _GEN_372 = 4'h4 == select_r ? level : pte_level_4; // @[playground/src/noop/tlb.scala 225:{45,45} 43:30]
  wire [1:0] _GEN_373 = 4'h5 == select_r ? level : pte_level_5; // @[playground/src/noop/tlb.scala 225:{45,45} 43:30]
  wire [1:0] _GEN_374 = 4'h6 == select_r ? level : pte_level_6; // @[playground/src/noop/tlb.scala 225:{45,45} 43:30]
  wire [1:0] _GEN_375 = 4'h7 == select_r ? level : pte_level_7; // @[playground/src/noop/tlb.scala 225:{45,45} 43:30]
  wire [1:0] _GEN_376 = 4'h8 == select_r ? level : pte_level_8; // @[playground/src/noop/tlb.scala 225:{45,45} 43:30]
  wire [1:0] _GEN_377 = 4'h9 == select_r ? level : pte_level_9; // @[playground/src/noop/tlb.scala 225:{45,45} 43:30]
  wire [1:0] _GEN_378 = 4'ha == select_r ? level : pte_level_10; // @[playground/src/noop/tlb.scala 225:{45,45} 43:30]
  wire [1:0] _GEN_379 = 4'hb == select_r ? level : pte_level_11; // @[playground/src/noop/tlb.scala 225:{45,45} 43:30]
  wire [1:0] _GEN_380 = 4'hc == select_r ? level : pte_level_12; // @[playground/src/noop/tlb.scala 225:{45,45} 43:30]
  wire [1:0] _GEN_381 = 4'hd == select_r ? level : pte_level_13; // @[playground/src/noop/tlb.scala 225:{45,45} 43:30]
  wire [1:0] _GEN_382 = 4'he == select_r ? level : pte_level_14; // @[playground/src/noop/tlb.scala 225:{45,45} 43:30]
  wire [1:0] _GEN_383 = 4'hf == select_r ? level : pte_level_15; // @[playground/src/noop/tlb.scala 225:{45,45} 43:30]
  wire [9:0] _GEN_384 = 4'h0 == select_r ? io_dcacheRW_rdata[9:0] : info_0; // @[playground/src/noop/tlb.scala 226:{40,40} 41:26]
  wire [9:0] _GEN_385 = 4'h1 == select_r ? io_dcacheRW_rdata[9:0] : info_1; // @[playground/src/noop/tlb.scala 226:{40,40} 41:26]
  wire [9:0] _GEN_386 = 4'h2 == select_r ? io_dcacheRW_rdata[9:0] : info_2; // @[playground/src/noop/tlb.scala 226:{40,40} 41:26]
  wire [9:0] _GEN_387 = 4'h3 == select_r ? io_dcacheRW_rdata[9:0] : info_3; // @[playground/src/noop/tlb.scala 226:{40,40} 41:26]
  wire [9:0] _GEN_388 = 4'h4 == select_r ? io_dcacheRW_rdata[9:0] : info_4; // @[playground/src/noop/tlb.scala 226:{40,40} 41:26]
  wire [9:0] _GEN_389 = 4'h5 == select_r ? io_dcacheRW_rdata[9:0] : info_5; // @[playground/src/noop/tlb.scala 226:{40,40} 41:26]
  wire [9:0] _GEN_390 = 4'h6 == select_r ? io_dcacheRW_rdata[9:0] : info_6; // @[playground/src/noop/tlb.scala 226:{40,40} 41:26]
  wire [9:0] _GEN_391 = 4'h7 == select_r ? io_dcacheRW_rdata[9:0] : info_7; // @[playground/src/noop/tlb.scala 226:{40,40} 41:26]
  wire [9:0] _GEN_392 = 4'h8 == select_r ? io_dcacheRW_rdata[9:0] : info_8; // @[playground/src/noop/tlb.scala 226:{40,40} 41:26]
  wire [9:0] _GEN_393 = 4'h9 == select_r ? io_dcacheRW_rdata[9:0] : info_9; // @[playground/src/noop/tlb.scala 226:{40,40} 41:26]
  wire [9:0] _GEN_394 = 4'ha == select_r ? io_dcacheRW_rdata[9:0] : info_10; // @[playground/src/noop/tlb.scala 226:{40,40} 41:26]
  wire [9:0] _GEN_395 = 4'hb == select_r ? io_dcacheRW_rdata[9:0] : info_11; // @[playground/src/noop/tlb.scala 226:{40,40} 41:26]
  wire [9:0] _GEN_396 = 4'hc == select_r ? io_dcacheRW_rdata[9:0] : info_12; // @[playground/src/noop/tlb.scala 226:{40,40} 41:26]
  wire [9:0] _GEN_397 = 4'hd == select_r ? io_dcacheRW_rdata[9:0] : info_13; // @[playground/src/noop/tlb.scala 226:{40,40} 41:26]
  wire [9:0] _GEN_398 = 4'he == select_r ? io_dcacheRW_rdata[9:0] : info_14; // @[playground/src/noop/tlb.scala 226:{40,40} 41:26]
  wire [9:0] _GEN_399 = 4'hf == select_r ? io_dcacheRW_rdata[9:0] : info_15; // @[playground/src/noop/tlb.scala 226:{40,40} 41:26]
  wire  _GEN_401 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     | _GEN_151; // @[playground/src/noop/tlb.scala 213:117 216:40]
  wire [51:0] _GEN_402 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? tag_0 : _GEN_304; // @[playground/src/noop/tlb.scala 213:117 39:26]
  wire [51:0] _GEN_403 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? tag_1 : _GEN_305; // @[playground/src/noop/tlb.scala 213:117 39:26]
  wire [51:0] _GEN_404 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? tag_2 : _GEN_306; // @[playground/src/noop/tlb.scala 213:117 39:26]
  wire [51:0] _GEN_405 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? tag_3 : _GEN_307; // @[playground/src/noop/tlb.scala 213:117 39:26]
  wire [51:0] _GEN_406 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? tag_4 : _GEN_308; // @[playground/src/noop/tlb.scala 213:117 39:26]
  wire [51:0] _GEN_407 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? tag_5 : _GEN_309; // @[playground/src/noop/tlb.scala 213:117 39:26]
  wire [51:0] _GEN_408 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? tag_6 : _GEN_310; // @[playground/src/noop/tlb.scala 213:117 39:26]
  wire [51:0] _GEN_409 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? tag_7 : _GEN_311; // @[playground/src/noop/tlb.scala 213:117 39:26]
  wire [51:0] _GEN_410 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? tag_8 : _GEN_312; // @[playground/src/noop/tlb.scala 213:117 39:26]
  wire [51:0] _GEN_411 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? tag_9 : _GEN_313; // @[playground/src/noop/tlb.scala 213:117 39:26]
  wire [51:0] _GEN_412 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? tag_10 : _GEN_314; // @[playground/src/noop/tlb.scala 213:117 39:26]
  wire [51:0] _GEN_413 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? tag_11 : _GEN_315; // @[playground/src/noop/tlb.scala 213:117 39:26]
  wire [51:0] _GEN_414 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? tag_12 : _GEN_316; // @[playground/src/noop/tlb.scala 213:117 39:26]
  wire [51:0] _GEN_415 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? tag_13 : _GEN_317; // @[playground/src/noop/tlb.scala 213:117 39:26]
  wire [51:0] _GEN_416 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? tag_14 : _GEN_318; // @[playground/src/noop/tlb.scala 213:117 39:26]
  wire [51:0] _GEN_417 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? tag_15 : _GEN_319; // @[playground/src/noop/tlb.scala 213:117 39:26]
  wire  _GEN_418 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? _GEN_130 : _GEN_320; // @[playground/src/noop/tlb.scala 213:117]
  wire  _GEN_419 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? _GEN_131 : _GEN_321; // @[playground/src/noop/tlb.scala 213:117]
  wire  _GEN_420 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? _GEN_132 : _GEN_322; // @[playground/src/noop/tlb.scala 213:117]
  wire  _GEN_421 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? _GEN_133 : _GEN_323; // @[playground/src/noop/tlb.scala 213:117]
  wire  _GEN_422 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? _GEN_134 : _GEN_324; // @[playground/src/noop/tlb.scala 213:117]
  wire  _GEN_423 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? _GEN_135 : _GEN_325; // @[playground/src/noop/tlb.scala 213:117]
  wire  _GEN_424 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? _GEN_136 : _GEN_326; // @[playground/src/noop/tlb.scala 213:117]
  wire  _GEN_425 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? _GEN_137 : _GEN_327; // @[playground/src/noop/tlb.scala 213:117]
  wire  _GEN_426 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? _GEN_138 : _GEN_328; // @[playground/src/noop/tlb.scala 213:117]
  wire  _GEN_427 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? _GEN_139 : _GEN_329; // @[playground/src/noop/tlb.scala 213:117]
  wire  _GEN_428 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? _GEN_140 : _GEN_330; // @[playground/src/noop/tlb.scala 213:117]
  wire  _GEN_429 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? _GEN_141 : _GEN_331; // @[playground/src/noop/tlb.scala 213:117]
  wire  _GEN_430 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? _GEN_142 : _GEN_332; // @[playground/src/noop/tlb.scala 213:117]
  wire  _GEN_431 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? _GEN_143 : _GEN_333; // @[playground/src/noop/tlb.scala 213:117]
  wire  _GEN_432 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? _GEN_144 : _GEN_334; // @[playground/src/noop/tlb.scala 213:117]
  wire  _GEN_433 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? _GEN_145 : _GEN_335; // @[playground/src/noop/tlb.scala 213:117]
  wire [19:0] _GEN_434 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? paddr_0 : _GEN_336; // @[playground/src/noop/tlb.scala 213:117 40:26]
  wire [19:0] _GEN_435 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? paddr_1 : _GEN_337; // @[playground/src/noop/tlb.scala 213:117 40:26]
  wire [19:0] _GEN_436 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? paddr_2 : _GEN_338; // @[playground/src/noop/tlb.scala 213:117 40:26]
  wire [19:0] _GEN_437 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? paddr_3 : _GEN_339; // @[playground/src/noop/tlb.scala 213:117 40:26]
  wire [19:0] _GEN_438 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? paddr_4 : _GEN_340; // @[playground/src/noop/tlb.scala 213:117 40:26]
  wire [19:0] _GEN_439 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? paddr_5 : _GEN_341; // @[playground/src/noop/tlb.scala 213:117 40:26]
  wire [19:0] _GEN_440 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? paddr_6 : _GEN_342; // @[playground/src/noop/tlb.scala 213:117 40:26]
  wire [19:0] _GEN_441 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? paddr_7 : _GEN_343; // @[playground/src/noop/tlb.scala 213:117 40:26]
  wire [19:0] _GEN_442 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? paddr_8 : _GEN_344; // @[playground/src/noop/tlb.scala 213:117 40:26]
  wire [19:0] _GEN_443 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? paddr_9 : _GEN_345; // @[playground/src/noop/tlb.scala 213:117 40:26]
  wire [19:0] _GEN_444 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? paddr_10 : _GEN_346; // @[playground/src/noop/tlb.scala 213:117 40:26]
  wire [19:0] _GEN_445 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? paddr_11 : _GEN_347; // @[playground/src/noop/tlb.scala 213:117 40:26]
  wire [19:0] _GEN_446 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? paddr_12 : _GEN_348; // @[playground/src/noop/tlb.scala 213:117 40:26]
  wire [19:0] _GEN_447 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? paddr_13 : _GEN_349; // @[playground/src/noop/tlb.scala 213:117 40:26]
  wire [19:0] _GEN_448 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? paddr_14 : _GEN_350; // @[playground/src/noop/tlb.scala 213:117 40:26]
  wire [19:0] _GEN_449 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? paddr_15 : _GEN_351; // @[playground/src/noop/tlb.scala 213:117 40:26]
  wire [31:0] _GEN_450 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? pte_addr_0 : _GEN_352; // @[playground/src/noop/tlb.scala 213:117 42:30]
  wire [31:0] _GEN_451 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? pte_addr_1 : _GEN_353; // @[playground/src/noop/tlb.scala 213:117 42:30]
  wire [31:0] _GEN_452 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? pte_addr_2 : _GEN_354; // @[playground/src/noop/tlb.scala 213:117 42:30]
  wire [31:0] _GEN_453 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? pte_addr_3 : _GEN_355; // @[playground/src/noop/tlb.scala 213:117 42:30]
  wire [31:0] _GEN_454 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? pte_addr_4 : _GEN_356; // @[playground/src/noop/tlb.scala 213:117 42:30]
  wire [31:0] _GEN_455 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? pte_addr_5 : _GEN_357; // @[playground/src/noop/tlb.scala 213:117 42:30]
  wire [31:0] _GEN_456 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? pte_addr_6 : _GEN_358; // @[playground/src/noop/tlb.scala 213:117 42:30]
  wire [31:0] _GEN_457 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? pte_addr_7 : _GEN_359; // @[playground/src/noop/tlb.scala 213:117 42:30]
  wire [31:0] _GEN_458 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? pte_addr_8 : _GEN_360; // @[playground/src/noop/tlb.scala 213:117 42:30]
  wire [31:0] _GEN_459 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? pte_addr_9 : _GEN_361; // @[playground/src/noop/tlb.scala 213:117 42:30]
  wire [31:0] _GEN_460 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? pte_addr_10 : _GEN_362; // @[playground/src/noop/tlb.scala 213:117 42:30]
  wire [31:0] _GEN_461 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? pte_addr_11 : _GEN_363; // @[playground/src/noop/tlb.scala 213:117 42:30]
  wire [31:0] _GEN_462 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? pte_addr_12 : _GEN_364; // @[playground/src/noop/tlb.scala 213:117 42:30]
  wire [31:0] _GEN_463 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? pte_addr_13 : _GEN_365; // @[playground/src/noop/tlb.scala 213:117 42:30]
  wire [31:0] _GEN_464 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? pte_addr_14 : _GEN_366; // @[playground/src/noop/tlb.scala 213:117 42:30]
  wire [31:0] _GEN_465 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? pte_addr_15 : _GEN_367; // @[playground/src/noop/tlb.scala 213:117 42:30]
  wire [1:0] _GEN_466 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? pte_level_0 : _GEN_368; // @[playground/src/noop/tlb.scala 213:117 43:30]
  wire [1:0] _GEN_467 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? pte_level_1 : _GEN_369; // @[playground/src/noop/tlb.scala 213:117 43:30]
  wire [1:0] _GEN_468 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? pte_level_2 : _GEN_370; // @[playground/src/noop/tlb.scala 213:117 43:30]
  wire [1:0] _GEN_469 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? pte_level_3 : _GEN_371; // @[playground/src/noop/tlb.scala 213:117 43:30]
  wire [1:0] _GEN_470 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? pte_level_4 : _GEN_372; // @[playground/src/noop/tlb.scala 213:117 43:30]
  wire [1:0] _GEN_471 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? pte_level_5 : _GEN_373; // @[playground/src/noop/tlb.scala 213:117 43:30]
  wire [1:0] _GEN_472 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? pte_level_6 : _GEN_374; // @[playground/src/noop/tlb.scala 213:117 43:30]
  wire [1:0] _GEN_473 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? pte_level_7 : _GEN_375; // @[playground/src/noop/tlb.scala 213:117 43:30]
  wire [1:0] _GEN_474 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? pte_level_8 : _GEN_376; // @[playground/src/noop/tlb.scala 213:117 43:30]
  wire [1:0] _GEN_475 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? pte_level_9 : _GEN_377; // @[playground/src/noop/tlb.scala 213:117 43:30]
  wire [1:0] _GEN_476 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? pte_level_10 : _GEN_378; // @[playground/src/noop/tlb.scala 213:117 43:30]
  wire [1:0] _GEN_477 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? pte_level_11 : _GEN_379; // @[playground/src/noop/tlb.scala 213:117 43:30]
  wire [1:0] _GEN_478 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? pte_level_12 : _GEN_380; // @[playground/src/noop/tlb.scala 213:117 43:30]
  wire [1:0] _GEN_479 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? pte_level_13 : _GEN_381; // @[playground/src/noop/tlb.scala 213:117 43:30]
  wire [1:0] _GEN_480 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? pte_level_14 : _GEN_382; // @[playground/src/noop/tlb.scala 213:117 43:30]
  wire [1:0] _GEN_481 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? pte_level_15 : _GEN_383; // @[playground/src/noop/tlb.scala 213:117 43:30]
  wire [9:0] _GEN_482 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? info_0 : _GEN_384; // @[playground/src/noop/tlb.scala 213:117 41:26]
  wire [9:0] _GEN_483 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? info_1 : _GEN_385; // @[playground/src/noop/tlb.scala 213:117 41:26]
  wire [9:0] _GEN_484 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? info_2 : _GEN_386; // @[playground/src/noop/tlb.scala 213:117 41:26]
  wire [9:0] _GEN_485 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? info_3 : _GEN_387; // @[playground/src/noop/tlb.scala 213:117 41:26]
  wire [9:0] _GEN_486 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? info_4 : _GEN_388; // @[playground/src/noop/tlb.scala 213:117 41:26]
  wire [9:0] _GEN_487 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? info_5 : _GEN_389; // @[playground/src/noop/tlb.scala 213:117 41:26]
  wire [9:0] _GEN_488 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? info_6 : _GEN_390; // @[playground/src/noop/tlb.scala 213:117 41:26]
  wire [9:0] _GEN_489 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? info_7 : _GEN_391; // @[playground/src/noop/tlb.scala 213:117 41:26]
  wire [9:0] _GEN_490 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? info_8 : _GEN_392; // @[playground/src/noop/tlb.scala 213:117 41:26]
  wire [9:0] _GEN_491 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? info_9 : _GEN_393; // @[playground/src/noop/tlb.scala 213:117 41:26]
  wire [9:0] _GEN_492 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? info_10 : _GEN_394; // @[playground/src/noop/tlb.scala 213:117 41:26]
  wire [9:0] _GEN_493 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? info_11 : _GEN_395; // @[playground/src/noop/tlb.scala 213:117 41:26]
  wire [9:0] _GEN_494 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? info_12 : _GEN_396; // @[playground/src/noop/tlb.scala 213:117 41:26]
  wire [9:0] _GEN_495 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? info_13 : _GEN_397; // @[playground/src/noop/tlb.scala 213:117 41:26]
  wire [9:0] _GEN_496 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? info_14 : _GEN_398; // @[playground/src/noop/tlb.scala 213:117 41:26]
  wire [9:0] _GEN_497 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? info_15 : _GEN_399; // @[playground/src/noop/tlb.scala 213:117 41:26]
  wire  _GEN_499 = _T_112 | _GEN_401; // @[playground/src/noop/tlb.scala 209:99 212:40]
  wire [51:0] _GEN_500 = _T_112 ? tag_0 : _GEN_402; // @[playground/src/noop/tlb.scala 209:99 39:26]
  wire [51:0] _GEN_501 = _T_112 ? tag_1 : _GEN_403; // @[playground/src/noop/tlb.scala 209:99 39:26]
  wire [51:0] _GEN_502 = _T_112 ? tag_2 : _GEN_404; // @[playground/src/noop/tlb.scala 209:99 39:26]
  wire [51:0] _GEN_503 = _T_112 ? tag_3 : _GEN_405; // @[playground/src/noop/tlb.scala 209:99 39:26]
  wire [51:0] _GEN_504 = _T_112 ? tag_4 : _GEN_406; // @[playground/src/noop/tlb.scala 209:99 39:26]
  wire [51:0] _GEN_505 = _T_112 ? tag_5 : _GEN_407; // @[playground/src/noop/tlb.scala 209:99 39:26]
  wire [51:0] _GEN_506 = _T_112 ? tag_6 : _GEN_408; // @[playground/src/noop/tlb.scala 209:99 39:26]
  wire [51:0] _GEN_507 = _T_112 ? tag_7 : _GEN_409; // @[playground/src/noop/tlb.scala 209:99 39:26]
  wire [51:0] _GEN_508 = _T_112 ? tag_8 : _GEN_410; // @[playground/src/noop/tlb.scala 209:99 39:26]
  wire [51:0] _GEN_509 = _T_112 ? tag_9 : _GEN_411; // @[playground/src/noop/tlb.scala 209:99 39:26]
  wire [51:0] _GEN_510 = _T_112 ? tag_10 : _GEN_412; // @[playground/src/noop/tlb.scala 209:99 39:26]
  wire [51:0] _GEN_511 = _T_112 ? tag_11 : _GEN_413; // @[playground/src/noop/tlb.scala 209:99 39:26]
  wire [51:0] _GEN_512 = _T_112 ? tag_12 : _GEN_414; // @[playground/src/noop/tlb.scala 209:99 39:26]
  wire [51:0] _GEN_513 = _T_112 ? tag_13 : _GEN_415; // @[playground/src/noop/tlb.scala 209:99 39:26]
  wire [51:0] _GEN_514 = _T_112 ? tag_14 : _GEN_416; // @[playground/src/noop/tlb.scala 209:99 39:26]
  wire [51:0] _GEN_515 = _T_112 ? tag_15 : _GEN_417; // @[playground/src/noop/tlb.scala 209:99 39:26]
  wire  _GEN_516 = _T_112 ? _GEN_130 : _GEN_418; // @[playground/src/noop/tlb.scala 209:99]
  wire  _GEN_517 = _T_112 ? _GEN_131 : _GEN_419; // @[playground/src/noop/tlb.scala 209:99]
  wire  _GEN_518 = _T_112 ? _GEN_132 : _GEN_420; // @[playground/src/noop/tlb.scala 209:99]
  wire  _GEN_519 = _T_112 ? _GEN_133 : _GEN_421; // @[playground/src/noop/tlb.scala 209:99]
  wire  _GEN_520 = _T_112 ? _GEN_134 : _GEN_422; // @[playground/src/noop/tlb.scala 209:99]
  wire  _GEN_521 = _T_112 ? _GEN_135 : _GEN_423; // @[playground/src/noop/tlb.scala 209:99]
  wire  _GEN_522 = _T_112 ? _GEN_136 : _GEN_424; // @[playground/src/noop/tlb.scala 209:99]
  wire  _GEN_523 = _T_112 ? _GEN_137 : _GEN_425; // @[playground/src/noop/tlb.scala 209:99]
  wire  _GEN_524 = _T_112 ? _GEN_138 : _GEN_426; // @[playground/src/noop/tlb.scala 209:99]
  wire  _GEN_525 = _T_112 ? _GEN_139 : _GEN_427; // @[playground/src/noop/tlb.scala 209:99]
  wire  _GEN_526 = _T_112 ? _GEN_140 : _GEN_428; // @[playground/src/noop/tlb.scala 209:99]
  wire  _GEN_527 = _T_112 ? _GEN_141 : _GEN_429; // @[playground/src/noop/tlb.scala 209:99]
  wire  _GEN_528 = _T_112 ? _GEN_142 : _GEN_430; // @[playground/src/noop/tlb.scala 209:99]
  wire  _GEN_529 = _T_112 ? _GEN_143 : _GEN_431; // @[playground/src/noop/tlb.scala 209:99]
  wire  _GEN_530 = _T_112 ? _GEN_144 : _GEN_432; // @[playground/src/noop/tlb.scala 209:99]
  wire  _GEN_531 = _T_112 ? _GEN_145 : _GEN_433; // @[playground/src/noop/tlb.scala 209:99]
  wire [19:0] _GEN_532 = _T_112 ? paddr_0 : _GEN_434; // @[playground/src/noop/tlb.scala 209:99 40:26]
  wire [19:0] _GEN_533 = _T_112 ? paddr_1 : _GEN_435; // @[playground/src/noop/tlb.scala 209:99 40:26]
  wire [19:0] _GEN_534 = _T_112 ? paddr_2 : _GEN_436; // @[playground/src/noop/tlb.scala 209:99 40:26]
  wire [19:0] _GEN_535 = _T_112 ? paddr_3 : _GEN_437; // @[playground/src/noop/tlb.scala 209:99 40:26]
  wire [19:0] _GEN_536 = _T_112 ? paddr_4 : _GEN_438; // @[playground/src/noop/tlb.scala 209:99 40:26]
  wire [19:0] _GEN_537 = _T_112 ? paddr_5 : _GEN_439; // @[playground/src/noop/tlb.scala 209:99 40:26]
  wire [19:0] _GEN_538 = _T_112 ? paddr_6 : _GEN_440; // @[playground/src/noop/tlb.scala 209:99 40:26]
  wire [19:0] _GEN_539 = _T_112 ? paddr_7 : _GEN_441; // @[playground/src/noop/tlb.scala 209:99 40:26]
  wire [19:0] _GEN_540 = _T_112 ? paddr_8 : _GEN_442; // @[playground/src/noop/tlb.scala 209:99 40:26]
  wire [19:0] _GEN_541 = _T_112 ? paddr_9 : _GEN_443; // @[playground/src/noop/tlb.scala 209:99 40:26]
  wire [19:0] _GEN_542 = _T_112 ? paddr_10 : _GEN_444; // @[playground/src/noop/tlb.scala 209:99 40:26]
  wire [19:0] _GEN_543 = _T_112 ? paddr_11 : _GEN_445; // @[playground/src/noop/tlb.scala 209:99 40:26]
  wire [19:0] _GEN_544 = _T_112 ? paddr_12 : _GEN_446; // @[playground/src/noop/tlb.scala 209:99 40:26]
  wire [19:0] _GEN_545 = _T_112 ? paddr_13 : _GEN_447; // @[playground/src/noop/tlb.scala 209:99 40:26]
  wire [19:0] _GEN_546 = _T_112 ? paddr_14 : _GEN_448; // @[playground/src/noop/tlb.scala 209:99 40:26]
  wire [19:0] _GEN_547 = _T_112 ? paddr_15 : _GEN_449; // @[playground/src/noop/tlb.scala 209:99 40:26]
  wire [31:0] _GEN_548 = _T_112 ? pte_addr_0 : _GEN_450; // @[playground/src/noop/tlb.scala 209:99 42:30]
  wire [31:0] _GEN_549 = _T_112 ? pte_addr_1 : _GEN_451; // @[playground/src/noop/tlb.scala 209:99 42:30]
  wire [31:0] _GEN_550 = _T_112 ? pte_addr_2 : _GEN_452; // @[playground/src/noop/tlb.scala 209:99 42:30]
  wire [31:0] _GEN_551 = _T_112 ? pte_addr_3 : _GEN_453; // @[playground/src/noop/tlb.scala 209:99 42:30]
  wire [31:0] _GEN_552 = _T_112 ? pte_addr_4 : _GEN_454; // @[playground/src/noop/tlb.scala 209:99 42:30]
  wire [31:0] _GEN_553 = _T_112 ? pte_addr_5 : _GEN_455; // @[playground/src/noop/tlb.scala 209:99 42:30]
  wire [31:0] _GEN_554 = _T_112 ? pte_addr_6 : _GEN_456; // @[playground/src/noop/tlb.scala 209:99 42:30]
  wire [31:0] _GEN_555 = _T_112 ? pte_addr_7 : _GEN_457; // @[playground/src/noop/tlb.scala 209:99 42:30]
  wire [31:0] _GEN_556 = _T_112 ? pte_addr_8 : _GEN_458; // @[playground/src/noop/tlb.scala 209:99 42:30]
  wire [31:0] _GEN_557 = _T_112 ? pte_addr_9 : _GEN_459; // @[playground/src/noop/tlb.scala 209:99 42:30]
  wire [31:0] _GEN_558 = _T_112 ? pte_addr_10 : _GEN_460; // @[playground/src/noop/tlb.scala 209:99 42:30]
  wire [31:0] _GEN_559 = _T_112 ? pte_addr_11 : _GEN_461; // @[playground/src/noop/tlb.scala 209:99 42:30]
  wire [31:0] _GEN_560 = _T_112 ? pte_addr_12 : _GEN_462; // @[playground/src/noop/tlb.scala 209:99 42:30]
  wire [31:0] _GEN_561 = _T_112 ? pte_addr_13 : _GEN_463; // @[playground/src/noop/tlb.scala 209:99 42:30]
  wire [31:0] _GEN_562 = _T_112 ? pte_addr_14 : _GEN_464; // @[playground/src/noop/tlb.scala 209:99 42:30]
  wire [31:0] _GEN_563 = _T_112 ? pte_addr_15 : _GEN_465; // @[playground/src/noop/tlb.scala 209:99 42:30]
  wire [1:0] _GEN_564 = _T_112 ? pte_level_0 : _GEN_466; // @[playground/src/noop/tlb.scala 209:99 43:30]
  wire [1:0] _GEN_565 = _T_112 ? pte_level_1 : _GEN_467; // @[playground/src/noop/tlb.scala 209:99 43:30]
  wire [1:0] _GEN_566 = _T_112 ? pte_level_2 : _GEN_468; // @[playground/src/noop/tlb.scala 209:99 43:30]
  wire [1:0] _GEN_567 = _T_112 ? pte_level_3 : _GEN_469; // @[playground/src/noop/tlb.scala 209:99 43:30]
  wire [1:0] _GEN_568 = _T_112 ? pte_level_4 : _GEN_470; // @[playground/src/noop/tlb.scala 209:99 43:30]
  wire [1:0] _GEN_569 = _T_112 ? pte_level_5 : _GEN_471; // @[playground/src/noop/tlb.scala 209:99 43:30]
  wire [1:0] _GEN_570 = _T_112 ? pte_level_6 : _GEN_472; // @[playground/src/noop/tlb.scala 209:99 43:30]
  wire [1:0] _GEN_571 = _T_112 ? pte_level_7 : _GEN_473; // @[playground/src/noop/tlb.scala 209:99 43:30]
  wire [1:0] _GEN_572 = _T_112 ? pte_level_8 : _GEN_474; // @[playground/src/noop/tlb.scala 209:99 43:30]
  wire [1:0] _GEN_573 = _T_112 ? pte_level_9 : _GEN_475; // @[playground/src/noop/tlb.scala 209:99 43:30]
  wire [1:0] _GEN_574 = _T_112 ? pte_level_10 : _GEN_476; // @[playground/src/noop/tlb.scala 209:99 43:30]
  wire [1:0] _GEN_575 = _T_112 ? pte_level_11 : _GEN_477; // @[playground/src/noop/tlb.scala 209:99 43:30]
  wire [1:0] _GEN_576 = _T_112 ? pte_level_12 : _GEN_478; // @[playground/src/noop/tlb.scala 209:99 43:30]
  wire [1:0] _GEN_577 = _T_112 ? pte_level_13 : _GEN_479; // @[playground/src/noop/tlb.scala 209:99 43:30]
  wire [1:0] _GEN_578 = _T_112 ? pte_level_14 : _GEN_480; // @[playground/src/noop/tlb.scala 209:99 43:30]
  wire [1:0] _GEN_579 = _T_112 ? pte_level_15 : _GEN_481; // @[playground/src/noop/tlb.scala 209:99 43:30]
  wire [9:0] _GEN_580 = _T_112 ? info_0 : _GEN_482; // @[playground/src/noop/tlb.scala 209:99 41:26]
  wire [9:0] _GEN_581 = _T_112 ? info_1 : _GEN_483; // @[playground/src/noop/tlb.scala 209:99 41:26]
  wire [9:0] _GEN_582 = _T_112 ? info_2 : _GEN_484; // @[playground/src/noop/tlb.scala 209:99 41:26]
  wire [9:0] _GEN_583 = _T_112 ? info_3 : _GEN_485; // @[playground/src/noop/tlb.scala 209:99 41:26]
  wire [9:0] _GEN_584 = _T_112 ? info_4 : _GEN_486; // @[playground/src/noop/tlb.scala 209:99 41:26]
  wire [9:0] _GEN_585 = _T_112 ? info_5 : _GEN_487; // @[playground/src/noop/tlb.scala 209:99 41:26]
  wire [9:0] _GEN_586 = _T_112 ? info_6 : _GEN_488; // @[playground/src/noop/tlb.scala 209:99 41:26]
  wire [9:0] _GEN_587 = _T_112 ? info_7 : _GEN_489; // @[playground/src/noop/tlb.scala 209:99 41:26]
  wire [9:0] _GEN_588 = _T_112 ? info_8 : _GEN_490; // @[playground/src/noop/tlb.scala 209:99 41:26]
  wire [9:0] _GEN_589 = _T_112 ? info_9 : _GEN_491; // @[playground/src/noop/tlb.scala 209:99 41:26]
  wire [9:0] _GEN_590 = _T_112 ? info_10 : _GEN_492; // @[playground/src/noop/tlb.scala 209:99 41:26]
  wire [9:0] _GEN_591 = _T_112 ? info_11 : _GEN_493; // @[playground/src/noop/tlb.scala 209:99 41:26]
  wire [9:0] _GEN_592 = _T_112 ? info_12 : _GEN_494; // @[playground/src/noop/tlb.scala 209:99 41:26]
  wire [9:0] _GEN_593 = _T_112 ? info_13 : _GEN_495; // @[playground/src/noop/tlb.scala 209:99 41:26]
  wire [9:0] _GEN_594 = _T_112 ? info_14 : _GEN_496; // @[playground/src/noop/tlb.scala 209:99 41:26]
  wire [9:0] _GEN_595 = _T_112 ? info_15 : _GEN_497; // @[playground/src/noop/tlb.scala 209:99 41:26]
  wire  _GEN_597 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] | _GEN_499; // @[playground/src/noop/tlb.scala 203:87 206:40]
  wire [51:0] _GEN_598 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? tag_0 : _GEN_500; // @[playground/src/noop/tlb.scala 203:87 39:26]
  wire [51:0] _GEN_599 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? tag_1 : _GEN_501; // @[playground/src/noop/tlb.scala 203:87 39:26]
  wire [51:0] _GEN_600 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? tag_2 : _GEN_502; // @[playground/src/noop/tlb.scala 203:87 39:26]
  wire [51:0] _GEN_601 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? tag_3 : _GEN_503; // @[playground/src/noop/tlb.scala 203:87 39:26]
  wire [51:0] _GEN_602 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? tag_4 : _GEN_504; // @[playground/src/noop/tlb.scala 203:87 39:26]
  wire [51:0] _GEN_603 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? tag_5 : _GEN_505; // @[playground/src/noop/tlb.scala 203:87 39:26]
  wire [51:0] _GEN_604 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? tag_6 : _GEN_506; // @[playground/src/noop/tlb.scala 203:87 39:26]
  wire [51:0] _GEN_605 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? tag_7 : _GEN_507; // @[playground/src/noop/tlb.scala 203:87 39:26]
  wire [51:0] _GEN_606 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? tag_8 : _GEN_508; // @[playground/src/noop/tlb.scala 203:87 39:26]
  wire [51:0] _GEN_607 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? tag_9 : _GEN_509; // @[playground/src/noop/tlb.scala 203:87 39:26]
  wire [51:0] _GEN_608 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? tag_10 : _GEN_510; // @[playground/src/noop/tlb.scala 203:87 39:26]
  wire [51:0] _GEN_609 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? tag_11 : _GEN_511; // @[playground/src/noop/tlb.scala 203:87 39:26]
  wire [51:0] _GEN_610 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? tag_12 : _GEN_512; // @[playground/src/noop/tlb.scala 203:87 39:26]
  wire [51:0] _GEN_611 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? tag_13 : _GEN_513; // @[playground/src/noop/tlb.scala 203:87 39:26]
  wire [51:0] _GEN_612 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? tag_14 : _GEN_514; // @[playground/src/noop/tlb.scala 203:87 39:26]
  wire [51:0] _GEN_613 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? tag_15 : _GEN_515; // @[playground/src/noop/tlb.scala 203:87 39:26]
  wire  _GEN_614 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? _GEN_130 : _GEN_516; // @[playground/src/noop/tlb.scala 203:87]
  wire  _GEN_615 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? _GEN_131 : _GEN_517; // @[playground/src/noop/tlb.scala 203:87]
  wire  _GEN_616 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? _GEN_132 : _GEN_518; // @[playground/src/noop/tlb.scala 203:87]
  wire  _GEN_617 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? _GEN_133 : _GEN_519; // @[playground/src/noop/tlb.scala 203:87]
  wire  _GEN_618 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? _GEN_134 : _GEN_520; // @[playground/src/noop/tlb.scala 203:87]
  wire  _GEN_619 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? _GEN_135 : _GEN_521; // @[playground/src/noop/tlb.scala 203:87]
  wire  _GEN_620 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? _GEN_136 : _GEN_522; // @[playground/src/noop/tlb.scala 203:87]
  wire  _GEN_621 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? _GEN_137 : _GEN_523; // @[playground/src/noop/tlb.scala 203:87]
  wire  _GEN_622 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? _GEN_138 : _GEN_524; // @[playground/src/noop/tlb.scala 203:87]
  wire  _GEN_623 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? _GEN_139 : _GEN_525; // @[playground/src/noop/tlb.scala 203:87]
  wire  _GEN_624 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? _GEN_140 : _GEN_526; // @[playground/src/noop/tlb.scala 203:87]
  wire  _GEN_625 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? _GEN_141 : _GEN_527; // @[playground/src/noop/tlb.scala 203:87]
  wire  _GEN_626 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? _GEN_142 : _GEN_528; // @[playground/src/noop/tlb.scala 203:87]
  wire  _GEN_627 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? _GEN_143 : _GEN_529; // @[playground/src/noop/tlb.scala 203:87]
  wire  _GEN_628 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? _GEN_144 : _GEN_530; // @[playground/src/noop/tlb.scala 203:87]
  wire  _GEN_629 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? _GEN_145 : _GEN_531; // @[playground/src/noop/tlb.scala 203:87]
  wire [19:0] _GEN_630 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? paddr_0 : _GEN_532; // @[playground/src/noop/tlb.scala 203:87 40:26]
  wire [19:0] _GEN_631 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? paddr_1 : _GEN_533; // @[playground/src/noop/tlb.scala 203:87 40:26]
  wire [19:0] _GEN_632 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? paddr_2 : _GEN_534; // @[playground/src/noop/tlb.scala 203:87 40:26]
  wire [19:0] _GEN_633 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? paddr_3 : _GEN_535; // @[playground/src/noop/tlb.scala 203:87 40:26]
  wire [19:0] _GEN_634 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? paddr_4 : _GEN_536; // @[playground/src/noop/tlb.scala 203:87 40:26]
  wire [19:0] _GEN_635 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? paddr_5 : _GEN_537; // @[playground/src/noop/tlb.scala 203:87 40:26]
  wire [19:0] _GEN_636 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? paddr_6 : _GEN_538; // @[playground/src/noop/tlb.scala 203:87 40:26]
  wire [19:0] _GEN_637 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? paddr_7 : _GEN_539; // @[playground/src/noop/tlb.scala 203:87 40:26]
  wire [19:0] _GEN_638 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? paddr_8 : _GEN_540; // @[playground/src/noop/tlb.scala 203:87 40:26]
  wire [19:0] _GEN_639 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? paddr_9 : _GEN_541; // @[playground/src/noop/tlb.scala 203:87 40:26]
  wire [19:0] _GEN_640 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? paddr_10 : _GEN_542; // @[playground/src/noop/tlb.scala 203:87 40:26]
  wire [19:0] _GEN_641 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? paddr_11 : _GEN_543; // @[playground/src/noop/tlb.scala 203:87 40:26]
  wire [19:0] _GEN_642 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? paddr_12 : _GEN_544; // @[playground/src/noop/tlb.scala 203:87 40:26]
  wire [19:0] _GEN_643 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? paddr_13 : _GEN_545; // @[playground/src/noop/tlb.scala 203:87 40:26]
  wire [19:0] _GEN_644 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? paddr_14 : _GEN_546; // @[playground/src/noop/tlb.scala 203:87 40:26]
  wire [19:0] _GEN_645 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? paddr_15 : _GEN_547; // @[playground/src/noop/tlb.scala 203:87 40:26]
  wire [31:0] _GEN_646 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? pte_addr_0 : _GEN_548; // @[playground/src/noop/tlb.scala 203:87 42:30]
  wire [31:0] _GEN_647 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? pte_addr_1 : _GEN_549; // @[playground/src/noop/tlb.scala 203:87 42:30]
  wire [31:0] _GEN_648 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? pte_addr_2 : _GEN_550; // @[playground/src/noop/tlb.scala 203:87 42:30]
  wire [31:0] _GEN_649 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? pte_addr_3 : _GEN_551; // @[playground/src/noop/tlb.scala 203:87 42:30]
  wire [31:0] _GEN_650 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? pte_addr_4 : _GEN_552; // @[playground/src/noop/tlb.scala 203:87 42:30]
  wire [31:0] _GEN_651 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? pte_addr_5 : _GEN_553; // @[playground/src/noop/tlb.scala 203:87 42:30]
  wire [31:0] _GEN_652 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? pte_addr_6 : _GEN_554; // @[playground/src/noop/tlb.scala 203:87 42:30]
  wire [31:0] _GEN_653 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? pte_addr_7 : _GEN_555; // @[playground/src/noop/tlb.scala 203:87 42:30]
  wire [31:0] _GEN_654 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? pte_addr_8 : _GEN_556; // @[playground/src/noop/tlb.scala 203:87 42:30]
  wire [31:0] _GEN_655 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? pte_addr_9 : _GEN_557; // @[playground/src/noop/tlb.scala 203:87 42:30]
  wire [31:0] _GEN_656 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? pte_addr_10 : _GEN_558; // @[playground/src/noop/tlb.scala 203:87 42:30]
  wire [31:0] _GEN_657 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? pte_addr_11 : _GEN_559; // @[playground/src/noop/tlb.scala 203:87 42:30]
  wire [31:0] _GEN_658 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? pte_addr_12 : _GEN_560; // @[playground/src/noop/tlb.scala 203:87 42:30]
  wire [31:0] _GEN_659 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? pte_addr_13 : _GEN_561; // @[playground/src/noop/tlb.scala 203:87 42:30]
  wire [31:0] _GEN_660 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? pte_addr_14 : _GEN_562; // @[playground/src/noop/tlb.scala 203:87 42:30]
  wire [31:0] _GEN_661 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? pte_addr_15 : _GEN_563; // @[playground/src/noop/tlb.scala 203:87 42:30]
  wire [1:0] _GEN_662 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? pte_level_0 : _GEN_564; // @[playground/src/noop/tlb.scala 203:87 43:30]
  wire [1:0] _GEN_663 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? pte_level_1 : _GEN_565; // @[playground/src/noop/tlb.scala 203:87 43:30]
  wire [1:0] _GEN_664 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? pte_level_2 : _GEN_566; // @[playground/src/noop/tlb.scala 203:87 43:30]
  wire [1:0] _GEN_665 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? pte_level_3 : _GEN_567; // @[playground/src/noop/tlb.scala 203:87 43:30]
  wire [1:0] _GEN_666 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? pte_level_4 : _GEN_568; // @[playground/src/noop/tlb.scala 203:87 43:30]
  wire [1:0] _GEN_667 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? pte_level_5 : _GEN_569; // @[playground/src/noop/tlb.scala 203:87 43:30]
  wire [1:0] _GEN_668 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? pte_level_6 : _GEN_570; // @[playground/src/noop/tlb.scala 203:87 43:30]
  wire [1:0] _GEN_669 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? pte_level_7 : _GEN_571; // @[playground/src/noop/tlb.scala 203:87 43:30]
  wire [1:0] _GEN_670 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? pte_level_8 : _GEN_572; // @[playground/src/noop/tlb.scala 203:87 43:30]
  wire [1:0] _GEN_671 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? pte_level_9 : _GEN_573; // @[playground/src/noop/tlb.scala 203:87 43:30]
  wire [1:0] _GEN_672 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? pte_level_10 : _GEN_574; // @[playground/src/noop/tlb.scala 203:87 43:30]
  wire [1:0] _GEN_673 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? pte_level_11 : _GEN_575; // @[playground/src/noop/tlb.scala 203:87 43:30]
  wire [1:0] _GEN_674 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? pte_level_12 : _GEN_576; // @[playground/src/noop/tlb.scala 203:87 43:30]
  wire [1:0] _GEN_675 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? pte_level_13 : _GEN_577; // @[playground/src/noop/tlb.scala 203:87 43:30]
  wire [1:0] _GEN_676 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? pte_level_14 : _GEN_578; // @[playground/src/noop/tlb.scala 203:87 43:30]
  wire [1:0] _GEN_677 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? pte_level_15 : _GEN_579; // @[playground/src/noop/tlb.scala 203:87 43:30]
  wire [9:0] _GEN_678 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? info_0 : _GEN_580; // @[playground/src/noop/tlb.scala 203:87 41:26]
  wire [9:0] _GEN_679 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? info_1 : _GEN_581; // @[playground/src/noop/tlb.scala 203:87 41:26]
  wire [9:0] _GEN_680 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? info_2 : _GEN_582; // @[playground/src/noop/tlb.scala 203:87 41:26]
  wire [9:0] _GEN_681 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? info_3 : _GEN_583; // @[playground/src/noop/tlb.scala 203:87 41:26]
  wire [9:0] _GEN_682 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? info_4 : _GEN_584; // @[playground/src/noop/tlb.scala 203:87 41:26]
  wire [9:0] _GEN_683 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? info_5 : _GEN_585; // @[playground/src/noop/tlb.scala 203:87 41:26]
  wire [9:0] _GEN_684 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? info_6 : _GEN_586; // @[playground/src/noop/tlb.scala 203:87 41:26]
  wire [9:0] _GEN_685 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? info_7 : _GEN_587; // @[playground/src/noop/tlb.scala 203:87 41:26]
  wire [9:0] _GEN_686 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? info_8 : _GEN_588; // @[playground/src/noop/tlb.scala 203:87 41:26]
  wire [9:0] _GEN_687 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? info_9 : _GEN_589; // @[playground/src/noop/tlb.scala 203:87 41:26]
  wire [9:0] _GEN_688 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? info_10 : _GEN_590; // @[playground/src/noop/tlb.scala 203:87 41:26]
  wire [9:0] _GEN_689 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? info_11 : _GEN_591; // @[playground/src/noop/tlb.scala 203:87 41:26]
  wire [9:0] _GEN_690 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? info_12 : _GEN_592; // @[playground/src/noop/tlb.scala 203:87 41:26]
  wire [9:0] _GEN_691 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? info_13 : _GEN_593; // @[playground/src/noop/tlb.scala 203:87 41:26]
  wire [9:0] _GEN_692 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? info_14 : _GEN_594; // @[playground/src/noop/tlb.scala 203:87 41:26]
  wire [9:0] _GEN_693 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? info_15 : _GEN_595; // @[playground/src/noop/tlb.scala 203:87 41:26]
  wire  _GEN_695 = _T_87 | _GEN_597; // @[playground/src/noop/tlb.scala 199:193 202:40]
  wire [51:0] _GEN_696 = _T_87 ? tag_0 : _GEN_598; // @[playground/src/noop/tlb.scala 199:193 39:26]
  wire [51:0] _GEN_697 = _T_87 ? tag_1 : _GEN_599; // @[playground/src/noop/tlb.scala 199:193 39:26]
  wire [51:0] _GEN_698 = _T_87 ? tag_2 : _GEN_600; // @[playground/src/noop/tlb.scala 199:193 39:26]
  wire [51:0] _GEN_699 = _T_87 ? tag_3 : _GEN_601; // @[playground/src/noop/tlb.scala 199:193 39:26]
  wire [51:0] _GEN_700 = _T_87 ? tag_4 : _GEN_602; // @[playground/src/noop/tlb.scala 199:193 39:26]
  wire [51:0] _GEN_701 = _T_87 ? tag_5 : _GEN_603; // @[playground/src/noop/tlb.scala 199:193 39:26]
  wire [51:0] _GEN_702 = _T_87 ? tag_6 : _GEN_604; // @[playground/src/noop/tlb.scala 199:193 39:26]
  wire [51:0] _GEN_703 = _T_87 ? tag_7 : _GEN_605; // @[playground/src/noop/tlb.scala 199:193 39:26]
  wire [51:0] _GEN_704 = _T_87 ? tag_8 : _GEN_606; // @[playground/src/noop/tlb.scala 199:193 39:26]
  wire [51:0] _GEN_705 = _T_87 ? tag_9 : _GEN_607; // @[playground/src/noop/tlb.scala 199:193 39:26]
  wire [51:0] _GEN_706 = _T_87 ? tag_10 : _GEN_608; // @[playground/src/noop/tlb.scala 199:193 39:26]
  wire [51:0] _GEN_707 = _T_87 ? tag_11 : _GEN_609; // @[playground/src/noop/tlb.scala 199:193 39:26]
  wire [51:0] _GEN_708 = _T_87 ? tag_12 : _GEN_610; // @[playground/src/noop/tlb.scala 199:193 39:26]
  wire [51:0] _GEN_709 = _T_87 ? tag_13 : _GEN_611; // @[playground/src/noop/tlb.scala 199:193 39:26]
  wire [51:0] _GEN_710 = _T_87 ? tag_14 : _GEN_612; // @[playground/src/noop/tlb.scala 199:193 39:26]
  wire [51:0] _GEN_711 = _T_87 ? tag_15 : _GEN_613; // @[playground/src/noop/tlb.scala 199:193 39:26]
  wire  _GEN_712 = _T_87 ? _GEN_130 : _GEN_614; // @[playground/src/noop/tlb.scala 199:193]
  wire  _GEN_713 = _T_87 ? _GEN_131 : _GEN_615; // @[playground/src/noop/tlb.scala 199:193]
  wire  _GEN_714 = _T_87 ? _GEN_132 : _GEN_616; // @[playground/src/noop/tlb.scala 199:193]
  wire  _GEN_715 = _T_87 ? _GEN_133 : _GEN_617; // @[playground/src/noop/tlb.scala 199:193]
  wire  _GEN_716 = _T_87 ? _GEN_134 : _GEN_618; // @[playground/src/noop/tlb.scala 199:193]
  wire  _GEN_717 = _T_87 ? _GEN_135 : _GEN_619; // @[playground/src/noop/tlb.scala 199:193]
  wire  _GEN_718 = _T_87 ? _GEN_136 : _GEN_620; // @[playground/src/noop/tlb.scala 199:193]
  wire  _GEN_719 = _T_87 ? _GEN_137 : _GEN_621; // @[playground/src/noop/tlb.scala 199:193]
  wire  _GEN_720 = _T_87 ? _GEN_138 : _GEN_622; // @[playground/src/noop/tlb.scala 199:193]
  wire  _GEN_721 = _T_87 ? _GEN_139 : _GEN_623; // @[playground/src/noop/tlb.scala 199:193]
  wire  _GEN_722 = _T_87 ? _GEN_140 : _GEN_624; // @[playground/src/noop/tlb.scala 199:193]
  wire  _GEN_723 = _T_87 ? _GEN_141 : _GEN_625; // @[playground/src/noop/tlb.scala 199:193]
  wire  _GEN_724 = _T_87 ? _GEN_142 : _GEN_626; // @[playground/src/noop/tlb.scala 199:193]
  wire  _GEN_725 = _T_87 ? _GEN_143 : _GEN_627; // @[playground/src/noop/tlb.scala 199:193]
  wire  _GEN_726 = _T_87 ? _GEN_144 : _GEN_628; // @[playground/src/noop/tlb.scala 199:193]
  wire  _GEN_727 = _T_87 ? _GEN_145 : _GEN_629; // @[playground/src/noop/tlb.scala 199:193]
  wire [19:0] _GEN_728 = _T_87 ? paddr_0 : _GEN_630; // @[playground/src/noop/tlb.scala 199:193 40:26]
  wire [19:0] _GEN_729 = _T_87 ? paddr_1 : _GEN_631; // @[playground/src/noop/tlb.scala 199:193 40:26]
  wire [19:0] _GEN_730 = _T_87 ? paddr_2 : _GEN_632; // @[playground/src/noop/tlb.scala 199:193 40:26]
  wire [19:0] _GEN_731 = _T_87 ? paddr_3 : _GEN_633; // @[playground/src/noop/tlb.scala 199:193 40:26]
  wire [19:0] _GEN_732 = _T_87 ? paddr_4 : _GEN_634; // @[playground/src/noop/tlb.scala 199:193 40:26]
  wire [19:0] _GEN_733 = _T_87 ? paddr_5 : _GEN_635; // @[playground/src/noop/tlb.scala 199:193 40:26]
  wire [19:0] _GEN_734 = _T_87 ? paddr_6 : _GEN_636; // @[playground/src/noop/tlb.scala 199:193 40:26]
  wire [19:0] _GEN_735 = _T_87 ? paddr_7 : _GEN_637; // @[playground/src/noop/tlb.scala 199:193 40:26]
  wire [19:0] _GEN_736 = _T_87 ? paddr_8 : _GEN_638; // @[playground/src/noop/tlb.scala 199:193 40:26]
  wire [19:0] _GEN_737 = _T_87 ? paddr_9 : _GEN_639; // @[playground/src/noop/tlb.scala 199:193 40:26]
  wire [19:0] _GEN_738 = _T_87 ? paddr_10 : _GEN_640; // @[playground/src/noop/tlb.scala 199:193 40:26]
  wire [19:0] _GEN_739 = _T_87 ? paddr_11 : _GEN_641; // @[playground/src/noop/tlb.scala 199:193 40:26]
  wire [19:0] _GEN_740 = _T_87 ? paddr_12 : _GEN_642; // @[playground/src/noop/tlb.scala 199:193 40:26]
  wire [19:0] _GEN_741 = _T_87 ? paddr_13 : _GEN_643; // @[playground/src/noop/tlb.scala 199:193 40:26]
  wire [19:0] _GEN_742 = _T_87 ? paddr_14 : _GEN_644; // @[playground/src/noop/tlb.scala 199:193 40:26]
  wire [19:0] _GEN_743 = _T_87 ? paddr_15 : _GEN_645; // @[playground/src/noop/tlb.scala 199:193 40:26]
  wire [31:0] _GEN_744 = _T_87 ? pte_addr_0 : _GEN_646; // @[playground/src/noop/tlb.scala 199:193 42:30]
  wire [31:0] _GEN_745 = _T_87 ? pte_addr_1 : _GEN_647; // @[playground/src/noop/tlb.scala 199:193 42:30]
  wire [31:0] _GEN_746 = _T_87 ? pte_addr_2 : _GEN_648; // @[playground/src/noop/tlb.scala 199:193 42:30]
  wire [31:0] _GEN_747 = _T_87 ? pte_addr_3 : _GEN_649; // @[playground/src/noop/tlb.scala 199:193 42:30]
  wire [31:0] _GEN_748 = _T_87 ? pte_addr_4 : _GEN_650; // @[playground/src/noop/tlb.scala 199:193 42:30]
  wire [31:0] _GEN_749 = _T_87 ? pte_addr_5 : _GEN_651; // @[playground/src/noop/tlb.scala 199:193 42:30]
  wire [31:0] _GEN_750 = _T_87 ? pte_addr_6 : _GEN_652; // @[playground/src/noop/tlb.scala 199:193 42:30]
  wire [31:0] _GEN_751 = _T_87 ? pte_addr_7 : _GEN_653; // @[playground/src/noop/tlb.scala 199:193 42:30]
  wire [31:0] _GEN_752 = _T_87 ? pte_addr_8 : _GEN_654; // @[playground/src/noop/tlb.scala 199:193 42:30]
  wire [31:0] _GEN_753 = _T_87 ? pte_addr_9 : _GEN_655; // @[playground/src/noop/tlb.scala 199:193 42:30]
  wire [31:0] _GEN_754 = _T_87 ? pte_addr_10 : _GEN_656; // @[playground/src/noop/tlb.scala 199:193 42:30]
  wire [31:0] _GEN_755 = _T_87 ? pte_addr_11 : _GEN_657; // @[playground/src/noop/tlb.scala 199:193 42:30]
  wire [31:0] _GEN_756 = _T_87 ? pte_addr_12 : _GEN_658; // @[playground/src/noop/tlb.scala 199:193 42:30]
  wire [31:0] _GEN_757 = _T_87 ? pte_addr_13 : _GEN_659; // @[playground/src/noop/tlb.scala 199:193 42:30]
  wire [31:0] _GEN_758 = _T_87 ? pte_addr_14 : _GEN_660; // @[playground/src/noop/tlb.scala 199:193 42:30]
  wire [31:0] _GEN_759 = _T_87 ? pte_addr_15 : _GEN_661; // @[playground/src/noop/tlb.scala 199:193 42:30]
  wire [1:0] _GEN_760 = _T_87 ? pte_level_0 : _GEN_662; // @[playground/src/noop/tlb.scala 199:193 43:30]
  wire [1:0] _GEN_761 = _T_87 ? pte_level_1 : _GEN_663; // @[playground/src/noop/tlb.scala 199:193 43:30]
  wire [1:0] _GEN_762 = _T_87 ? pte_level_2 : _GEN_664; // @[playground/src/noop/tlb.scala 199:193 43:30]
  wire [1:0] _GEN_763 = _T_87 ? pte_level_3 : _GEN_665; // @[playground/src/noop/tlb.scala 199:193 43:30]
  wire [1:0] _GEN_764 = _T_87 ? pte_level_4 : _GEN_666; // @[playground/src/noop/tlb.scala 199:193 43:30]
  wire [1:0] _GEN_765 = _T_87 ? pte_level_5 : _GEN_667; // @[playground/src/noop/tlb.scala 199:193 43:30]
  wire [1:0] _GEN_766 = _T_87 ? pte_level_6 : _GEN_668; // @[playground/src/noop/tlb.scala 199:193 43:30]
  wire [1:0] _GEN_767 = _T_87 ? pte_level_7 : _GEN_669; // @[playground/src/noop/tlb.scala 199:193 43:30]
  wire [1:0] _GEN_768 = _T_87 ? pte_level_8 : _GEN_670; // @[playground/src/noop/tlb.scala 199:193 43:30]
  wire [1:0] _GEN_769 = _T_87 ? pte_level_9 : _GEN_671; // @[playground/src/noop/tlb.scala 199:193 43:30]
  wire [1:0] _GEN_770 = _T_87 ? pte_level_10 : _GEN_672; // @[playground/src/noop/tlb.scala 199:193 43:30]
  wire [1:0] _GEN_771 = _T_87 ? pte_level_11 : _GEN_673; // @[playground/src/noop/tlb.scala 199:193 43:30]
  wire [1:0] _GEN_772 = _T_87 ? pte_level_12 : _GEN_674; // @[playground/src/noop/tlb.scala 199:193 43:30]
  wire [1:0] _GEN_773 = _T_87 ? pte_level_13 : _GEN_675; // @[playground/src/noop/tlb.scala 199:193 43:30]
  wire [1:0] _GEN_774 = _T_87 ? pte_level_14 : _GEN_676; // @[playground/src/noop/tlb.scala 199:193 43:30]
  wire [1:0] _GEN_775 = _T_87 ? pte_level_15 : _GEN_677; // @[playground/src/noop/tlb.scala 199:193 43:30]
  wire [9:0] _GEN_776 = _T_87 ? info_0 : _GEN_678; // @[playground/src/noop/tlb.scala 199:193 41:26]
  wire [9:0] _GEN_777 = _T_87 ? info_1 : _GEN_679; // @[playground/src/noop/tlb.scala 199:193 41:26]
  wire [9:0] _GEN_778 = _T_87 ? info_2 : _GEN_680; // @[playground/src/noop/tlb.scala 199:193 41:26]
  wire [9:0] _GEN_779 = _T_87 ? info_3 : _GEN_681; // @[playground/src/noop/tlb.scala 199:193 41:26]
  wire [9:0] _GEN_780 = _T_87 ? info_4 : _GEN_682; // @[playground/src/noop/tlb.scala 199:193 41:26]
  wire [9:0] _GEN_781 = _T_87 ? info_5 : _GEN_683; // @[playground/src/noop/tlb.scala 199:193 41:26]
  wire [9:0] _GEN_782 = _T_87 ? info_6 : _GEN_684; // @[playground/src/noop/tlb.scala 199:193 41:26]
  wire [9:0] _GEN_783 = _T_87 ? info_7 : _GEN_685; // @[playground/src/noop/tlb.scala 199:193 41:26]
  wire [9:0] _GEN_784 = _T_87 ? info_8 : _GEN_686; // @[playground/src/noop/tlb.scala 199:193 41:26]
  wire [9:0] _GEN_785 = _T_87 ? info_9 : _GEN_687; // @[playground/src/noop/tlb.scala 199:193 41:26]
  wire [9:0] _GEN_786 = _T_87 ? info_10 : _GEN_688; // @[playground/src/noop/tlb.scala 199:193 41:26]
  wire [9:0] _GEN_787 = _T_87 ? info_11 : _GEN_689; // @[playground/src/noop/tlb.scala 199:193 41:26]
  wire [9:0] _GEN_788 = _T_87 ? info_12 : _GEN_690; // @[playground/src/noop/tlb.scala 199:193 41:26]
  wire [9:0] _GEN_789 = _T_87 ? info_13 : _GEN_691; // @[playground/src/noop/tlb.scala 199:193 41:26]
  wire [9:0] _GEN_790 = _T_87 ? info_14 : _GEN_692; // @[playground/src/noop/tlb.scala 199:193 41:26]
  wire [9:0] _GEN_791 = _T_87 ? info_15 : _GEN_693; // @[playground/src/noop/tlb.scala 199:193 41:26]
  wire [1:0] _GEN_792 = _T_73 == 64'h1 ? _GEN_300 : 2'h0; // @[playground/src/noop/tlb.scala 191:76]
  wire  _GEN_793 = _T_73 == 64'h1 ? _GEN_301 : _GEN_695; // @[playground/src/noop/tlb.scala 191:76]
  wire [55:0] _GEN_794 = _T_73 == 64'h1 ? _GEN_302 : {{24'd0}, pte_addr_r}; // @[playground/src/noop/tlb.scala 191:76 47:30]
  wire [4:0] _GEN_795 = _T_73 == 64'h1 ? _GEN_303 : _GEN_297; // @[playground/src/noop/tlb.scala 191:76]
  wire [51:0] _GEN_796 = _T_73 == 64'h1 ? tag_0 : _GEN_696; // @[playground/src/noop/tlb.scala 191:76 39:26]
  wire [51:0] _GEN_797 = _T_73 == 64'h1 ? tag_1 : _GEN_697; // @[playground/src/noop/tlb.scala 191:76 39:26]
  wire [51:0] _GEN_798 = _T_73 == 64'h1 ? tag_2 : _GEN_698; // @[playground/src/noop/tlb.scala 191:76 39:26]
  wire [51:0] _GEN_799 = _T_73 == 64'h1 ? tag_3 : _GEN_699; // @[playground/src/noop/tlb.scala 191:76 39:26]
  wire [51:0] _GEN_800 = _T_73 == 64'h1 ? tag_4 : _GEN_700; // @[playground/src/noop/tlb.scala 191:76 39:26]
  wire [51:0] _GEN_801 = _T_73 == 64'h1 ? tag_5 : _GEN_701; // @[playground/src/noop/tlb.scala 191:76 39:26]
  wire [51:0] _GEN_802 = _T_73 == 64'h1 ? tag_6 : _GEN_702; // @[playground/src/noop/tlb.scala 191:76 39:26]
  wire [51:0] _GEN_803 = _T_73 == 64'h1 ? tag_7 : _GEN_703; // @[playground/src/noop/tlb.scala 191:76 39:26]
  wire [51:0] _GEN_804 = _T_73 == 64'h1 ? tag_8 : _GEN_704; // @[playground/src/noop/tlb.scala 191:76 39:26]
  wire [51:0] _GEN_805 = _T_73 == 64'h1 ? tag_9 : _GEN_705; // @[playground/src/noop/tlb.scala 191:76 39:26]
  wire [51:0] _GEN_806 = _T_73 == 64'h1 ? tag_10 : _GEN_706; // @[playground/src/noop/tlb.scala 191:76 39:26]
  wire [51:0] _GEN_807 = _T_73 == 64'h1 ? tag_11 : _GEN_707; // @[playground/src/noop/tlb.scala 191:76 39:26]
  wire [51:0] _GEN_808 = _T_73 == 64'h1 ? tag_12 : _GEN_708; // @[playground/src/noop/tlb.scala 191:76 39:26]
  wire [51:0] _GEN_809 = _T_73 == 64'h1 ? tag_13 : _GEN_709; // @[playground/src/noop/tlb.scala 191:76 39:26]
  wire [51:0] _GEN_810 = _T_73 == 64'h1 ? tag_14 : _GEN_710; // @[playground/src/noop/tlb.scala 191:76 39:26]
  wire [51:0] _GEN_811 = _T_73 == 64'h1 ? tag_15 : _GEN_711; // @[playground/src/noop/tlb.scala 191:76 39:26]
  wire  _GEN_812 = _T_73 == 64'h1 ? _GEN_130 : _GEN_712; // @[playground/src/noop/tlb.scala 191:76]
  wire  _GEN_813 = _T_73 == 64'h1 ? _GEN_131 : _GEN_713; // @[playground/src/noop/tlb.scala 191:76]
  wire  _GEN_814 = _T_73 == 64'h1 ? _GEN_132 : _GEN_714; // @[playground/src/noop/tlb.scala 191:76]
  wire  _GEN_815 = _T_73 == 64'h1 ? _GEN_133 : _GEN_715; // @[playground/src/noop/tlb.scala 191:76]
  wire  _GEN_816 = _T_73 == 64'h1 ? _GEN_134 : _GEN_716; // @[playground/src/noop/tlb.scala 191:76]
  wire  _GEN_817 = _T_73 == 64'h1 ? _GEN_135 : _GEN_717; // @[playground/src/noop/tlb.scala 191:76]
  wire  _GEN_818 = _T_73 == 64'h1 ? _GEN_136 : _GEN_718; // @[playground/src/noop/tlb.scala 191:76]
  wire  _GEN_819 = _T_73 == 64'h1 ? _GEN_137 : _GEN_719; // @[playground/src/noop/tlb.scala 191:76]
  wire  _GEN_820 = _T_73 == 64'h1 ? _GEN_138 : _GEN_720; // @[playground/src/noop/tlb.scala 191:76]
  wire  _GEN_821 = _T_73 == 64'h1 ? _GEN_139 : _GEN_721; // @[playground/src/noop/tlb.scala 191:76]
  wire  _GEN_822 = _T_73 == 64'h1 ? _GEN_140 : _GEN_722; // @[playground/src/noop/tlb.scala 191:76]
  wire  _GEN_823 = _T_73 == 64'h1 ? _GEN_141 : _GEN_723; // @[playground/src/noop/tlb.scala 191:76]
  wire  _GEN_824 = _T_73 == 64'h1 ? _GEN_142 : _GEN_724; // @[playground/src/noop/tlb.scala 191:76]
  wire  _GEN_825 = _T_73 == 64'h1 ? _GEN_143 : _GEN_725; // @[playground/src/noop/tlb.scala 191:76]
  wire  _GEN_826 = _T_73 == 64'h1 ? _GEN_144 : _GEN_726; // @[playground/src/noop/tlb.scala 191:76]
  wire  _GEN_827 = _T_73 == 64'h1 ? _GEN_145 : _GEN_727; // @[playground/src/noop/tlb.scala 191:76]
  wire [19:0] _GEN_828 = _T_73 == 64'h1 ? paddr_0 : _GEN_728; // @[playground/src/noop/tlb.scala 191:76 40:26]
  wire [19:0] _GEN_829 = _T_73 == 64'h1 ? paddr_1 : _GEN_729; // @[playground/src/noop/tlb.scala 191:76 40:26]
  wire [19:0] _GEN_830 = _T_73 == 64'h1 ? paddr_2 : _GEN_730; // @[playground/src/noop/tlb.scala 191:76 40:26]
  wire [19:0] _GEN_831 = _T_73 == 64'h1 ? paddr_3 : _GEN_731; // @[playground/src/noop/tlb.scala 191:76 40:26]
  wire [19:0] _GEN_832 = _T_73 == 64'h1 ? paddr_4 : _GEN_732; // @[playground/src/noop/tlb.scala 191:76 40:26]
  wire [19:0] _GEN_833 = _T_73 == 64'h1 ? paddr_5 : _GEN_733; // @[playground/src/noop/tlb.scala 191:76 40:26]
  wire [19:0] _GEN_834 = _T_73 == 64'h1 ? paddr_6 : _GEN_734; // @[playground/src/noop/tlb.scala 191:76 40:26]
  wire [19:0] _GEN_835 = _T_73 == 64'h1 ? paddr_7 : _GEN_735; // @[playground/src/noop/tlb.scala 191:76 40:26]
  wire [19:0] _GEN_836 = _T_73 == 64'h1 ? paddr_8 : _GEN_736; // @[playground/src/noop/tlb.scala 191:76 40:26]
  wire [19:0] _GEN_837 = _T_73 == 64'h1 ? paddr_9 : _GEN_737; // @[playground/src/noop/tlb.scala 191:76 40:26]
  wire [19:0] _GEN_838 = _T_73 == 64'h1 ? paddr_10 : _GEN_738; // @[playground/src/noop/tlb.scala 191:76 40:26]
  wire [19:0] _GEN_839 = _T_73 == 64'h1 ? paddr_11 : _GEN_739; // @[playground/src/noop/tlb.scala 191:76 40:26]
  wire [19:0] _GEN_840 = _T_73 == 64'h1 ? paddr_12 : _GEN_740; // @[playground/src/noop/tlb.scala 191:76 40:26]
  wire [19:0] _GEN_841 = _T_73 == 64'h1 ? paddr_13 : _GEN_741; // @[playground/src/noop/tlb.scala 191:76 40:26]
  wire [19:0] _GEN_842 = _T_73 == 64'h1 ? paddr_14 : _GEN_742; // @[playground/src/noop/tlb.scala 191:76 40:26]
  wire [19:0] _GEN_843 = _T_73 == 64'h1 ? paddr_15 : _GEN_743; // @[playground/src/noop/tlb.scala 191:76 40:26]
  wire [31:0] _GEN_844 = _T_73 == 64'h1 ? pte_addr_0 : _GEN_744; // @[playground/src/noop/tlb.scala 191:76 42:30]
  wire [31:0] _GEN_845 = _T_73 == 64'h1 ? pte_addr_1 : _GEN_745; // @[playground/src/noop/tlb.scala 191:76 42:30]
  wire [31:0] _GEN_846 = _T_73 == 64'h1 ? pte_addr_2 : _GEN_746; // @[playground/src/noop/tlb.scala 191:76 42:30]
  wire [31:0] _GEN_847 = _T_73 == 64'h1 ? pte_addr_3 : _GEN_747; // @[playground/src/noop/tlb.scala 191:76 42:30]
  wire [31:0] _GEN_848 = _T_73 == 64'h1 ? pte_addr_4 : _GEN_748; // @[playground/src/noop/tlb.scala 191:76 42:30]
  wire [31:0] _GEN_849 = _T_73 == 64'h1 ? pte_addr_5 : _GEN_749; // @[playground/src/noop/tlb.scala 191:76 42:30]
  wire [31:0] _GEN_850 = _T_73 == 64'h1 ? pte_addr_6 : _GEN_750; // @[playground/src/noop/tlb.scala 191:76 42:30]
  wire [31:0] _GEN_851 = _T_73 == 64'h1 ? pte_addr_7 : _GEN_751; // @[playground/src/noop/tlb.scala 191:76 42:30]
  wire [31:0] _GEN_852 = _T_73 == 64'h1 ? pte_addr_8 : _GEN_752; // @[playground/src/noop/tlb.scala 191:76 42:30]
  wire [31:0] _GEN_853 = _T_73 == 64'h1 ? pte_addr_9 : _GEN_753; // @[playground/src/noop/tlb.scala 191:76 42:30]
  wire [31:0] _GEN_854 = _T_73 == 64'h1 ? pte_addr_10 : _GEN_754; // @[playground/src/noop/tlb.scala 191:76 42:30]
  wire [31:0] _GEN_855 = _T_73 == 64'h1 ? pte_addr_11 : _GEN_755; // @[playground/src/noop/tlb.scala 191:76 42:30]
  wire [31:0] _GEN_856 = _T_73 == 64'h1 ? pte_addr_12 : _GEN_756; // @[playground/src/noop/tlb.scala 191:76 42:30]
  wire [31:0] _GEN_857 = _T_73 == 64'h1 ? pte_addr_13 : _GEN_757; // @[playground/src/noop/tlb.scala 191:76 42:30]
  wire [31:0] _GEN_858 = _T_73 == 64'h1 ? pte_addr_14 : _GEN_758; // @[playground/src/noop/tlb.scala 191:76 42:30]
  wire [31:0] _GEN_859 = _T_73 == 64'h1 ? pte_addr_15 : _GEN_759; // @[playground/src/noop/tlb.scala 191:76 42:30]
  wire [1:0] _GEN_860 = _T_73 == 64'h1 ? pte_level_0 : _GEN_760; // @[playground/src/noop/tlb.scala 191:76 43:30]
  wire [1:0] _GEN_861 = _T_73 == 64'h1 ? pte_level_1 : _GEN_761; // @[playground/src/noop/tlb.scala 191:76 43:30]
  wire [1:0] _GEN_862 = _T_73 == 64'h1 ? pte_level_2 : _GEN_762; // @[playground/src/noop/tlb.scala 191:76 43:30]
  wire [1:0] _GEN_863 = _T_73 == 64'h1 ? pte_level_3 : _GEN_763; // @[playground/src/noop/tlb.scala 191:76 43:30]
  wire [1:0] _GEN_864 = _T_73 == 64'h1 ? pte_level_4 : _GEN_764; // @[playground/src/noop/tlb.scala 191:76 43:30]
  wire [1:0] _GEN_865 = _T_73 == 64'h1 ? pte_level_5 : _GEN_765; // @[playground/src/noop/tlb.scala 191:76 43:30]
  wire [1:0] _GEN_866 = _T_73 == 64'h1 ? pte_level_6 : _GEN_766; // @[playground/src/noop/tlb.scala 191:76 43:30]
  wire [1:0] _GEN_867 = _T_73 == 64'h1 ? pte_level_7 : _GEN_767; // @[playground/src/noop/tlb.scala 191:76 43:30]
  wire [1:0] _GEN_868 = _T_73 == 64'h1 ? pte_level_8 : _GEN_768; // @[playground/src/noop/tlb.scala 191:76 43:30]
  wire [1:0] _GEN_869 = _T_73 == 64'h1 ? pte_level_9 : _GEN_769; // @[playground/src/noop/tlb.scala 191:76 43:30]
  wire [1:0] _GEN_870 = _T_73 == 64'h1 ? pte_level_10 : _GEN_770; // @[playground/src/noop/tlb.scala 191:76 43:30]
  wire [1:0] _GEN_871 = _T_73 == 64'h1 ? pte_level_11 : _GEN_771; // @[playground/src/noop/tlb.scala 191:76 43:30]
  wire [1:0] _GEN_872 = _T_73 == 64'h1 ? pte_level_12 : _GEN_772; // @[playground/src/noop/tlb.scala 191:76 43:30]
  wire [1:0] _GEN_873 = _T_73 == 64'h1 ? pte_level_13 : _GEN_773; // @[playground/src/noop/tlb.scala 191:76 43:30]
  wire [1:0] _GEN_874 = _T_73 == 64'h1 ? pte_level_14 : _GEN_774; // @[playground/src/noop/tlb.scala 191:76 43:30]
  wire [1:0] _GEN_875 = _T_73 == 64'h1 ? pte_level_15 : _GEN_775; // @[playground/src/noop/tlb.scala 191:76 43:30]
  wire [9:0] _GEN_876 = _T_73 == 64'h1 ? info_0 : _GEN_776; // @[playground/src/noop/tlb.scala 191:76 41:26]
  wire [9:0] _GEN_877 = _T_73 == 64'h1 ? info_1 : _GEN_777; // @[playground/src/noop/tlb.scala 191:76 41:26]
  wire [9:0] _GEN_878 = _T_73 == 64'h1 ? info_2 : _GEN_778; // @[playground/src/noop/tlb.scala 191:76 41:26]
  wire [9:0] _GEN_879 = _T_73 == 64'h1 ? info_3 : _GEN_779; // @[playground/src/noop/tlb.scala 191:76 41:26]
  wire [9:0] _GEN_880 = _T_73 == 64'h1 ? info_4 : _GEN_780; // @[playground/src/noop/tlb.scala 191:76 41:26]
  wire [9:0] _GEN_881 = _T_73 == 64'h1 ? info_5 : _GEN_781; // @[playground/src/noop/tlb.scala 191:76 41:26]
  wire [9:0] _GEN_882 = _T_73 == 64'h1 ? info_6 : _GEN_782; // @[playground/src/noop/tlb.scala 191:76 41:26]
  wire [9:0] _GEN_883 = _T_73 == 64'h1 ? info_7 : _GEN_783; // @[playground/src/noop/tlb.scala 191:76 41:26]
  wire [9:0] _GEN_884 = _T_73 == 64'h1 ? info_8 : _GEN_784; // @[playground/src/noop/tlb.scala 191:76 41:26]
  wire [9:0] _GEN_885 = _T_73 == 64'h1 ? info_9 : _GEN_785; // @[playground/src/noop/tlb.scala 191:76 41:26]
  wire [9:0] _GEN_886 = _T_73 == 64'h1 ? info_10 : _GEN_786; // @[playground/src/noop/tlb.scala 191:76 41:26]
  wire [9:0] _GEN_887 = _T_73 == 64'h1 ? info_11 : _GEN_787; // @[playground/src/noop/tlb.scala 191:76 41:26]
  wire [9:0] _GEN_888 = _T_73 == 64'h1 ? info_12 : _GEN_788; // @[playground/src/noop/tlb.scala 191:76 41:26]
  wire [9:0] _GEN_889 = _T_73 == 64'h1 ? info_13 : _GEN_789; // @[playground/src/noop/tlb.scala 191:76 41:26]
  wire [9:0] _GEN_890 = _T_73 == 64'h1 ? info_14 : _GEN_790; // @[playground/src/noop/tlb.scala 191:76 41:26]
  wire [9:0] _GEN_891 = _T_73 == 64'h1 ? info_15 : _GEN_791; // @[playground/src/noop/tlb.scala 191:76 41:26]
  wire [1:0] _GEN_892 = io_dcacheRW_rvalid ? _GEN_792 : state; // @[playground/src/noop/tlb.scala 190:41 84:24]
  wire  _GEN_893 = io_dcacheRW_rvalid ? _GEN_793 : _GEN_151; // @[playground/src/noop/tlb.scala 190:41]
  wire [55:0] _GEN_894 = io_dcacheRW_rvalid ? _GEN_794 : {{24'd0}, pte_addr_r}; // @[playground/src/noop/tlb.scala 190:41 47:30]
  wire [4:0] _GEN_895 = io_dcacheRW_rvalid ? _GEN_795 : _GEN_297; // @[playground/src/noop/tlb.scala 190:41]
  wire [51:0] _GEN_896 = io_dcacheRW_rvalid ? _GEN_796 : tag_0; // @[playground/src/noop/tlb.scala 190:41 39:26]
  wire [51:0] _GEN_897 = io_dcacheRW_rvalid ? _GEN_797 : tag_1; // @[playground/src/noop/tlb.scala 190:41 39:26]
  wire [51:0] _GEN_898 = io_dcacheRW_rvalid ? _GEN_798 : tag_2; // @[playground/src/noop/tlb.scala 190:41 39:26]
  wire [51:0] _GEN_899 = io_dcacheRW_rvalid ? _GEN_799 : tag_3; // @[playground/src/noop/tlb.scala 190:41 39:26]
  wire [51:0] _GEN_900 = io_dcacheRW_rvalid ? _GEN_800 : tag_4; // @[playground/src/noop/tlb.scala 190:41 39:26]
  wire [51:0] _GEN_901 = io_dcacheRW_rvalid ? _GEN_801 : tag_5; // @[playground/src/noop/tlb.scala 190:41 39:26]
  wire [51:0] _GEN_902 = io_dcacheRW_rvalid ? _GEN_802 : tag_6; // @[playground/src/noop/tlb.scala 190:41 39:26]
  wire [51:0] _GEN_903 = io_dcacheRW_rvalid ? _GEN_803 : tag_7; // @[playground/src/noop/tlb.scala 190:41 39:26]
  wire [51:0] _GEN_904 = io_dcacheRW_rvalid ? _GEN_804 : tag_8; // @[playground/src/noop/tlb.scala 190:41 39:26]
  wire [51:0] _GEN_905 = io_dcacheRW_rvalid ? _GEN_805 : tag_9; // @[playground/src/noop/tlb.scala 190:41 39:26]
  wire [51:0] _GEN_906 = io_dcacheRW_rvalid ? _GEN_806 : tag_10; // @[playground/src/noop/tlb.scala 190:41 39:26]
  wire [51:0] _GEN_907 = io_dcacheRW_rvalid ? _GEN_807 : tag_11; // @[playground/src/noop/tlb.scala 190:41 39:26]
  wire [51:0] _GEN_908 = io_dcacheRW_rvalid ? _GEN_808 : tag_12; // @[playground/src/noop/tlb.scala 190:41 39:26]
  wire [51:0] _GEN_909 = io_dcacheRW_rvalid ? _GEN_809 : tag_13; // @[playground/src/noop/tlb.scala 190:41 39:26]
  wire [51:0] _GEN_910 = io_dcacheRW_rvalid ? _GEN_810 : tag_14; // @[playground/src/noop/tlb.scala 190:41 39:26]
  wire [51:0] _GEN_911 = io_dcacheRW_rvalid ? _GEN_811 : tag_15; // @[playground/src/noop/tlb.scala 190:41 39:26]
  wire  _GEN_912 = io_dcacheRW_rvalid ? _GEN_812 : _GEN_130; // @[playground/src/noop/tlb.scala 190:41]
  wire  _GEN_913 = io_dcacheRW_rvalid ? _GEN_813 : _GEN_131; // @[playground/src/noop/tlb.scala 190:41]
  wire  _GEN_914 = io_dcacheRW_rvalid ? _GEN_814 : _GEN_132; // @[playground/src/noop/tlb.scala 190:41]
  wire  _GEN_915 = io_dcacheRW_rvalid ? _GEN_815 : _GEN_133; // @[playground/src/noop/tlb.scala 190:41]
  wire  _GEN_916 = io_dcacheRW_rvalid ? _GEN_816 : _GEN_134; // @[playground/src/noop/tlb.scala 190:41]
  wire  _GEN_917 = io_dcacheRW_rvalid ? _GEN_817 : _GEN_135; // @[playground/src/noop/tlb.scala 190:41]
  wire  _GEN_918 = io_dcacheRW_rvalid ? _GEN_818 : _GEN_136; // @[playground/src/noop/tlb.scala 190:41]
  wire  _GEN_919 = io_dcacheRW_rvalid ? _GEN_819 : _GEN_137; // @[playground/src/noop/tlb.scala 190:41]
  wire  _GEN_920 = io_dcacheRW_rvalid ? _GEN_820 : _GEN_138; // @[playground/src/noop/tlb.scala 190:41]
  wire  _GEN_921 = io_dcacheRW_rvalid ? _GEN_821 : _GEN_139; // @[playground/src/noop/tlb.scala 190:41]
  wire  _GEN_922 = io_dcacheRW_rvalid ? _GEN_822 : _GEN_140; // @[playground/src/noop/tlb.scala 190:41]
  wire  _GEN_923 = io_dcacheRW_rvalid ? _GEN_823 : _GEN_141; // @[playground/src/noop/tlb.scala 190:41]
  wire  _GEN_924 = io_dcacheRW_rvalid ? _GEN_824 : _GEN_142; // @[playground/src/noop/tlb.scala 190:41]
  wire  _GEN_925 = io_dcacheRW_rvalid ? _GEN_825 : _GEN_143; // @[playground/src/noop/tlb.scala 190:41]
  wire  _GEN_926 = io_dcacheRW_rvalid ? _GEN_826 : _GEN_144; // @[playground/src/noop/tlb.scala 190:41]
  wire  _GEN_927 = io_dcacheRW_rvalid ? _GEN_827 : _GEN_145; // @[playground/src/noop/tlb.scala 190:41]
  wire [19:0] _GEN_928 = io_dcacheRW_rvalid ? _GEN_828 : paddr_0; // @[playground/src/noop/tlb.scala 190:41 40:26]
  wire [19:0] _GEN_929 = io_dcacheRW_rvalid ? _GEN_829 : paddr_1; // @[playground/src/noop/tlb.scala 190:41 40:26]
  wire [19:0] _GEN_930 = io_dcacheRW_rvalid ? _GEN_830 : paddr_2; // @[playground/src/noop/tlb.scala 190:41 40:26]
  wire [19:0] _GEN_931 = io_dcacheRW_rvalid ? _GEN_831 : paddr_3; // @[playground/src/noop/tlb.scala 190:41 40:26]
  wire [19:0] _GEN_932 = io_dcacheRW_rvalid ? _GEN_832 : paddr_4; // @[playground/src/noop/tlb.scala 190:41 40:26]
  wire [19:0] _GEN_933 = io_dcacheRW_rvalid ? _GEN_833 : paddr_5; // @[playground/src/noop/tlb.scala 190:41 40:26]
  wire [19:0] _GEN_934 = io_dcacheRW_rvalid ? _GEN_834 : paddr_6; // @[playground/src/noop/tlb.scala 190:41 40:26]
  wire [19:0] _GEN_935 = io_dcacheRW_rvalid ? _GEN_835 : paddr_7; // @[playground/src/noop/tlb.scala 190:41 40:26]
  wire [19:0] _GEN_936 = io_dcacheRW_rvalid ? _GEN_836 : paddr_8; // @[playground/src/noop/tlb.scala 190:41 40:26]
  wire [19:0] _GEN_937 = io_dcacheRW_rvalid ? _GEN_837 : paddr_9; // @[playground/src/noop/tlb.scala 190:41 40:26]
  wire [19:0] _GEN_938 = io_dcacheRW_rvalid ? _GEN_838 : paddr_10; // @[playground/src/noop/tlb.scala 190:41 40:26]
  wire [19:0] _GEN_939 = io_dcacheRW_rvalid ? _GEN_839 : paddr_11; // @[playground/src/noop/tlb.scala 190:41 40:26]
  wire [19:0] _GEN_940 = io_dcacheRW_rvalid ? _GEN_840 : paddr_12; // @[playground/src/noop/tlb.scala 190:41 40:26]
  wire [19:0] _GEN_941 = io_dcacheRW_rvalid ? _GEN_841 : paddr_13; // @[playground/src/noop/tlb.scala 190:41 40:26]
  wire [19:0] _GEN_942 = io_dcacheRW_rvalid ? _GEN_842 : paddr_14; // @[playground/src/noop/tlb.scala 190:41 40:26]
  wire [19:0] _GEN_943 = io_dcacheRW_rvalid ? _GEN_843 : paddr_15; // @[playground/src/noop/tlb.scala 190:41 40:26]
  wire [31:0] _GEN_944 = io_dcacheRW_rvalid ? _GEN_844 : pte_addr_0; // @[playground/src/noop/tlb.scala 190:41 42:30]
  wire [31:0] _GEN_945 = io_dcacheRW_rvalid ? _GEN_845 : pte_addr_1; // @[playground/src/noop/tlb.scala 190:41 42:30]
  wire [31:0] _GEN_946 = io_dcacheRW_rvalid ? _GEN_846 : pte_addr_2; // @[playground/src/noop/tlb.scala 190:41 42:30]
  wire [31:0] _GEN_947 = io_dcacheRW_rvalid ? _GEN_847 : pte_addr_3; // @[playground/src/noop/tlb.scala 190:41 42:30]
  wire [31:0] _GEN_948 = io_dcacheRW_rvalid ? _GEN_848 : pte_addr_4; // @[playground/src/noop/tlb.scala 190:41 42:30]
  wire [31:0] _GEN_949 = io_dcacheRW_rvalid ? _GEN_849 : pte_addr_5; // @[playground/src/noop/tlb.scala 190:41 42:30]
  wire [31:0] _GEN_950 = io_dcacheRW_rvalid ? _GEN_850 : pte_addr_6; // @[playground/src/noop/tlb.scala 190:41 42:30]
  wire [31:0] _GEN_951 = io_dcacheRW_rvalid ? _GEN_851 : pte_addr_7; // @[playground/src/noop/tlb.scala 190:41 42:30]
  wire [31:0] _GEN_952 = io_dcacheRW_rvalid ? _GEN_852 : pte_addr_8; // @[playground/src/noop/tlb.scala 190:41 42:30]
  wire [31:0] _GEN_953 = io_dcacheRW_rvalid ? _GEN_853 : pte_addr_9; // @[playground/src/noop/tlb.scala 190:41 42:30]
  wire [31:0] _GEN_954 = io_dcacheRW_rvalid ? _GEN_854 : pte_addr_10; // @[playground/src/noop/tlb.scala 190:41 42:30]
  wire [31:0] _GEN_955 = io_dcacheRW_rvalid ? _GEN_855 : pte_addr_11; // @[playground/src/noop/tlb.scala 190:41 42:30]
  wire [31:0] _GEN_956 = io_dcacheRW_rvalid ? _GEN_856 : pte_addr_12; // @[playground/src/noop/tlb.scala 190:41 42:30]
  wire [31:0] _GEN_957 = io_dcacheRW_rvalid ? _GEN_857 : pte_addr_13; // @[playground/src/noop/tlb.scala 190:41 42:30]
  wire [31:0] _GEN_958 = io_dcacheRW_rvalid ? _GEN_858 : pte_addr_14; // @[playground/src/noop/tlb.scala 190:41 42:30]
  wire [31:0] _GEN_959 = io_dcacheRW_rvalid ? _GEN_859 : pte_addr_15; // @[playground/src/noop/tlb.scala 190:41 42:30]
  wire [1:0] _GEN_960 = io_dcacheRW_rvalid ? _GEN_860 : pte_level_0; // @[playground/src/noop/tlb.scala 190:41 43:30]
  wire [1:0] _GEN_961 = io_dcacheRW_rvalid ? _GEN_861 : pte_level_1; // @[playground/src/noop/tlb.scala 190:41 43:30]
  wire [1:0] _GEN_962 = io_dcacheRW_rvalid ? _GEN_862 : pte_level_2; // @[playground/src/noop/tlb.scala 190:41 43:30]
  wire [1:0] _GEN_963 = io_dcacheRW_rvalid ? _GEN_863 : pte_level_3; // @[playground/src/noop/tlb.scala 190:41 43:30]
  wire [1:0] _GEN_964 = io_dcacheRW_rvalid ? _GEN_864 : pte_level_4; // @[playground/src/noop/tlb.scala 190:41 43:30]
  wire [1:0] _GEN_965 = io_dcacheRW_rvalid ? _GEN_865 : pte_level_5; // @[playground/src/noop/tlb.scala 190:41 43:30]
  wire [1:0] _GEN_966 = io_dcacheRW_rvalid ? _GEN_866 : pte_level_6; // @[playground/src/noop/tlb.scala 190:41 43:30]
  wire [1:0] _GEN_967 = io_dcacheRW_rvalid ? _GEN_867 : pte_level_7; // @[playground/src/noop/tlb.scala 190:41 43:30]
  wire [1:0] _GEN_968 = io_dcacheRW_rvalid ? _GEN_868 : pte_level_8; // @[playground/src/noop/tlb.scala 190:41 43:30]
  wire [1:0] _GEN_969 = io_dcacheRW_rvalid ? _GEN_869 : pte_level_9; // @[playground/src/noop/tlb.scala 190:41 43:30]
  wire [1:0] _GEN_970 = io_dcacheRW_rvalid ? _GEN_870 : pte_level_10; // @[playground/src/noop/tlb.scala 190:41 43:30]
  wire [1:0] _GEN_971 = io_dcacheRW_rvalid ? _GEN_871 : pte_level_11; // @[playground/src/noop/tlb.scala 190:41 43:30]
  wire [1:0] _GEN_972 = io_dcacheRW_rvalid ? _GEN_872 : pte_level_12; // @[playground/src/noop/tlb.scala 190:41 43:30]
  wire [1:0] _GEN_973 = io_dcacheRW_rvalid ? _GEN_873 : pte_level_13; // @[playground/src/noop/tlb.scala 190:41 43:30]
  wire [1:0] _GEN_974 = io_dcacheRW_rvalid ? _GEN_874 : pte_level_14; // @[playground/src/noop/tlb.scala 190:41 43:30]
  wire [1:0] _GEN_975 = io_dcacheRW_rvalid ? _GEN_875 : pte_level_15; // @[playground/src/noop/tlb.scala 190:41 43:30]
  wire [9:0] _GEN_976 = io_dcacheRW_rvalid ? _GEN_876 : info_0; // @[playground/src/noop/tlb.scala 190:41 41:26]
  wire [9:0] _GEN_977 = io_dcacheRW_rvalid ? _GEN_877 : info_1; // @[playground/src/noop/tlb.scala 190:41 41:26]
  wire [9:0] _GEN_978 = io_dcacheRW_rvalid ? _GEN_878 : info_2; // @[playground/src/noop/tlb.scala 190:41 41:26]
  wire [9:0] _GEN_979 = io_dcacheRW_rvalid ? _GEN_879 : info_3; // @[playground/src/noop/tlb.scala 190:41 41:26]
  wire [9:0] _GEN_980 = io_dcacheRW_rvalid ? _GEN_880 : info_4; // @[playground/src/noop/tlb.scala 190:41 41:26]
  wire [9:0] _GEN_981 = io_dcacheRW_rvalid ? _GEN_881 : info_5; // @[playground/src/noop/tlb.scala 190:41 41:26]
  wire [9:0] _GEN_982 = io_dcacheRW_rvalid ? _GEN_882 : info_6; // @[playground/src/noop/tlb.scala 190:41 41:26]
  wire [9:0] _GEN_983 = io_dcacheRW_rvalid ? _GEN_883 : info_7; // @[playground/src/noop/tlb.scala 190:41 41:26]
  wire [9:0] _GEN_984 = io_dcacheRW_rvalid ? _GEN_884 : info_8; // @[playground/src/noop/tlb.scala 190:41 41:26]
  wire [9:0] _GEN_985 = io_dcacheRW_rvalid ? _GEN_885 : info_9; // @[playground/src/noop/tlb.scala 190:41 41:26]
  wire [9:0] _GEN_986 = io_dcacheRW_rvalid ? _GEN_886 : info_10; // @[playground/src/noop/tlb.scala 190:41 41:26]
  wire [9:0] _GEN_987 = io_dcacheRW_rvalid ? _GEN_887 : info_11; // @[playground/src/noop/tlb.scala 190:41 41:26]
  wire [9:0] _GEN_988 = io_dcacheRW_rvalid ? _GEN_888 : info_12; // @[playground/src/noop/tlb.scala 190:41 41:26]
  wire [9:0] _GEN_989 = io_dcacheRW_rvalid ? _GEN_889 : info_13; // @[playground/src/noop/tlb.scala 190:41 41:26]
  wire [9:0] _GEN_990 = io_dcacheRW_rvalid ? _GEN_890 : info_14; // @[playground/src/noop/tlb.scala 190:41 41:26]
  wire [9:0] _GEN_991 = io_dcacheRW_rvalid ? _GEN_891 : info_15; // @[playground/src/noop/tlb.scala 190:41 41:26]
  wire [4:0] _GEN_992 = 2'h1 == state ? _GEN_895 : dc_mode_r; // @[playground/src/noop/tlb.scala 136:22 49:30]
  wire [7:0] _GEN_993 = 2'h1 == state ? _GEN_298 : offset; // @[playground/src/noop/tlb.scala 136:22 131:26]
  wire [1:0] _GEN_994 = 2'h1 == state ? _GEN_299 : level; // @[playground/src/noop/tlb.scala 136:22 132:26]
  wire [1:0] _GEN_995 = 2'h1 == state ? _GEN_892 : state; // @[playground/src/noop/tlb.scala 136:22 84:24]
  wire  _GEN_996 = 2'h1 == state ? _GEN_893 : _GEN_151; // @[playground/src/noop/tlb.scala 136:22]
  wire [55:0] _GEN_997 = 2'h1 == state ? _GEN_894 : {{24'd0}, pte_addr_r}; // @[playground/src/noop/tlb.scala 136:22 47:30]
  wire [51:0] _GEN_998 = 2'h1 == state ? _GEN_896 : tag_0; // @[playground/src/noop/tlb.scala 136:22 39:26]
  wire [51:0] _GEN_999 = 2'h1 == state ? _GEN_897 : tag_1; // @[playground/src/noop/tlb.scala 136:22 39:26]
  wire [51:0] _GEN_1000 = 2'h1 == state ? _GEN_898 : tag_2; // @[playground/src/noop/tlb.scala 136:22 39:26]
  wire [51:0] _GEN_1001 = 2'h1 == state ? _GEN_899 : tag_3; // @[playground/src/noop/tlb.scala 136:22 39:26]
  wire [51:0] _GEN_1002 = 2'h1 == state ? _GEN_900 : tag_4; // @[playground/src/noop/tlb.scala 136:22 39:26]
  wire [51:0] _GEN_1003 = 2'h1 == state ? _GEN_901 : tag_5; // @[playground/src/noop/tlb.scala 136:22 39:26]
  wire [51:0] _GEN_1004 = 2'h1 == state ? _GEN_902 : tag_6; // @[playground/src/noop/tlb.scala 136:22 39:26]
  wire [51:0] _GEN_1005 = 2'h1 == state ? _GEN_903 : tag_7; // @[playground/src/noop/tlb.scala 136:22 39:26]
  wire [51:0] _GEN_1006 = 2'h1 == state ? _GEN_904 : tag_8; // @[playground/src/noop/tlb.scala 136:22 39:26]
  wire [51:0] _GEN_1007 = 2'h1 == state ? _GEN_905 : tag_9; // @[playground/src/noop/tlb.scala 136:22 39:26]
  wire [51:0] _GEN_1008 = 2'h1 == state ? _GEN_906 : tag_10; // @[playground/src/noop/tlb.scala 136:22 39:26]
  wire [51:0] _GEN_1009 = 2'h1 == state ? _GEN_907 : tag_11; // @[playground/src/noop/tlb.scala 136:22 39:26]
  wire [51:0] _GEN_1010 = 2'h1 == state ? _GEN_908 : tag_12; // @[playground/src/noop/tlb.scala 136:22 39:26]
  wire [51:0] _GEN_1011 = 2'h1 == state ? _GEN_909 : tag_13; // @[playground/src/noop/tlb.scala 136:22 39:26]
  wire [51:0] _GEN_1012 = 2'h1 == state ? _GEN_910 : tag_14; // @[playground/src/noop/tlb.scala 136:22 39:26]
  wire [51:0] _GEN_1013 = 2'h1 == state ? _GEN_911 : tag_15; // @[playground/src/noop/tlb.scala 136:22 39:26]
  wire  _GEN_1014 = 2'h1 == state ? _GEN_912 : _GEN_130; // @[playground/src/noop/tlb.scala 136:22]
  wire  _GEN_1015 = 2'h1 == state ? _GEN_913 : _GEN_131; // @[playground/src/noop/tlb.scala 136:22]
  wire  _GEN_1016 = 2'h1 == state ? _GEN_914 : _GEN_132; // @[playground/src/noop/tlb.scala 136:22]
  wire  _GEN_1017 = 2'h1 == state ? _GEN_915 : _GEN_133; // @[playground/src/noop/tlb.scala 136:22]
  wire  _GEN_1018 = 2'h1 == state ? _GEN_916 : _GEN_134; // @[playground/src/noop/tlb.scala 136:22]
  wire  _GEN_1019 = 2'h1 == state ? _GEN_917 : _GEN_135; // @[playground/src/noop/tlb.scala 136:22]
  wire  _GEN_1020 = 2'h1 == state ? _GEN_918 : _GEN_136; // @[playground/src/noop/tlb.scala 136:22]
  wire  _GEN_1021 = 2'h1 == state ? _GEN_919 : _GEN_137; // @[playground/src/noop/tlb.scala 136:22]
  wire  _GEN_1022 = 2'h1 == state ? _GEN_920 : _GEN_138; // @[playground/src/noop/tlb.scala 136:22]
  wire  _GEN_1023 = 2'h1 == state ? _GEN_921 : _GEN_139; // @[playground/src/noop/tlb.scala 136:22]
  wire  _GEN_1024 = 2'h1 == state ? _GEN_922 : _GEN_140; // @[playground/src/noop/tlb.scala 136:22]
  wire  _GEN_1025 = 2'h1 == state ? _GEN_923 : _GEN_141; // @[playground/src/noop/tlb.scala 136:22]
  wire  _GEN_1026 = 2'h1 == state ? _GEN_924 : _GEN_142; // @[playground/src/noop/tlb.scala 136:22]
  wire  _GEN_1027 = 2'h1 == state ? _GEN_925 : _GEN_143; // @[playground/src/noop/tlb.scala 136:22]
  wire  _GEN_1028 = 2'h1 == state ? _GEN_926 : _GEN_144; // @[playground/src/noop/tlb.scala 136:22]
  wire  _GEN_1029 = 2'h1 == state ? _GEN_927 : _GEN_145; // @[playground/src/noop/tlb.scala 136:22]
  wire [19:0] _GEN_1030 = 2'h1 == state ? _GEN_928 : paddr_0; // @[playground/src/noop/tlb.scala 136:22 40:26]
  wire [19:0] _GEN_1031 = 2'h1 == state ? _GEN_929 : paddr_1; // @[playground/src/noop/tlb.scala 136:22 40:26]
  wire [19:0] _GEN_1032 = 2'h1 == state ? _GEN_930 : paddr_2; // @[playground/src/noop/tlb.scala 136:22 40:26]
  wire [19:0] _GEN_1033 = 2'h1 == state ? _GEN_931 : paddr_3; // @[playground/src/noop/tlb.scala 136:22 40:26]
  wire [19:0] _GEN_1034 = 2'h1 == state ? _GEN_932 : paddr_4; // @[playground/src/noop/tlb.scala 136:22 40:26]
  wire [19:0] _GEN_1035 = 2'h1 == state ? _GEN_933 : paddr_5; // @[playground/src/noop/tlb.scala 136:22 40:26]
  wire [19:0] _GEN_1036 = 2'h1 == state ? _GEN_934 : paddr_6; // @[playground/src/noop/tlb.scala 136:22 40:26]
  wire [19:0] _GEN_1037 = 2'h1 == state ? _GEN_935 : paddr_7; // @[playground/src/noop/tlb.scala 136:22 40:26]
  wire [19:0] _GEN_1038 = 2'h1 == state ? _GEN_936 : paddr_8; // @[playground/src/noop/tlb.scala 136:22 40:26]
  wire [19:0] _GEN_1039 = 2'h1 == state ? _GEN_937 : paddr_9; // @[playground/src/noop/tlb.scala 136:22 40:26]
  wire [19:0] _GEN_1040 = 2'h1 == state ? _GEN_938 : paddr_10; // @[playground/src/noop/tlb.scala 136:22 40:26]
  wire [19:0] _GEN_1041 = 2'h1 == state ? _GEN_939 : paddr_11; // @[playground/src/noop/tlb.scala 136:22 40:26]
  wire [19:0] _GEN_1042 = 2'h1 == state ? _GEN_940 : paddr_12; // @[playground/src/noop/tlb.scala 136:22 40:26]
  wire [19:0] _GEN_1043 = 2'h1 == state ? _GEN_941 : paddr_13; // @[playground/src/noop/tlb.scala 136:22 40:26]
  wire [19:0] _GEN_1044 = 2'h1 == state ? _GEN_942 : paddr_14; // @[playground/src/noop/tlb.scala 136:22 40:26]
  wire [19:0] _GEN_1045 = 2'h1 == state ? _GEN_943 : paddr_15; // @[playground/src/noop/tlb.scala 136:22 40:26]
  wire [31:0] _GEN_1046 = 2'h1 == state ? _GEN_944 : pte_addr_0; // @[playground/src/noop/tlb.scala 136:22 42:30]
  wire [31:0] _GEN_1047 = 2'h1 == state ? _GEN_945 : pte_addr_1; // @[playground/src/noop/tlb.scala 136:22 42:30]
  wire [31:0] _GEN_1048 = 2'h1 == state ? _GEN_946 : pte_addr_2; // @[playground/src/noop/tlb.scala 136:22 42:30]
  wire [31:0] _GEN_1049 = 2'h1 == state ? _GEN_947 : pte_addr_3; // @[playground/src/noop/tlb.scala 136:22 42:30]
  wire [31:0] _GEN_1050 = 2'h1 == state ? _GEN_948 : pte_addr_4; // @[playground/src/noop/tlb.scala 136:22 42:30]
  wire [31:0] _GEN_1051 = 2'h1 == state ? _GEN_949 : pte_addr_5; // @[playground/src/noop/tlb.scala 136:22 42:30]
  wire [31:0] _GEN_1052 = 2'h1 == state ? _GEN_950 : pte_addr_6; // @[playground/src/noop/tlb.scala 136:22 42:30]
  wire [31:0] _GEN_1053 = 2'h1 == state ? _GEN_951 : pte_addr_7; // @[playground/src/noop/tlb.scala 136:22 42:30]
  wire [31:0] _GEN_1054 = 2'h1 == state ? _GEN_952 : pte_addr_8; // @[playground/src/noop/tlb.scala 136:22 42:30]
  wire [31:0] _GEN_1055 = 2'h1 == state ? _GEN_953 : pte_addr_9; // @[playground/src/noop/tlb.scala 136:22 42:30]
  wire [31:0] _GEN_1056 = 2'h1 == state ? _GEN_954 : pte_addr_10; // @[playground/src/noop/tlb.scala 136:22 42:30]
  wire [31:0] _GEN_1057 = 2'h1 == state ? _GEN_955 : pte_addr_11; // @[playground/src/noop/tlb.scala 136:22 42:30]
  wire [31:0] _GEN_1058 = 2'h1 == state ? _GEN_956 : pte_addr_12; // @[playground/src/noop/tlb.scala 136:22 42:30]
  wire [31:0] _GEN_1059 = 2'h1 == state ? _GEN_957 : pte_addr_13; // @[playground/src/noop/tlb.scala 136:22 42:30]
  wire [31:0] _GEN_1060 = 2'h1 == state ? _GEN_958 : pte_addr_14; // @[playground/src/noop/tlb.scala 136:22 42:30]
  wire [31:0] _GEN_1061 = 2'h1 == state ? _GEN_959 : pte_addr_15; // @[playground/src/noop/tlb.scala 136:22 42:30]
  wire [1:0] _GEN_1062 = 2'h1 == state ? _GEN_960 : pte_level_0; // @[playground/src/noop/tlb.scala 136:22 43:30]
  wire [1:0] _GEN_1063 = 2'h1 == state ? _GEN_961 : pte_level_1; // @[playground/src/noop/tlb.scala 136:22 43:30]
  wire [1:0] _GEN_1064 = 2'h1 == state ? _GEN_962 : pte_level_2; // @[playground/src/noop/tlb.scala 136:22 43:30]
  wire [1:0] _GEN_1065 = 2'h1 == state ? _GEN_963 : pte_level_3; // @[playground/src/noop/tlb.scala 136:22 43:30]
  wire [1:0] _GEN_1066 = 2'h1 == state ? _GEN_964 : pte_level_4; // @[playground/src/noop/tlb.scala 136:22 43:30]
  wire [1:0] _GEN_1067 = 2'h1 == state ? _GEN_965 : pte_level_5; // @[playground/src/noop/tlb.scala 136:22 43:30]
  wire [1:0] _GEN_1068 = 2'h1 == state ? _GEN_966 : pte_level_6; // @[playground/src/noop/tlb.scala 136:22 43:30]
  wire [1:0] _GEN_1069 = 2'h1 == state ? _GEN_967 : pte_level_7; // @[playground/src/noop/tlb.scala 136:22 43:30]
  wire [1:0] _GEN_1070 = 2'h1 == state ? _GEN_968 : pte_level_8; // @[playground/src/noop/tlb.scala 136:22 43:30]
  wire [1:0] _GEN_1071 = 2'h1 == state ? _GEN_969 : pte_level_9; // @[playground/src/noop/tlb.scala 136:22 43:30]
  wire [1:0] _GEN_1072 = 2'h1 == state ? _GEN_970 : pte_level_10; // @[playground/src/noop/tlb.scala 136:22 43:30]
  wire [1:0] _GEN_1073 = 2'h1 == state ? _GEN_971 : pte_level_11; // @[playground/src/noop/tlb.scala 136:22 43:30]
  wire [1:0] _GEN_1074 = 2'h1 == state ? _GEN_972 : pte_level_12; // @[playground/src/noop/tlb.scala 136:22 43:30]
  wire [1:0] _GEN_1075 = 2'h1 == state ? _GEN_973 : pte_level_13; // @[playground/src/noop/tlb.scala 136:22 43:30]
  wire [1:0] _GEN_1076 = 2'h1 == state ? _GEN_974 : pte_level_14; // @[playground/src/noop/tlb.scala 136:22 43:30]
  wire [1:0] _GEN_1077 = 2'h1 == state ? _GEN_975 : pte_level_15; // @[playground/src/noop/tlb.scala 136:22 43:30]
  wire [9:0] _GEN_1078 = 2'h1 == state ? _GEN_976 : info_0; // @[playground/src/noop/tlb.scala 136:22 41:26]
  wire [9:0] _GEN_1079 = 2'h1 == state ? _GEN_977 : info_1; // @[playground/src/noop/tlb.scala 136:22 41:26]
  wire [9:0] _GEN_1080 = 2'h1 == state ? _GEN_978 : info_2; // @[playground/src/noop/tlb.scala 136:22 41:26]
  wire [9:0] _GEN_1081 = 2'h1 == state ? _GEN_979 : info_3; // @[playground/src/noop/tlb.scala 136:22 41:26]
  wire [9:0] _GEN_1082 = 2'h1 == state ? _GEN_980 : info_4; // @[playground/src/noop/tlb.scala 136:22 41:26]
  wire [9:0] _GEN_1083 = 2'h1 == state ? _GEN_981 : info_5; // @[playground/src/noop/tlb.scala 136:22 41:26]
  wire [9:0] _GEN_1084 = 2'h1 == state ? _GEN_982 : info_6; // @[playground/src/noop/tlb.scala 136:22 41:26]
  wire [9:0] _GEN_1085 = 2'h1 == state ? _GEN_983 : info_7; // @[playground/src/noop/tlb.scala 136:22 41:26]
  wire [9:0] _GEN_1086 = 2'h1 == state ? _GEN_984 : info_8; // @[playground/src/noop/tlb.scala 136:22 41:26]
  wire [9:0] _GEN_1087 = 2'h1 == state ? _GEN_985 : info_9; // @[playground/src/noop/tlb.scala 136:22 41:26]
  wire [9:0] _GEN_1088 = 2'h1 == state ? _GEN_986 : info_10; // @[playground/src/noop/tlb.scala 136:22 41:26]
  wire [9:0] _GEN_1089 = 2'h1 == state ? _GEN_987 : info_11; // @[playground/src/noop/tlb.scala 136:22 41:26]
  wire [9:0] _GEN_1090 = 2'h1 == state ? _GEN_988 : info_12; // @[playground/src/noop/tlb.scala 136:22 41:26]
  wire [9:0] _GEN_1091 = 2'h1 == state ? _GEN_989 : info_13; // @[playground/src/noop/tlb.scala 136:22 41:26]
  wire [9:0] _GEN_1092 = 2'h1 == state ? _GEN_990 : info_14; // @[playground/src/noop/tlb.scala 136:22 41:26]
  wire [9:0] _GEN_1093 = 2'h1 == state ? _GEN_991 : info_15; // @[playground/src/noop/tlb.scala 136:22 41:26]
  wire [55:0] _GEN_1100 = 2'h3 == state ? {{24'd0}, pte_addr_r} : _GEN_997; // @[playground/src/noop/tlb.scala 136:22 47:30]
  wire [63:0] _GEN_1202 = 2'h0 == state ? _GEN_268 : {{32'd0}, out_paddr_r}; // @[playground/src/noop/tlb.scala 136:22 52:30]
  wire [55:0] _GEN_1205 = 2'h0 == state ? _GEN_271 : _GEN_1100; // @[playground/src/noop/tlb.scala 136:22]
  wire [63:0] _GEN_1312 = is_Sv39 | state != 2'h0 ? _GEN_1202 : io_va2pa_vaddr; // @[playground/src/noop/tlb.scala 135:37 233:21]
  wire [55:0] _GEN_1315 = is_Sv39 | state != 2'h0 ? _GEN_1205 : {{24'd0}, pte_addr_r}; // @[playground/src/noop/tlb.scala 135:37 47:30]
  wire [55:0] _GEN_1418 = reset ? 56'h0 : _GEN_1315; // @[playground/src/noop/tlb.scala 47:{30,30}]
  wire [63:0] _GEN_1419 = reset ? 64'h0 : _GEN_1312; // @[playground/src/noop/tlb.scala 52:{30,30}]
  MaxPeriodFibonacciLFSR_2 select_prng ( // @[src/main/scala/chisel3/util/random/PRNG.scala 91:22]
    .clock(select_prng_clock),
    .reset(select_prng_reset),
    .io_out_0(select_prng_io_out_0),
    .io_out_1(select_prng_io_out_1),
    .io_out_2(select_prng_io_out_2),
    .io_out_3(select_prng_io_out_3)
  );
  assign io_va2pa_ready = io_va2pa_vvalid & _T_50 & ~io_flush & ~flush_r; // @[playground/src/noop/tlb.scala 98:74]
  assign io_va2pa_paddr = out_paddr_r; // @[playground/src/noop/tlb.scala 113:20]
  assign io_va2pa_pvalid = out_valid_r; // @[playground/src/noop/tlb.scala 114:21]
  assign io_va2pa_tlb_excep_cause = out_excep_r_cause; // @[playground/src/noop/tlb.scala 115:24]
  assign io_va2pa_tlb_excep_tval = out_excep_r_tval; // @[playground/src/noop/tlb.scala 115:24]
  assign io_va2pa_tlb_excep_en = out_excep_r_en; // @[playground/src/noop/tlb.scala 115:24]
  assign io_dcacheRW_addr = pte_addr_r; // @[playground/src/noop/tlb.scala 117:22]
  assign io_dcacheRW_wdata = wpte_data_r; // @[playground/src/noop/tlb.scala 118:23]
  assign io_dcacheRW_dc_mode = dc_mode_r; // @[playground/src/noop/tlb.scala 119:25]
  assign select_prng_clock = clock;
  assign select_prng_reset = reset;
  always @(posedge clock) begin
    if (reset) begin // @[playground/src/noop/tlb.scala 39:26]
      tag_0 <= 52'h0; // @[playground/src/noop/tlb.scala 39:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (!(2'h0 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
        if (!(2'h3 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
          tag_0 <= _GEN_998;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 39:26]
      tag_1 <= 52'h0; // @[playground/src/noop/tlb.scala 39:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (!(2'h0 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
        if (!(2'h3 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
          tag_1 <= _GEN_999;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 39:26]
      tag_2 <= 52'h0; // @[playground/src/noop/tlb.scala 39:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (!(2'h0 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
        if (!(2'h3 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
          tag_2 <= _GEN_1000;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 39:26]
      tag_3 <= 52'h0; // @[playground/src/noop/tlb.scala 39:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (!(2'h0 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
        if (!(2'h3 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
          tag_3 <= _GEN_1001;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 39:26]
      tag_4 <= 52'h0; // @[playground/src/noop/tlb.scala 39:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (!(2'h0 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
        if (!(2'h3 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
          tag_4 <= _GEN_1002;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 39:26]
      tag_5 <= 52'h0; // @[playground/src/noop/tlb.scala 39:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (!(2'h0 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
        if (!(2'h3 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
          tag_5 <= _GEN_1003;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 39:26]
      tag_6 <= 52'h0; // @[playground/src/noop/tlb.scala 39:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (!(2'h0 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
        if (!(2'h3 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
          tag_6 <= _GEN_1004;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 39:26]
      tag_7 <= 52'h0; // @[playground/src/noop/tlb.scala 39:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (!(2'h0 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
        if (!(2'h3 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
          tag_7 <= _GEN_1005;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 39:26]
      tag_8 <= 52'h0; // @[playground/src/noop/tlb.scala 39:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (!(2'h0 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
        if (!(2'h3 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
          tag_8 <= _GEN_1006;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 39:26]
      tag_9 <= 52'h0; // @[playground/src/noop/tlb.scala 39:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (!(2'h0 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
        if (!(2'h3 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
          tag_9 <= _GEN_1007;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 39:26]
      tag_10 <= 52'h0; // @[playground/src/noop/tlb.scala 39:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (!(2'h0 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
        if (!(2'h3 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
          tag_10 <= _GEN_1008;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 39:26]
      tag_11 <= 52'h0; // @[playground/src/noop/tlb.scala 39:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (!(2'h0 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
        if (!(2'h3 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
          tag_11 <= _GEN_1009;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 39:26]
      tag_12 <= 52'h0; // @[playground/src/noop/tlb.scala 39:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (!(2'h0 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
        if (!(2'h3 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
          tag_12 <= _GEN_1010;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 39:26]
      tag_13 <= 52'h0; // @[playground/src/noop/tlb.scala 39:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (!(2'h0 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
        if (!(2'h3 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
          tag_13 <= _GEN_1011;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 39:26]
      tag_14 <= 52'h0; // @[playground/src/noop/tlb.scala 39:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (!(2'h0 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
        if (!(2'h3 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
          tag_14 <= _GEN_1012;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 39:26]
      tag_15 <= 52'h0; // @[playground/src/noop/tlb.scala 39:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (!(2'h0 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
        if (!(2'h3 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
          tag_15 <= _GEN_1013;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 40:26]
      paddr_0 <= 20'h0; // @[playground/src/noop/tlb.scala 40:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (!(2'h0 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
        if (!(2'h3 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
          paddr_0 <= _GEN_1030;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 40:26]
      paddr_1 <= 20'h0; // @[playground/src/noop/tlb.scala 40:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (!(2'h0 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
        if (!(2'h3 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
          paddr_1 <= _GEN_1031;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 40:26]
      paddr_2 <= 20'h0; // @[playground/src/noop/tlb.scala 40:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (!(2'h0 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
        if (!(2'h3 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
          paddr_2 <= _GEN_1032;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 40:26]
      paddr_3 <= 20'h0; // @[playground/src/noop/tlb.scala 40:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (!(2'h0 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
        if (!(2'h3 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
          paddr_3 <= _GEN_1033;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 40:26]
      paddr_4 <= 20'h0; // @[playground/src/noop/tlb.scala 40:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (!(2'h0 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
        if (!(2'h3 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
          paddr_4 <= _GEN_1034;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 40:26]
      paddr_5 <= 20'h0; // @[playground/src/noop/tlb.scala 40:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (!(2'h0 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
        if (!(2'h3 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
          paddr_5 <= _GEN_1035;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 40:26]
      paddr_6 <= 20'h0; // @[playground/src/noop/tlb.scala 40:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (!(2'h0 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
        if (!(2'h3 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
          paddr_6 <= _GEN_1036;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 40:26]
      paddr_7 <= 20'h0; // @[playground/src/noop/tlb.scala 40:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (!(2'h0 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
        if (!(2'h3 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
          paddr_7 <= _GEN_1037;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 40:26]
      paddr_8 <= 20'h0; // @[playground/src/noop/tlb.scala 40:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (!(2'h0 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
        if (!(2'h3 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
          paddr_8 <= _GEN_1038;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 40:26]
      paddr_9 <= 20'h0; // @[playground/src/noop/tlb.scala 40:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (!(2'h0 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
        if (!(2'h3 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
          paddr_9 <= _GEN_1039;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 40:26]
      paddr_10 <= 20'h0; // @[playground/src/noop/tlb.scala 40:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (!(2'h0 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
        if (!(2'h3 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
          paddr_10 <= _GEN_1040;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 40:26]
      paddr_11 <= 20'h0; // @[playground/src/noop/tlb.scala 40:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (!(2'h0 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
        if (!(2'h3 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
          paddr_11 <= _GEN_1041;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 40:26]
      paddr_12 <= 20'h0; // @[playground/src/noop/tlb.scala 40:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (!(2'h0 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
        if (!(2'h3 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
          paddr_12 <= _GEN_1042;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 40:26]
      paddr_13 <= 20'h0; // @[playground/src/noop/tlb.scala 40:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (!(2'h0 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
        if (!(2'h3 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
          paddr_13 <= _GEN_1043;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 40:26]
      paddr_14 <= 20'h0; // @[playground/src/noop/tlb.scala 40:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (!(2'h0 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
        if (!(2'h3 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
          paddr_14 <= _GEN_1044;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 40:26]
      paddr_15 <= 20'h0; // @[playground/src/noop/tlb.scala 40:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (!(2'h0 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
        if (!(2'h3 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
          paddr_15 <= _GEN_1045;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 41:26]
      info_0 <= 10'h0; // @[playground/src/noop/tlb.scala 41:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (2'h0 == state) begin // @[playground/src/noop/tlb.scala 136:22]
        if (!(~handshake)) begin // @[playground/src/noop/tlb.scala 139:33]
          info_0 <= _GEN_243;
        end
      end else if (!(2'h3 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
        info_0 <= _GEN_1078;
      end
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 41:26]
      info_1 <= 10'h0; // @[playground/src/noop/tlb.scala 41:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (2'h0 == state) begin // @[playground/src/noop/tlb.scala 136:22]
        if (!(~handshake)) begin // @[playground/src/noop/tlb.scala 139:33]
          info_1 <= _GEN_244;
        end
      end else if (!(2'h3 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
        info_1 <= _GEN_1079;
      end
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 41:26]
      info_2 <= 10'h0; // @[playground/src/noop/tlb.scala 41:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (2'h0 == state) begin // @[playground/src/noop/tlb.scala 136:22]
        if (!(~handshake)) begin // @[playground/src/noop/tlb.scala 139:33]
          info_2 <= _GEN_245;
        end
      end else if (!(2'h3 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
        info_2 <= _GEN_1080;
      end
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 41:26]
      info_3 <= 10'h0; // @[playground/src/noop/tlb.scala 41:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (2'h0 == state) begin // @[playground/src/noop/tlb.scala 136:22]
        if (!(~handshake)) begin // @[playground/src/noop/tlb.scala 139:33]
          info_3 <= _GEN_246;
        end
      end else if (!(2'h3 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
        info_3 <= _GEN_1081;
      end
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 41:26]
      info_4 <= 10'h0; // @[playground/src/noop/tlb.scala 41:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (2'h0 == state) begin // @[playground/src/noop/tlb.scala 136:22]
        if (!(~handshake)) begin // @[playground/src/noop/tlb.scala 139:33]
          info_4 <= _GEN_247;
        end
      end else if (!(2'h3 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
        info_4 <= _GEN_1082;
      end
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 41:26]
      info_5 <= 10'h0; // @[playground/src/noop/tlb.scala 41:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (2'h0 == state) begin // @[playground/src/noop/tlb.scala 136:22]
        if (!(~handshake)) begin // @[playground/src/noop/tlb.scala 139:33]
          info_5 <= _GEN_248;
        end
      end else if (!(2'h3 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
        info_5 <= _GEN_1083;
      end
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 41:26]
      info_6 <= 10'h0; // @[playground/src/noop/tlb.scala 41:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (2'h0 == state) begin // @[playground/src/noop/tlb.scala 136:22]
        if (!(~handshake)) begin // @[playground/src/noop/tlb.scala 139:33]
          info_6 <= _GEN_249;
        end
      end else if (!(2'h3 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
        info_6 <= _GEN_1084;
      end
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 41:26]
      info_7 <= 10'h0; // @[playground/src/noop/tlb.scala 41:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (2'h0 == state) begin // @[playground/src/noop/tlb.scala 136:22]
        if (!(~handshake)) begin // @[playground/src/noop/tlb.scala 139:33]
          info_7 <= _GEN_250;
        end
      end else if (!(2'h3 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
        info_7 <= _GEN_1085;
      end
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 41:26]
      info_8 <= 10'h0; // @[playground/src/noop/tlb.scala 41:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (2'h0 == state) begin // @[playground/src/noop/tlb.scala 136:22]
        if (!(~handshake)) begin // @[playground/src/noop/tlb.scala 139:33]
          info_8 <= _GEN_251;
        end
      end else if (!(2'h3 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
        info_8 <= _GEN_1086;
      end
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 41:26]
      info_9 <= 10'h0; // @[playground/src/noop/tlb.scala 41:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (2'h0 == state) begin // @[playground/src/noop/tlb.scala 136:22]
        if (!(~handshake)) begin // @[playground/src/noop/tlb.scala 139:33]
          info_9 <= _GEN_252;
        end
      end else if (!(2'h3 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
        info_9 <= _GEN_1087;
      end
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 41:26]
      info_10 <= 10'h0; // @[playground/src/noop/tlb.scala 41:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (2'h0 == state) begin // @[playground/src/noop/tlb.scala 136:22]
        if (!(~handshake)) begin // @[playground/src/noop/tlb.scala 139:33]
          info_10 <= _GEN_253;
        end
      end else if (!(2'h3 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
        info_10 <= _GEN_1088;
      end
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 41:26]
      info_11 <= 10'h0; // @[playground/src/noop/tlb.scala 41:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (2'h0 == state) begin // @[playground/src/noop/tlb.scala 136:22]
        if (!(~handshake)) begin // @[playground/src/noop/tlb.scala 139:33]
          info_11 <= _GEN_254;
        end
      end else if (!(2'h3 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
        info_11 <= _GEN_1089;
      end
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 41:26]
      info_12 <= 10'h0; // @[playground/src/noop/tlb.scala 41:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (2'h0 == state) begin // @[playground/src/noop/tlb.scala 136:22]
        if (!(~handshake)) begin // @[playground/src/noop/tlb.scala 139:33]
          info_12 <= _GEN_255;
        end
      end else if (!(2'h3 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
        info_12 <= _GEN_1090;
      end
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 41:26]
      info_13 <= 10'h0; // @[playground/src/noop/tlb.scala 41:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (2'h0 == state) begin // @[playground/src/noop/tlb.scala 136:22]
        if (!(~handshake)) begin // @[playground/src/noop/tlb.scala 139:33]
          info_13 <= _GEN_256;
        end
      end else if (!(2'h3 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
        info_13 <= _GEN_1091;
      end
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 41:26]
      info_14 <= 10'h0; // @[playground/src/noop/tlb.scala 41:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (2'h0 == state) begin // @[playground/src/noop/tlb.scala 136:22]
        if (!(~handshake)) begin // @[playground/src/noop/tlb.scala 139:33]
          info_14 <= _GEN_257;
        end
      end else if (!(2'h3 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
        info_14 <= _GEN_1092;
      end
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 41:26]
      info_15 <= 10'h0; // @[playground/src/noop/tlb.scala 41:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (2'h0 == state) begin // @[playground/src/noop/tlb.scala 136:22]
        if (!(~handshake)) begin // @[playground/src/noop/tlb.scala 139:33]
          info_15 <= _GEN_258;
        end
      end else if (!(2'h3 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
        info_15 <= _GEN_1093;
      end
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 42:30]
      pte_addr_0 <= 32'h0; // @[playground/src/noop/tlb.scala 42:30]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (!(2'h0 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
        if (!(2'h3 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
          pte_addr_0 <= _GEN_1046;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 42:30]
      pte_addr_1 <= 32'h0; // @[playground/src/noop/tlb.scala 42:30]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (!(2'h0 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
        if (!(2'h3 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
          pte_addr_1 <= _GEN_1047;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 42:30]
      pte_addr_2 <= 32'h0; // @[playground/src/noop/tlb.scala 42:30]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (!(2'h0 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
        if (!(2'h3 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
          pte_addr_2 <= _GEN_1048;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 42:30]
      pte_addr_3 <= 32'h0; // @[playground/src/noop/tlb.scala 42:30]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (!(2'h0 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
        if (!(2'h3 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
          pte_addr_3 <= _GEN_1049;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 42:30]
      pte_addr_4 <= 32'h0; // @[playground/src/noop/tlb.scala 42:30]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (!(2'h0 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
        if (!(2'h3 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
          pte_addr_4 <= _GEN_1050;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 42:30]
      pte_addr_5 <= 32'h0; // @[playground/src/noop/tlb.scala 42:30]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (!(2'h0 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
        if (!(2'h3 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
          pte_addr_5 <= _GEN_1051;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 42:30]
      pte_addr_6 <= 32'h0; // @[playground/src/noop/tlb.scala 42:30]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (!(2'h0 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
        if (!(2'h3 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
          pte_addr_6 <= _GEN_1052;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 42:30]
      pte_addr_7 <= 32'h0; // @[playground/src/noop/tlb.scala 42:30]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (!(2'h0 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
        if (!(2'h3 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
          pte_addr_7 <= _GEN_1053;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 42:30]
      pte_addr_8 <= 32'h0; // @[playground/src/noop/tlb.scala 42:30]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (!(2'h0 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
        if (!(2'h3 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
          pte_addr_8 <= _GEN_1054;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 42:30]
      pte_addr_9 <= 32'h0; // @[playground/src/noop/tlb.scala 42:30]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (!(2'h0 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
        if (!(2'h3 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
          pte_addr_9 <= _GEN_1055;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 42:30]
      pte_addr_10 <= 32'h0; // @[playground/src/noop/tlb.scala 42:30]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (!(2'h0 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
        if (!(2'h3 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
          pte_addr_10 <= _GEN_1056;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 42:30]
      pte_addr_11 <= 32'h0; // @[playground/src/noop/tlb.scala 42:30]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (!(2'h0 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
        if (!(2'h3 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
          pte_addr_11 <= _GEN_1057;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 42:30]
      pte_addr_12 <= 32'h0; // @[playground/src/noop/tlb.scala 42:30]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (!(2'h0 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
        if (!(2'h3 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
          pte_addr_12 <= _GEN_1058;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 42:30]
      pte_addr_13 <= 32'h0; // @[playground/src/noop/tlb.scala 42:30]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (!(2'h0 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
        if (!(2'h3 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
          pte_addr_13 <= _GEN_1059;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 42:30]
      pte_addr_14 <= 32'h0; // @[playground/src/noop/tlb.scala 42:30]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (!(2'h0 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
        if (!(2'h3 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
          pte_addr_14 <= _GEN_1060;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 42:30]
      pte_addr_15 <= 32'h0; // @[playground/src/noop/tlb.scala 42:30]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (!(2'h0 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
        if (!(2'h3 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
          pte_addr_15 <= _GEN_1061;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 43:30]
      pte_level_0 <= 2'h0; // @[playground/src/noop/tlb.scala 43:30]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (!(2'h0 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
        if (!(2'h3 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
          pte_level_0 <= _GEN_1062;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 43:30]
      pte_level_1 <= 2'h0; // @[playground/src/noop/tlb.scala 43:30]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (!(2'h0 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
        if (!(2'h3 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
          pte_level_1 <= _GEN_1063;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 43:30]
      pte_level_2 <= 2'h0; // @[playground/src/noop/tlb.scala 43:30]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (!(2'h0 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
        if (!(2'h3 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
          pte_level_2 <= _GEN_1064;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 43:30]
      pte_level_3 <= 2'h0; // @[playground/src/noop/tlb.scala 43:30]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (!(2'h0 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
        if (!(2'h3 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
          pte_level_3 <= _GEN_1065;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 43:30]
      pte_level_4 <= 2'h0; // @[playground/src/noop/tlb.scala 43:30]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (!(2'h0 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
        if (!(2'h3 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
          pte_level_4 <= _GEN_1066;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 43:30]
      pte_level_5 <= 2'h0; // @[playground/src/noop/tlb.scala 43:30]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (!(2'h0 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
        if (!(2'h3 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
          pte_level_5 <= _GEN_1067;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 43:30]
      pte_level_6 <= 2'h0; // @[playground/src/noop/tlb.scala 43:30]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (!(2'h0 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
        if (!(2'h3 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
          pte_level_6 <= _GEN_1068;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 43:30]
      pte_level_7 <= 2'h0; // @[playground/src/noop/tlb.scala 43:30]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (!(2'h0 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
        if (!(2'h3 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
          pte_level_7 <= _GEN_1069;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 43:30]
      pte_level_8 <= 2'h0; // @[playground/src/noop/tlb.scala 43:30]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (!(2'h0 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
        if (!(2'h3 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
          pte_level_8 <= _GEN_1070;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 43:30]
      pte_level_9 <= 2'h0; // @[playground/src/noop/tlb.scala 43:30]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (!(2'h0 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
        if (!(2'h3 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
          pte_level_9 <= _GEN_1071;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 43:30]
      pte_level_10 <= 2'h0; // @[playground/src/noop/tlb.scala 43:30]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (!(2'h0 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
        if (!(2'h3 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
          pte_level_10 <= _GEN_1072;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 43:30]
      pte_level_11 <= 2'h0; // @[playground/src/noop/tlb.scala 43:30]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (!(2'h0 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
        if (!(2'h3 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
          pte_level_11 <= _GEN_1073;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 43:30]
      pte_level_12 <= 2'h0; // @[playground/src/noop/tlb.scala 43:30]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (!(2'h0 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
        if (!(2'h3 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
          pte_level_12 <= _GEN_1074;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 43:30]
      pte_level_13 <= 2'h0; // @[playground/src/noop/tlb.scala 43:30]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (!(2'h0 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
        if (!(2'h3 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
          pte_level_13 <= _GEN_1075;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 43:30]
      pte_level_14 <= 2'h0; // @[playground/src/noop/tlb.scala 43:30]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (!(2'h0 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
        if (!(2'h3 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
          pte_level_14 <= _GEN_1076;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 43:30]
      pte_level_15 <= 2'h0; // @[playground/src/noop/tlb.scala 43:30]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (!(2'h0 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
        if (!(2'h3 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
          pte_level_15 <= _GEN_1077;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 44:26]
      valid_0 <= 1'h0; // @[playground/src/noop/tlb.scala 44:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (2'h0 == state) begin // @[playground/src/noop/tlb.scala 136:22]
        valid_0 <= _GEN_130;
      end else if (2'h3 == state) begin // @[playground/src/noop/tlb.scala 136:22]
        valid_0 <= _GEN_130;
      end else begin
        valid_0 <= _GEN_1014;
      end
    end else begin
      valid_0 <= _GEN_130;
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 44:26]
      valid_1 <= 1'h0; // @[playground/src/noop/tlb.scala 44:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (2'h0 == state) begin // @[playground/src/noop/tlb.scala 136:22]
        valid_1 <= _GEN_131;
      end else if (2'h3 == state) begin // @[playground/src/noop/tlb.scala 136:22]
        valid_1 <= _GEN_131;
      end else begin
        valid_1 <= _GEN_1015;
      end
    end else begin
      valid_1 <= _GEN_131;
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 44:26]
      valid_2 <= 1'h0; // @[playground/src/noop/tlb.scala 44:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (2'h0 == state) begin // @[playground/src/noop/tlb.scala 136:22]
        valid_2 <= _GEN_132;
      end else if (2'h3 == state) begin // @[playground/src/noop/tlb.scala 136:22]
        valid_2 <= _GEN_132;
      end else begin
        valid_2 <= _GEN_1016;
      end
    end else begin
      valid_2 <= _GEN_132;
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 44:26]
      valid_3 <= 1'h0; // @[playground/src/noop/tlb.scala 44:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (2'h0 == state) begin // @[playground/src/noop/tlb.scala 136:22]
        valid_3 <= _GEN_133;
      end else if (2'h3 == state) begin // @[playground/src/noop/tlb.scala 136:22]
        valid_3 <= _GEN_133;
      end else begin
        valid_3 <= _GEN_1017;
      end
    end else begin
      valid_3 <= _GEN_133;
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 44:26]
      valid_4 <= 1'h0; // @[playground/src/noop/tlb.scala 44:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (2'h0 == state) begin // @[playground/src/noop/tlb.scala 136:22]
        valid_4 <= _GEN_134;
      end else if (2'h3 == state) begin // @[playground/src/noop/tlb.scala 136:22]
        valid_4 <= _GEN_134;
      end else begin
        valid_4 <= _GEN_1018;
      end
    end else begin
      valid_4 <= _GEN_134;
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 44:26]
      valid_5 <= 1'h0; // @[playground/src/noop/tlb.scala 44:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (2'h0 == state) begin // @[playground/src/noop/tlb.scala 136:22]
        valid_5 <= _GEN_135;
      end else if (2'h3 == state) begin // @[playground/src/noop/tlb.scala 136:22]
        valid_5 <= _GEN_135;
      end else begin
        valid_5 <= _GEN_1019;
      end
    end else begin
      valid_5 <= _GEN_135;
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 44:26]
      valid_6 <= 1'h0; // @[playground/src/noop/tlb.scala 44:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (2'h0 == state) begin // @[playground/src/noop/tlb.scala 136:22]
        valid_6 <= _GEN_136;
      end else if (2'h3 == state) begin // @[playground/src/noop/tlb.scala 136:22]
        valid_6 <= _GEN_136;
      end else begin
        valid_6 <= _GEN_1020;
      end
    end else begin
      valid_6 <= _GEN_136;
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 44:26]
      valid_7 <= 1'h0; // @[playground/src/noop/tlb.scala 44:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (2'h0 == state) begin // @[playground/src/noop/tlb.scala 136:22]
        valid_7 <= _GEN_137;
      end else if (2'h3 == state) begin // @[playground/src/noop/tlb.scala 136:22]
        valid_7 <= _GEN_137;
      end else begin
        valid_7 <= _GEN_1021;
      end
    end else begin
      valid_7 <= _GEN_137;
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 44:26]
      valid_8 <= 1'h0; // @[playground/src/noop/tlb.scala 44:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (2'h0 == state) begin // @[playground/src/noop/tlb.scala 136:22]
        valid_8 <= _GEN_138;
      end else if (2'h3 == state) begin // @[playground/src/noop/tlb.scala 136:22]
        valid_8 <= _GEN_138;
      end else begin
        valid_8 <= _GEN_1022;
      end
    end else begin
      valid_8 <= _GEN_138;
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 44:26]
      valid_9 <= 1'h0; // @[playground/src/noop/tlb.scala 44:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (2'h0 == state) begin // @[playground/src/noop/tlb.scala 136:22]
        valid_9 <= _GEN_139;
      end else if (2'h3 == state) begin // @[playground/src/noop/tlb.scala 136:22]
        valid_9 <= _GEN_139;
      end else begin
        valid_9 <= _GEN_1023;
      end
    end else begin
      valid_9 <= _GEN_139;
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 44:26]
      valid_10 <= 1'h0; // @[playground/src/noop/tlb.scala 44:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (2'h0 == state) begin // @[playground/src/noop/tlb.scala 136:22]
        valid_10 <= _GEN_140;
      end else if (2'h3 == state) begin // @[playground/src/noop/tlb.scala 136:22]
        valid_10 <= _GEN_140;
      end else begin
        valid_10 <= _GEN_1024;
      end
    end else begin
      valid_10 <= _GEN_140;
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 44:26]
      valid_11 <= 1'h0; // @[playground/src/noop/tlb.scala 44:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (2'h0 == state) begin // @[playground/src/noop/tlb.scala 136:22]
        valid_11 <= _GEN_141;
      end else if (2'h3 == state) begin // @[playground/src/noop/tlb.scala 136:22]
        valid_11 <= _GEN_141;
      end else begin
        valid_11 <= _GEN_1025;
      end
    end else begin
      valid_11 <= _GEN_141;
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 44:26]
      valid_12 <= 1'h0; // @[playground/src/noop/tlb.scala 44:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (2'h0 == state) begin // @[playground/src/noop/tlb.scala 136:22]
        valid_12 <= _GEN_142;
      end else if (2'h3 == state) begin // @[playground/src/noop/tlb.scala 136:22]
        valid_12 <= _GEN_142;
      end else begin
        valid_12 <= _GEN_1026;
      end
    end else begin
      valid_12 <= _GEN_142;
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 44:26]
      valid_13 <= 1'h0; // @[playground/src/noop/tlb.scala 44:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (2'h0 == state) begin // @[playground/src/noop/tlb.scala 136:22]
        valid_13 <= _GEN_143;
      end else if (2'h3 == state) begin // @[playground/src/noop/tlb.scala 136:22]
        valid_13 <= _GEN_143;
      end else begin
        valid_13 <= _GEN_1027;
      end
    end else begin
      valid_13 <= _GEN_143;
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 44:26]
      valid_14 <= 1'h0; // @[playground/src/noop/tlb.scala 44:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (2'h0 == state) begin // @[playground/src/noop/tlb.scala 136:22]
        valid_14 <= _GEN_144;
      end else if (2'h3 == state) begin // @[playground/src/noop/tlb.scala 136:22]
        valid_14 <= _GEN_144;
      end else begin
        valid_14 <= _GEN_1028;
      end
    end else begin
      valid_14 <= _GEN_144;
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 44:26]
      valid_15 <= 1'h0; // @[playground/src/noop/tlb.scala 44:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (2'h0 == state) begin // @[playground/src/noop/tlb.scala 136:22]
        valid_15 <= _GEN_145;
      end else if (2'h3 == state) begin // @[playground/src/noop/tlb.scala 136:22]
        valid_15 <= _GEN_145;
      end else begin
        valid_15 <= _GEN_1029;
      end
    end else begin
      valid_15 <= _GEN_145;
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 46:30]
      pre_addr <= 64'h0; // @[playground/src/noop/tlb.scala 46:30]
    end else if (handshake) begin // @[playground/src/noop/tlb.scala 101:20]
      pre_addr <= io_va2pa_vaddr; // @[playground/src/noop/tlb.scala 103:18]
    end else if (io_va2pa_ready & io_va2pa_vvalid) begin // @[playground/src/noop/tlb.scala 54:44]
      pre_addr <= io_va2pa_vaddr; // @[playground/src/noop/tlb.scala 55:18]
    end
    pte_addr_r <= _GEN_1418[31:0]; // @[playground/src/noop/tlb.scala 47:{30,30}]
    if (reset) begin // @[playground/src/noop/tlb.scala 48:30]
      wpte_data_r <= 64'h0; // @[playground/src/noop/tlb.scala 48:30]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (2'h0 == state) begin // @[playground/src/noop/tlb.scala 136:22]
        if (!(~handshake)) begin // @[playground/src/noop/tlb.scala 139:33]
          wpte_data_r <= _GEN_242;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 49:30]
      dc_mode_r <= 5'h0; // @[playground/src/noop/tlb.scala 49:30]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (2'h0 == state) begin // @[playground/src/noop/tlb.scala 136:22]
        if (~handshake) begin // @[playground/src/noop/tlb.scala 139:33]
          dc_mode_r <= 5'h0; // @[playground/src/noop/tlb.scala 138:27]
        end else begin
          dc_mode_r <= _GEN_261;
        end
      end else if (2'h3 == state) begin // @[playground/src/noop/tlb.scala 136:22]
        dc_mode_r <= _GEN_294;
      end else begin
        dc_mode_r <= _GEN_992;
      end
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 51:30]
      out_valid_r <= 1'h0; // @[playground/src/noop/tlb.scala 51:30]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (2'h0 == state) begin // @[playground/src/noop/tlb.scala 136:22]
        if (~handshake) begin // @[playground/src/noop/tlb.scala 139:33]
          out_valid_r <= _GEN_150;
        end else begin
          out_valid_r <= _GEN_237;
        end
      end else begin
        out_valid_r <= _GEN_150;
      end
    end else begin
      out_valid_r <= io_va2pa_vvalid; // @[playground/src/noop/tlb.scala 232:21]
    end
    out_paddr_r <= _GEN_1419[31:0]; // @[playground/src/noop/tlb.scala 52:{30,30}]
    if (reset) begin // @[playground/src/noop/tlb.scala 53:30]
      out_excep_r_cause <= 64'h0; // @[playground/src/noop/tlb.scala 53:30]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (2'h0 == state) begin // @[playground/src/noop/tlb.scala 136:22]
        if (!(~handshake)) begin // @[playground/src/noop/tlb.scala 139:33]
          out_excep_r_cause <= _GEN_235;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 53:30]
      out_excep_r_tval <= 64'h0; // @[playground/src/noop/tlb.scala 53:30]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (2'h0 == state) begin // @[playground/src/noop/tlb.scala 136:22]
        if (!(~handshake)) begin // @[playground/src/noop/tlb.scala 139:33]
          out_excep_r_tval <= _GEN_236;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 53:30]
      out_excep_r_en <= 1'h0; // @[playground/src/noop/tlb.scala 53:30]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (2'h0 == state) begin // @[playground/src/noop/tlb.scala 136:22]
        if (~handshake) begin // @[playground/src/noop/tlb.scala 139:33]
          out_excep_r_en <= _GEN_151;
        end else begin
          out_excep_r_en <= _GEN_234;
        end
      end else if (2'h3 == state) begin // @[playground/src/noop/tlb.scala 136:22]
        out_excep_r_en <= _GEN_151;
      end else begin
        out_excep_r_en <= _GEN_996;
      end
    end else begin
      out_excep_r_en <= _GEN_151;
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 84:24]
      state <= 2'h0; // @[playground/src/noop/tlb.scala 84:24]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (2'h0 == state) begin // @[playground/src/noop/tlb.scala 136:22]
        if (!(~handshake)) begin // @[playground/src/noop/tlb.scala 139:33]
          state <= _GEN_239;
        end
      end else if (2'h3 == state) begin // @[playground/src/noop/tlb.scala 136:22]
        state <= _GEN_296;
      end else begin
        state <= _GEN_995;
      end
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 85:26]
      flush_r <= 1'h0; // @[playground/src/noop/tlb.scala 85:26]
    end else if (io_flush | flush_r) begin // @[playground/src/noop/tlb.scala 86:30]
      if (state == 2'h0) begin // @[playground/src/noop/tlb.scala 87:30]
        flush_r <= 1'h0; // @[playground/src/noop/tlb.scala 89:21]
      end else begin
        flush_r <= 1'h1; // @[playground/src/noop/tlb.scala 91:21]
      end
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 95:27]
      m_type_r <= 2'h0; // @[playground/src/noop/tlb.scala 95:27]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (2'h0 == state) begin // @[playground/src/noop/tlb.scala 136:22]
        if (!(~handshake)) begin // @[playground/src/noop/tlb.scala 139:33]
          m_type_r <= _GEN_260;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 130:27]
      select_r <= 4'h0; // @[playground/src/noop/tlb.scala 130:27]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (2'h0 == state) begin // @[playground/src/noop/tlb.scala 136:22]
        if (!(~handshake)) begin // @[playground/src/noop/tlb.scala 139:33]
          select_r <= _GEN_259;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 131:26]
      offset <= 8'h0; // @[playground/src/noop/tlb.scala 131:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (2'h0 == state) begin // @[playground/src/noop/tlb.scala 136:22]
        if (!(~handshake)) begin // @[playground/src/noop/tlb.scala 139:33]
          offset <= _GEN_262;
        end
      end else if (!(2'h3 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
        offset <= _GEN_993;
      end
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 132:26]
      level <= 2'h0; // @[playground/src/noop/tlb.scala 132:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (2'h0 == state) begin // @[playground/src/noop/tlb.scala 136:22]
        if (!(~handshake)) begin // @[playground/src/noop/tlb.scala 139:33]
          level <= _GEN_263;
        end
      end else if (!(2'h3 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
        level <= _GEN_994;
      end
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 134:28]
      wpte_hs_r <= 1'h0; // @[playground/src/noop/tlb.scala 134:28]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (2'h0 == state) begin // @[playground/src/noop/tlb.scala 136:22]
        if (!(~handshake)) begin // @[playground/src/noop/tlb.scala 139:33]
          wpte_hs_r <= _GEN_240;
        end
      end else if (2'h3 == state) begin // @[playground/src/noop/tlb.scala 136:22]
        wpte_hs_r <= _GEN_295;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  tag_0 = _RAND_0[51:0];
  _RAND_1 = {2{`RANDOM}};
  tag_1 = _RAND_1[51:0];
  _RAND_2 = {2{`RANDOM}};
  tag_2 = _RAND_2[51:0];
  _RAND_3 = {2{`RANDOM}};
  tag_3 = _RAND_3[51:0];
  _RAND_4 = {2{`RANDOM}};
  tag_4 = _RAND_4[51:0];
  _RAND_5 = {2{`RANDOM}};
  tag_5 = _RAND_5[51:0];
  _RAND_6 = {2{`RANDOM}};
  tag_6 = _RAND_6[51:0];
  _RAND_7 = {2{`RANDOM}};
  tag_7 = _RAND_7[51:0];
  _RAND_8 = {2{`RANDOM}};
  tag_8 = _RAND_8[51:0];
  _RAND_9 = {2{`RANDOM}};
  tag_9 = _RAND_9[51:0];
  _RAND_10 = {2{`RANDOM}};
  tag_10 = _RAND_10[51:0];
  _RAND_11 = {2{`RANDOM}};
  tag_11 = _RAND_11[51:0];
  _RAND_12 = {2{`RANDOM}};
  tag_12 = _RAND_12[51:0];
  _RAND_13 = {2{`RANDOM}};
  tag_13 = _RAND_13[51:0];
  _RAND_14 = {2{`RANDOM}};
  tag_14 = _RAND_14[51:0];
  _RAND_15 = {2{`RANDOM}};
  tag_15 = _RAND_15[51:0];
  _RAND_16 = {1{`RANDOM}};
  paddr_0 = _RAND_16[19:0];
  _RAND_17 = {1{`RANDOM}};
  paddr_1 = _RAND_17[19:0];
  _RAND_18 = {1{`RANDOM}};
  paddr_2 = _RAND_18[19:0];
  _RAND_19 = {1{`RANDOM}};
  paddr_3 = _RAND_19[19:0];
  _RAND_20 = {1{`RANDOM}};
  paddr_4 = _RAND_20[19:0];
  _RAND_21 = {1{`RANDOM}};
  paddr_5 = _RAND_21[19:0];
  _RAND_22 = {1{`RANDOM}};
  paddr_6 = _RAND_22[19:0];
  _RAND_23 = {1{`RANDOM}};
  paddr_7 = _RAND_23[19:0];
  _RAND_24 = {1{`RANDOM}};
  paddr_8 = _RAND_24[19:0];
  _RAND_25 = {1{`RANDOM}};
  paddr_9 = _RAND_25[19:0];
  _RAND_26 = {1{`RANDOM}};
  paddr_10 = _RAND_26[19:0];
  _RAND_27 = {1{`RANDOM}};
  paddr_11 = _RAND_27[19:0];
  _RAND_28 = {1{`RANDOM}};
  paddr_12 = _RAND_28[19:0];
  _RAND_29 = {1{`RANDOM}};
  paddr_13 = _RAND_29[19:0];
  _RAND_30 = {1{`RANDOM}};
  paddr_14 = _RAND_30[19:0];
  _RAND_31 = {1{`RANDOM}};
  paddr_15 = _RAND_31[19:0];
  _RAND_32 = {1{`RANDOM}};
  info_0 = _RAND_32[9:0];
  _RAND_33 = {1{`RANDOM}};
  info_1 = _RAND_33[9:0];
  _RAND_34 = {1{`RANDOM}};
  info_2 = _RAND_34[9:0];
  _RAND_35 = {1{`RANDOM}};
  info_3 = _RAND_35[9:0];
  _RAND_36 = {1{`RANDOM}};
  info_4 = _RAND_36[9:0];
  _RAND_37 = {1{`RANDOM}};
  info_5 = _RAND_37[9:0];
  _RAND_38 = {1{`RANDOM}};
  info_6 = _RAND_38[9:0];
  _RAND_39 = {1{`RANDOM}};
  info_7 = _RAND_39[9:0];
  _RAND_40 = {1{`RANDOM}};
  info_8 = _RAND_40[9:0];
  _RAND_41 = {1{`RANDOM}};
  info_9 = _RAND_41[9:0];
  _RAND_42 = {1{`RANDOM}};
  info_10 = _RAND_42[9:0];
  _RAND_43 = {1{`RANDOM}};
  info_11 = _RAND_43[9:0];
  _RAND_44 = {1{`RANDOM}};
  info_12 = _RAND_44[9:0];
  _RAND_45 = {1{`RANDOM}};
  info_13 = _RAND_45[9:0];
  _RAND_46 = {1{`RANDOM}};
  info_14 = _RAND_46[9:0];
  _RAND_47 = {1{`RANDOM}};
  info_15 = _RAND_47[9:0];
  _RAND_48 = {1{`RANDOM}};
  pte_addr_0 = _RAND_48[31:0];
  _RAND_49 = {1{`RANDOM}};
  pte_addr_1 = _RAND_49[31:0];
  _RAND_50 = {1{`RANDOM}};
  pte_addr_2 = _RAND_50[31:0];
  _RAND_51 = {1{`RANDOM}};
  pte_addr_3 = _RAND_51[31:0];
  _RAND_52 = {1{`RANDOM}};
  pte_addr_4 = _RAND_52[31:0];
  _RAND_53 = {1{`RANDOM}};
  pte_addr_5 = _RAND_53[31:0];
  _RAND_54 = {1{`RANDOM}};
  pte_addr_6 = _RAND_54[31:0];
  _RAND_55 = {1{`RANDOM}};
  pte_addr_7 = _RAND_55[31:0];
  _RAND_56 = {1{`RANDOM}};
  pte_addr_8 = _RAND_56[31:0];
  _RAND_57 = {1{`RANDOM}};
  pte_addr_9 = _RAND_57[31:0];
  _RAND_58 = {1{`RANDOM}};
  pte_addr_10 = _RAND_58[31:0];
  _RAND_59 = {1{`RANDOM}};
  pte_addr_11 = _RAND_59[31:0];
  _RAND_60 = {1{`RANDOM}};
  pte_addr_12 = _RAND_60[31:0];
  _RAND_61 = {1{`RANDOM}};
  pte_addr_13 = _RAND_61[31:0];
  _RAND_62 = {1{`RANDOM}};
  pte_addr_14 = _RAND_62[31:0];
  _RAND_63 = {1{`RANDOM}};
  pte_addr_15 = _RAND_63[31:0];
  _RAND_64 = {1{`RANDOM}};
  pte_level_0 = _RAND_64[1:0];
  _RAND_65 = {1{`RANDOM}};
  pte_level_1 = _RAND_65[1:0];
  _RAND_66 = {1{`RANDOM}};
  pte_level_2 = _RAND_66[1:0];
  _RAND_67 = {1{`RANDOM}};
  pte_level_3 = _RAND_67[1:0];
  _RAND_68 = {1{`RANDOM}};
  pte_level_4 = _RAND_68[1:0];
  _RAND_69 = {1{`RANDOM}};
  pte_level_5 = _RAND_69[1:0];
  _RAND_70 = {1{`RANDOM}};
  pte_level_6 = _RAND_70[1:0];
  _RAND_71 = {1{`RANDOM}};
  pte_level_7 = _RAND_71[1:0];
  _RAND_72 = {1{`RANDOM}};
  pte_level_8 = _RAND_72[1:0];
  _RAND_73 = {1{`RANDOM}};
  pte_level_9 = _RAND_73[1:0];
  _RAND_74 = {1{`RANDOM}};
  pte_level_10 = _RAND_74[1:0];
  _RAND_75 = {1{`RANDOM}};
  pte_level_11 = _RAND_75[1:0];
  _RAND_76 = {1{`RANDOM}};
  pte_level_12 = _RAND_76[1:0];
  _RAND_77 = {1{`RANDOM}};
  pte_level_13 = _RAND_77[1:0];
  _RAND_78 = {1{`RANDOM}};
  pte_level_14 = _RAND_78[1:0];
  _RAND_79 = {1{`RANDOM}};
  pte_level_15 = _RAND_79[1:0];
  _RAND_80 = {1{`RANDOM}};
  valid_0 = _RAND_80[0:0];
  _RAND_81 = {1{`RANDOM}};
  valid_1 = _RAND_81[0:0];
  _RAND_82 = {1{`RANDOM}};
  valid_2 = _RAND_82[0:0];
  _RAND_83 = {1{`RANDOM}};
  valid_3 = _RAND_83[0:0];
  _RAND_84 = {1{`RANDOM}};
  valid_4 = _RAND_84[0:0];
  _RAND_85 = {1{`RANDOM}};
  valid_5 = _RAND_85[0:0];
  _RAND_86 = {1{`RANDOM}};
  valid_6 = _RAND_86[0:0];
  _RAND_87 = {1{`RANDOM}};
  valid_7 = _RAND_87[0:0];
  _RAND_88 = {1{`RANDOM}};
  valid_8 = _RAND_88[0:0];
  _RAND_89 = {1{`RANDOM}};
  valid_9 = _RAND_89[0:0];
  _RAND_90 = {1{`RANDOM}};
  valid_10 = _RAND_90[0:0];
  _RAND_91 = {1{`RANDOM}};
  valid_11 = _RAND_91[0:0];
  _RAND_92 = {1{`RANDOM}};
  valid_12 = _RAND_92[0:0];
  _RAND_93 = {1{`RANDOM}};
  valid_13 = _RAND_93[0:0];
  _RAND_94 = {1{`RANDOM}};
  valid_14 = _RAND_94[0:0];
  _RAND_95 = {1{`RANDOM}};
  valid_15 = _RAND_95[0:0];
  _RAND_96 = {2{`RANDOM}};
  pre_addr = _RAND_96[63:0];
  _RAND_97 = {1{`RANDOM}};
  pte_addr_r = _RAND_97[31:0];
  _RAND_98 = {2{`RANDOM}};
  wpte_data_r = _RAND_98[63:0];
  _RAND_99 = {1{`RANDOM}};
  dc_mode_r = _RAND_99[4:0];
  _RAND_100 = {1{`RANDOM}};
  out_valid_r = _RAND_100[0:0];
  _RAND_101 = {1{`RANDOM}};
  out_paddr_r = _RAND_101[31:0];
  _RAND_102 = {2{`RANDOM}};
  out_excep_r_cause = _RAND_102[63:0];
  _RAND_103 = {2{`RANDOM}};
  out_excep_r_tval = _RAND_103[63:0];
  _RAND_104 = {1{`RANDOM}};
  out_excep_r_en = _RAND_104[0:0];
  _RAND_105 = {1{`RANDOM}};
  state = _RAND_105[1:0];
  _RAND_106 = {1{`RANDOM}};
  flush_r = _RAND_106[0:0];
  _RAND_107 = {1{`RANDOM}};
  m_type_r = _RAND_107[1:0];
  _RAND_108 = {1{`RANDOM}};
  select_r = _RAND_108[3:0];
  _RAND_109 = {1{`RANDOM}};
  offset = _RAND_109[7:0];
  _RAND_110 = {1{`RANDOM}};
  level = _RAND_110[1:0];
  _RAND_111 = {1{`RANDOM}};
  wpte_hs_r = _RAND_111[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TLB_1(
  input         clock,
  input         reset,
  input  [63:0] io_va2pa_vaddr, // @[playground/src/noop/tlb.scala 33:16]
  input         io_va2pa_vvalid, // @[playground/src/noop/tlb.scala 33:16]
  input  [1:0]  io_va2pa_m_type, // @[playground/src/noop/tlb.scala 33:16]
  output        io_va2pa_ready, // @[playground/src/noop/tlb.scala 33:16]
  output [31:0] io_va2pa_paddr, // @[playground/src/noop/tlb.scala 33:16]
  output        io_va2pa_pvalid, // @[playground/src/noop/tlb.scala 33:16]
  output [63:0] io_va2pa_tlb_excep_cause, // @[playground/src/noop/tlb.scala 33:16]
  output [63:0] io_va2pa_tlb_excep_tval, // @[playground/src/noop/tlb.scala 33:16]
  output        io_va2pa_tlb_excep_en, // @[playground/src/noop/tlb.scala 33:16]
  input  [1:0]  io_mmuState_priv, // @[playground/src/noop/tlb.scala 33:16]
  input  [63:0] io_mmuState_mstatus, // @[playground/src/noop/tlb.scala 33:16]
  input  [63:0] io_mmuState_satp, // @[playground/src/noop/tlb.scala 33:16]
  input         io_flush, // @[playground/src/noop/tlb.scala 33:16]
  output [31:0] io_dcacheRW_addr, // @[playground/src/noop/tlb.scala 33:16]
  input  [63:0] io_dcacheRW_rdata, // @[playground/src/noop/tlb.scala 33:16]
  input         io_dcacheRW_rvalid, // @[playground/src/noop/tlb.scala 33:16]
  output [63:0] io_dcacheRW_wdata, // @[playground/src/noop/tlb.scala 33:16]
  output [4:0]  io_dcacheRW_dc_mode, // @[playground/src/noop/tlb.scala 33:16]
  input         io_dcacheRW_ready // @[playground/src/noop/tlb.scala 33:16]
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [63:0] _RAND_12;
  reg [63:0] _RAND_13;
  reg [63:0] _RAND_14;
  reg [63:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [63:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [63:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [63:0] _RAND_102;
  reg [63:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
`endif // RANDOMIZE_REG_INIT
  wire  select_prng_clock; // @[src/main/scala/chisel3/util/random/PRNG.scala 91:22]
  wire  select_prng_reset; // @[src/main/scala/chisel3/util/random/PRNG.scala 91:22]
  wire  select_prng_io_out_0; // @[src/main/scala/chisel3/util/random/PRNG.scala 91:22]
  wire  select_prng_io_out_1; // @[src/main/scala/chisel3/util/random/PRNG.scala 91:22]
  wire  select_prng_io_out_2; // @[src/main/scala/chisel3/util/random/PRNG.scala 91:22]
  wire  select_prng_io_out_3; // @[src/main/scala/chisel3/util/random/PRNG.scala 91:22]
  reg [51:0] tag_0; // @[playground/src/noop/tlb.scala 39:26]
  reg [51:0] tag_1; // @[playground/src/noop/tlb.scala 39:26]
  reg [51:0] tag_2; // @[playground/src/noop/tlb.scala 39:26]
  reg [51:0] tag_3; // @[playground/src/noop/tlb.scala 39:26]
  reg [51:0] tag_4; // @[playground/src/noop/tlb.scala 39:26]
  reg [51:0] tag_5; // @[playground/src/noop/tlb.scala 39:26]
  reg [51:0] tag_6; // @[playground/src/noop/tlb.scala 39:26]
  reg [51:0] tag_7; // @[playground/src/noop/tlb.scala 39:26]
  reg [51:0] tag_8; // @[playground/src/noop/tlb.scala 39:26]
  reg [51:0] tag_9; // @[playground/src/noop/tlb.scala 39:26]
  reg [51:0] tag_10; // @[playground/src/noop/tlb.scala 39:26]
  reg [51:0] tag_11; // @[playground/src/noop/tlb.scala 39:26]
  reg [51:0] tag_12; // @[playground/src/noop/tlb.scala 39:26]
  reg [51:0] tag_13; // @[playground/src/noop/tlb.scala 39:26]
  reg [51:0] tag_14; // @[playground/src/noop/tlb.scala 39:26]
  reg [51:0] tag_15; // @[playground/src/noop/tlb.scala 39:26]
  reg [19:0] paddr_0; // @[playground/src/noop/tlb.scala 40:26]
  reg [19:0] paddr_1; // @[playground/src/noop/tlb.scala 40:26]
  reg [19:0] paddr_2; // @[playground/src/noop/tlb.scala 40:26]
  reg [19:0] paddr_3; // @[playground/src/noop/tlb.scala 40:26]
  reg [19:0] paddr_4; // @[playground/src/noop/tlb.scala 40:26]
  reg [19:0] paddr_5; // @[playground/src/noop/tlb.scala 40:26]
  reg [19:0] paddr_6; // @[playground/src/noop/tlb.scala 40:26]
  reg [19:0] paddr_7; // @[playground/src/noop/tlb.scala 40:26]
  reg [19:0] paddr_8; // @[playground/src/noop/tlb.scala 40:26]
  reg [19:0] paddr_9; // @[playground/src/noop/tlb.scala 40:26]
  reg [19:0] paddr_10; // @[playground/src/noop/tlb.scala 40:26]
  reg [19:0] paddr_11; // @[playground/src/noop/tlb.scala 40:26]
  reg [19:0] paddr_12; // @[playground/src/noop/tlb.scala 40:26]
  reg [19:0] paddr_13; // @[playground/src/noop/tlb.scala 40:26]
  reg [19:0] paddr_14; // @[playground/src/noop/tlb.scala 40:26]
  reg [19:0] paddr_15; // @[playground/src/noop/tlb.scala 40:26]
  reg [9:0] info_0; // @[playground/src/noop/tlb.scala 41:26]
  reg [9:0] info_1; // @[playground/src/noop/tlb.scala 41:26]
  reg [9:0] info_2; // @[playground/src/noop/tlb.scala 41:26]
  reg [9:0] info_3; // @[playground/src/noop/tlb.scala 41:26]
  reg [9:0] info_4; // @[playground/src/noop/tlb.scala 41:26]
  reg [9:0] info_5; // @[playground/src/noop/tlb.scala 41:26]
  reg [9:0] info_6; // @[playground/src/noop/tlb.scala 41:26]
  reg [9:0] info_7; // @[playground/src/noop/tlb.scala 41:26]
  reg [9:0] info_8; // @[playground/src/noop/tlb.scala 41:26]
  reg [9:0] info_9; // @[playground/src/noop/tlb.scala 41:26]
  reg [9:0] info_10; // @[playground/src/noop/tlb.scala 41:26]
  reg [9:0] info_11; // @[playground/src/noop/tlb.scala 41:26]
  reg [9:0] info_12; // @[playground/src/noop/tlb.scala 41:26]
  reg [9:0] info_13; // @[playground/src/noop/tlb.scala 41:26]
  reg [9:0] info_14; // @[playground/src/noop/tlb.scala 41:26]
  reg [9:0] info_15; // @[playground/src/noop/tlb.scala 41:26]
  reg [31:0] pte_addr_0; // @[playground/src/noop/tlb.scala 42:30]
  reg [31:0] pte_addr_1; // @[playground/src/noop/tlb.scala 42:30]
  reg [31:0] pte_addr_2; // @[playground/src/noop/tlb.scala 42:30]
  reg [31:0] pte_addr_3; // @[playground/src/noop/tlb.scala 42:30]
  reg [31:0] pte_addr_4; // @[playground/src/noop/tlb.scala 42:30]
  reg [31:0] pte_addr_5; // @[playground/src/noop/tlb.scala 42:30]
  reg [31:0] pte_addr_6; // @[playground/src/noop/tlb.scala 42:30]
  reg [31:0] pte_addr_7; // @[playground/src/noop/tlb.scala 42:30]
  reg [31:0] pte_addr_8; // @[playground/src/noop/tlb.scala 42:30]
  reg [31:0] pte_addr_9; // @[playground/src/noop/tlb.scala 42:30]
  reg [31:0] pte_addr_10; // @[playground/src/noop/tlb.scala 42:30]
  reg [31:0] pte_addr_11; // @[playground/src/noop/tlb.scala 42:30]
  reg [31:0] pte_addr_12; // @[playground/src/noop/tlb.scala 42:30]
  reg [31:0] pte_addr_13; // @[playground/src/noop/tlb.scala 42:30]
  reg [31:0] pte_addr_14; // @[playground/src/noop/tlb.scala 42:30]
  reg [31:0] pte_addr_15; // @[playground/src/noop/tlb.scala 42:30]
  reg [1:0] pte_level_0; // @[playground/src/noop/tlb.scala 43:30]
  reg [1:0] pte_level_1; // @[playground/src/noop/tlb.scala 43:30]
  reg [1:0] pte_level_2; // @[playground/src/noop/tlb.scala 43:30]
  reg [1:0] pte_level_3; // @[playground/src/noop/tlb.scala 43:30]
  reg [1:0] pte_level_4; // @[playground/src/noop/tlb.scala 43:30]
  reg [1:0] pte_level_5; // @[playground/src/noop/tlb.scala 43:30]
  reg [1:0] pte_level_6; // @[playground/src/noop/tlb.scala 43:30]
  reg [1:0] pte_level_7; // @[playground/src/noop/tlb.scala 43:30]
  reg [1:0] pte_level_8; // @[playground/src/noop/tlb.scala 43:30]
  reg [1:0] pte_level_9; // @[playground/src/noop/tlb.scala 43:30]
  reg [1:0] pte_level_10; // @[playground/src/noop/tlb.scala 43:30]
  reg [1:0] pte_level_11; // @[playground/src/noop/tlb.scala 43:30]
  reg [1:0] pte_level_12; // @[playground/src/noop/tlb.scala 43:30]
  reg [1:0] pte_level_13; // @[playground/src/noop/tlb.scala 43:30]
  reg [1:0] pte_level_14; // @[playground/src/noop/tlb.scala 43:30]
  reg [1:0] pte_level_15; // @[playground/src/noop/tlb.scala 43:30]
  reg  valid_0; // @[playground/src/noop/tlb.scala 44:26]
  reg  valid_1; // @[playground/src/noop/tlb.scala 44:26]
  reg  valid_2; // @[playground/src/noop/tlb.scala 44:26]
  reg  valid_3; // @[playground/src/noop/tlb.scala 44:26]
  reg  valid_4; // @[playground/src/noop/tlb.scala 44:26]
  reg  valid_5; // @[playground/src/noop/tlb.scala 44:26]
  reg  valid_6; // @[playground/src/noop/tlb.scala 44:26]
  reg  valid_7; // @[playground/src/noop/tlb.scala 44:26]
  reg  valid_8; // @[playground/src/noop/tlb.scala 44:26]
  reg  valid_9; // @[playground/src/noop/tlb.scala 44:26]
  reg  valid_10; // @[playground/src/noop/tlb.scala 44:26]
  reg  valid_11; // @[playground/src/noop/tlb.scala 44:26]
  reg  valid_12; // @[playground/src/noop/tlb.scala 44:26]
  reg  valid_13; // @[playground/src/noop/tlb.scala 44:26]
  reg  valid_14; // @[playground/src/noop/tlb.scala 44:26]
  reg  valid_15; // @[playground/src/noop/tlb.scala 44:26]
  reg [63:0] pre_addr; // @[playground/src/noop/tlb.scala 46:30]
  reg [31:0] pte_addr_r; // @[playground/src/noop/tlb.scala 47:30]
  reg [63:0] wpte_data_r; // @[playground/src/noop/tlb.scala 48:30]
  reg [4:0] dc_mode_r; // @[playground/src/noop/tlb.scala 49:30]
  reg  out_valid_r; // @[playground/src/noop/tlb.scala 51:30]
  reg [31:0] out_paddr_r; // @[playground/src/noop/tlb.scala 52:30]
  reg [63:0] out_excep_r_cause; // @[playground/src/noop/tlb.scala 53:30]
  reg [63:0] out_excep_r_tval; // @[playground/src/noop/tlb.scala 53:30]
  reg  out_excep_r_en; // @[playground/src/noop/tlb.scala 53:30]
  wire [51:0] inp_tag = io_va2pa_vaddr[63:12]; // @[playground/src/noop/tlb.scala 58:33]
  wire  _mode_T = io_va2pa_m_type == 2'h1; // @[playground/src/noop/tlb.scala 61:26]
  wire [1:0] _mode_T_3 = io_mmuState_mstatus[17] ? io_mmuState_mstatus[12:11] : io_mmuState_priv; // @[src/main/scala/chisel3/util/Mux.scala 47:70]
  wire [1:0] mode = _mode_T ? io_mmuState_priv : _mode_T_3; // @[src/main/scala/chisel3/util/Mux.scala 47:70]
  wire [3:0] mmuMode = mode == 2'h3 ? 4'h0 : io_mmuState_satp[63:60]; // @[playground/src/noop/tlb.scala 65:22]
  wire  is_Sv39 = mmuMode == 4'h8; // @[playground/src/noop/tlb.scala 66:27]
  wire [51:0] _tlb_tag_mask_T_4 = 2'h0 == pte_level_0 ? 52'hfffffffffffff : 52'h0; // @[src/main/scala/chisel3/util/Mux.scala 81:58]
  wire [51:0] _tlb_tag_mask_T_6 = 2'h1 == pte_level_0 ? 52'hffffffffffe00 : _tlb_tag_mask_T_4; // @[src/main/scala/chisel3/util/Mux.scala 81:58]
  wire [51:0] tlb_tag_mask = 2'h2 == pte_level_0 ? 52'hffffffffc0000 : _tlb_tag_mask_T_6; // @[src/main/scala/chisel3/util/Mux.scala 81:58]
  wire [51:0] _T_1 = inp_tag & tlb_tag_mask; // @[playground/src/noop/tlb.scala 73:24]
  wire [19:0] _GEN_2 = _T_1 == tag_0 & valid_0 ? paddr_0 : 20'h0; // @[playground/src/noop/tlb.scala 73:64 75:28 68:40]
  wire [9:0] _GEN_4 = _T_1 == tag_0 & valid_0 ? info_0 : 10'h0; // @[playground/src/noop/tlb.scala 73:64 77:28 68:86]
  wire [31:0] _GEN_5 = _T_1 == tag_0 & valid_0 ? pte_addr_0 : 32'h0; // @[playground/src/noop/tlb.scala 69:23 73:64 78:31]
  wire [1:0] _GEN_7 = _T_1 == tag_0 & valid_0 ? pte_level_0 : 2'h0; // @[playground/src/noop/tlb.scala 73:64 80:31 69:69]
  wire [51:0] _tlb_tag_mask_T_12 = 2'h0 == pte_level_1 ? 52'hfffffffffffff : 52'h0; // @[src/main/scala/chisel3/util/Mux.scala 81:58]
  wire [51:0] _tlb_tag_mask_T_14 = 2'h1 == pte_level_1 ? 52'hffffffffffe00 : _tlb_tag_mask_T_12; // @[src/main/scala/chisel3/util/Mux.scala 81:58]
  wire [51:0] tlb_tag_mask_1 = 2'h2 == pte_level_1 ? 52'hffffffffc0000 : _tlb_tag_mask_T_14; // @[src/main/scala/chisel3/util/Mux.scala 81:58]
  wire [51:0] _T_4 = inp_tag & tlb_tag_mask_1; // @[playground/src/noop/tlb.scala 73:24]
  wire  _T_6 = _T_4 == tag_1 & valid_1; // @[playground/src/noop/tlb.scala 73:52]
  wire [19:0] _GEN_9 = _T_4 == tag_1 & valid_1 ? paddr_1 : _GEN_2; // @[playground/src/noop/tlb.scala 73:64 75:28]
  wire [9:0] _GEN_11 = _T_4 == tag_1 & valid_1 ? info_1 : _GEN_4; // @[playground/src/noop/tlb.scala 73:64 77:28]
  wire [31:0] _GEN_12 = _T_4 == tag_1 & valid_1 ? pte_addr_1 : _GEN_5; // @[playground/src/noop/tlb.scala 73:64 78:31]
  wire [1:0] _GEN_14 = _T_4 == tag_1 & valid_1 ? pte_level_1 : _GEN_7; // @[playground/src/noop/tlb.scala 73:64 80:31]
  wire [51:0] _tlb_tag_mask_T_20 = 2'h0 == pte_level_2 ? 52'hfffffffffffff : 52'h0; // @[src/main/scala/chisel3/util/Mux.scala 81:58]
  wire [51:0] _tlb_tag_mask_T_22 = 2'h1 == pte_level_2 ? 52'hffffffffffe00 : _tlb_tag_mask_T_20; // @[src/main/scala/chisel3/util/Mux.scala 81:58]
  wire [51:0] tlb_tag_mask_2 = 2'h2 == pte_level_2 ? 52'hffffffffc0000 : _tlb_tag_mask_T_22; // @[src/main/scala/chisel3/util/Mux.scala 81:58]
  wire [51:0] _T_7 = inp_tag & tlb_tag_mask_2; // @[playground/src/noop/tlb.scala 73:24]
  wire [19:0] _GEN_16 = _T_7 == tag_2 & valid_2 ? paddr_2 : _GEN_9; // @[playground/src/noop/tlb.scala 73:64 75:28]
  wire [9:0] _GEN_18 = _T_7 == tag_2 & valid_2 ? info_2 : _GEN_11; // @[playground/src/noop/tlb.scala 73:64 77:28]
  wire [31:0] _GEN_19 = _T_7 == tag_2 & valid_2 ? pte_addr_2 : _GEN_12; // @[playground/src/noop/tlb.scala 73:64 78:31]
  wire [1:0] _GEN_20 = _T_7 == tag_2 & valid_2 ? 2'h2 : {{1'd0}, _T_6}; // @[playground/src/noop/tlb.scala 73:64 79:28]
  wire [1:0] _GEN_21 = _T_7 == tag_2 & valid_2 ? pte_level_2 : _GEN_14; // @[playground/src/noop/tlb.scala 73:64 80:31]
  wire [51:0] _tlb_tag_mask_T_28 = 2'h0 == pte_level_3 ? 52'hfffffffffffff : 52'h0; // @[src/main/scala/chisel3/util/Mux.scala 81:58]
  wire [51:0] _tlb_tag_mask_T_30 = 2'h1 == pte_level_3 ? 52'hffffffffffe00 : _tlb_tag_mask_T_28; // @[src/main/scala/chisel3/util/Mux.scala 81:58]
  wire [51:0] tlb_tag_mask_3 = 2'h2 == pte_level_3 ? 52'hffffffffc0000 : _tlb_tag_mask_T_30; // @[src/main/scala/chisel3/util/Mux.scala 81:58]
  wire [51:0] _T_10 = inp_tag & tlb_tag_mask_3; // @[playground/src/noop/tlb.scala 73:24]
  wire [19:0] _GEN_23 = _T_10 == tag_3 & valid_3 ? paddr_3 : _GEN_16; // @[playground/src/noop/tlb.scala 73:64 75:28]
  wire [9:0] _GEN_25 = _T_10 == tag_3 & valid_3 ? info_3 : _GEN_18; // @[playground/src/noop/tlb.scala 73:64 77:28]
  wire [31:0] _GEN_26 = _T_10 == tag_3 & valid_3 ? pte_addr_3 : _GEN_19; // @[playground/src/noop/tlb.scala 73:64 78:31]
  wire [1:0] _GEN_27 = _T_10 == tag_3 & valid_3 ? 2'h3 : _GEN_20; // @[playground/src/noop/tlb.scala 73:64 79:28]
  wire [1:0] _GEN_28 = _T_10 == tag_3 & valid_3 ? pte_level_3 : _GEN_21; // @[playground/src/noop/tlb.scala 73:64 80:31]
  wire [51:0] _tlb_tag_mask_T_36 = 2'h0 == pte_level_4 ? 52'hfffffffffffff : 52'h0; // @[src/main/scala/chisel3/util/Mux.scala 81:58]
  wire [51:0] _tlb_tag_mask_T_38 = 2'h1 == pte_level_4 ? 52'hffffffffffe00 : _tlb_tag_mask_T_36; // @[src/main/scala/chisel3/util/Mux.scala 81:58]
  wire [51:0] tlb_tag_mask_4 = 2'h2 == pte_level_4 ? 52'hffffffffc0000 : _tlb_tag_mask_T_38; // @[src/main/scala/chisel3/util/Mux.scala 81:58]
  wire [51:0] _T_13 = inp_tag & tlb_tag_mask_4; // @[playground/src/noop/tlb.scala 73:24]
  wire [19:0] _GEN_30 = _T_13 == tag_4 & valid_4 ? paddr_4 : _GEN_23; // @[playground/src/noop/tlb.scala 73:64 75:28]
  wire [9:0] _GEN_32 = _T_13 == tag_4 & valid_4 ? info_4 : _GEN_25; // @[playground/src/noop/tlb.scala 73:64 77:28]
  wire [31:0] _GEN_33 = _T_13 == tag_4 & valid_4 ? pte_addr_4 : _GEN_26; // @[playground/src/noop/tlb.scala 73:64 78:31]
  wire [2:0] _GEN_34 = _T_13 == tag_4 & valid_4 ? 3'h4 : {{1'd0}, _GEN_27}; // @[playground/src/noop/tlb.scala 73:64 79:28]
  wire [1:0] _GEN_35 = _T_13 == tag_4 & valid_4 ? pte_level_4 : _GEN_28; // @[playground/src/noop/tlb.scala 73:64 80:31]
  wire [51:0] _tlb_tag_mask_T_44 = 2'h0 == pte_level_5 ? 52'hfffffffffffff : 52'h0; // @[src/main/scala/chisel3/util/Mux.scala 81:58]
  wire [51:0] _tlb_tag_mask_T_46 = 2'h1 == pte_level_5 ? 52'hffffffffffe00 : _tlb_tag_mask_T_44; // @[src/main/scala/chisel3/util/Mux.scala 81:58]
  wire [51:0] tlb_tag_mask_5 = 2'h2 == pte_level_5 ? 52'hffffffffc0000 : _tlb_tag_mask_T_46; // @[src/main/scala/chisel3/util/Mux.scala 81:58]
  wire [51:0] _T_16 = inp_tag & tlb_tag_mask_5; // @[playground/src/noop/tlb.scala 73:24]
  wire [19:0] _GEN_37 = _T_16 == tag_5 & valid_5 ? paddr_5 : _GEN_30; // @[playground/src/noop/tlb.scala 73:64 75:28]
  wire [9:0] _GEN_39 = _T_16 == tag_5 & valid_5 ? info_5 : _GEN_32; // @[playground/src/noop/tlb.scala 73:64 77:28]
  wire [31:0] _GEN_40 = _T_16 == tag_5 & valid_5 ? pte_addr_5 : _GEN_33; // @[playground/src/noop/tlb.scala 73:64 78:31]
  wire [2:0] _GEN_41 = _T_16 == tag_5 & valid_5 ? 3'h5 : _GEN_34; // @[playground/src/noop/tlb.scala 73:64 79:28]
  wire [1:0] _GEN_42 = _T_16 == tag_5 & valid_5 ? pte_level_5 : _GEN_35; // @[playground/src/noop/tlb.scala 73:64 80:31]
  wire [51:0] _tlb_tag_mask_T_52 = 2'h0 == pte_level_6 ? 52'hfffffffffffff : 52'h0; // @[src/main/scala/chisel3/util/Mux.scala 81:58]
  wire [51:0] _tlb_tag_mask_T_54 = 2'h1 == pte_level_6 ? 52'hffffffffffe00 : _tlb_tag_mask_T_52; // @[src/main/scala/chisel3/util/Mux.scala 81:58]
  wire [51:0] tlb_tag_mask_6 = 2'h2 == pte_level_6 ? 52'hffffffffc0000 : _tlb_tag_mask_T_54; // @[src/main/scala/chisel3/util/Mux.scala 81:58]
  wire [51:0] _T_19 = inp_tag & tlb_tag_mask_6; // @[playground/src/noop/tlb.scala 73:24]
  wire [19:0] _GEN_44 = _T_19 == tag_6 & valid_6 ? paddr_6 : _GEN_37; // @[playground/src/noop/tlb.scala 73:64 75:28]
  wire [9:0] _GEN_46 = _T_19 == tag_6 & valid_6 ? info_6 : _GEN_39; // @[playground/src/noop/tlb.scala 73:64 77:28]
  wire [31:0] _GEN_47 = _T_19 == tag_6 & valid_6 ? pte_addr_6 : _GEN_40; // @[playground/src/noop/tlb.scala 73:64 78:31]
  wire [2:0] _GEN_48 = _T_19 == tag_6 & valid_6 ? 3'h6 : _GEN_41; // @[playground/src/noop/tlb.scala 73:64 79:28]
  wire [1:0] _GEN_49 = _T_19 == tag_6 & valid_6 ? pte_level_6 : _GEN_42; // @[playground/src/noop/tlb.scala 73:64 80:31]
  wire [51:0] _tlb_tag_mask_T_60 = 2'h0 == pte_level_7 ? 52'hfffffffffffff : 52'h0; // @[src/main/scala/chisel3/util/Mux.scala 81:58]
  wire [51:0] _tlb_tag_mask_T_62 = 2'h1 == pte_level_7 ? 52'hffffffffffe00 : _tlb_tag_mask_T_60; // @[src/main/scala/chisel3/util/Mux.scala 81:58]
  wire [51:0] tlb_tag_mask_7 = 2'h2 == pte_level_7 ? 52'hffffffffc0000 : _tlb_tag_mask_T_62; // @[src/main/scala/chisel3/util/Mux.scala 81:58]
  wire [51:0] _T_22 = inp_tag & tlb_tag_mask_7; // @[playground/src/noop/tlb.scala 73:24]
  wire [19:0] _GEN_51 = _T_22 == tag_7 & valid_7 ? paddr_7 : _GEN_44; // @[playground/src/noop/tlb.scala 73:64 75:28]
  wire [9:0] _GEN_53 = _T_22 == tag_7 & valid_7 ? info_7 : _GEN_46; // @[playground/src/noop/tlb.scala 73:64 77:28]
  wire [31:0] _GEN_54 = _T_22 == tag_7 & valid_7 ? pte_addr_7 : _GEN_47; // @[playground/src/noop/tlb.scala 73:64 78:31]
  wire [2:0] _GEN_55 = _T_22 == tag_7 & valid_7 ? 3'h7 : _GEN_48; // @[playground/src/noop/tlb.scala 73:64 79:28]
  wire [1:0] _GEN_56 = _T_22 == tag_7 & valid_7 ? pte_level_7 : _GEN_49; // @[playground/src/noop/tlb.scala 73:64 80:31]
  wire [51:0] _tlb_tag_mask_T_68 = 2'h0 == pte_level_8 ? 52'hfffffffffffff : 52'h0; // @[src/main/scala/chisel3/util/Mux.scala 81:58]
  wire [51:0] _tlb_tag_mask_T_70 = 2'h1 == pte_level_8 ? 52'hffffffffffe00 : _tlb_tag_mask_T_68; // @[src/main/scala/chisel3/util/Mux.scala 81:58]
  wire [51:0] tlb_tag_mask_8 = 2'h2 == pte_level_8 ? 52'hffffffffc0000 : _tlb_tag_mask_T_70; // @[src/main/scala/chisel3/util/Mux.scala 81:58]
  wire [51:0] _T_25 = inp_tag & tlb_tag_mask_8; // @[playground/src/noop/tlb.scala 73:24]
  wire [19:0] _GEN_58 = _T_25 == tag_8 & valid_8 ? paddr_8 : _GEN_51; // @[playground/src/noop/tlb.scala 73:64 75:28]
  wire [9:0] _GEN_60 = _T_25 == tag_8 & valid_8 ? info_8 : _GEN_53; // @[playground/src/noop/tlb.scala 73:64 77:28]
  wire [31:0] _GEN_61 = _T_25 == tag_8 & valid_8 ? pte_addr_8 : _GEN_54; // @[playground/src/noop/tlb.scala 73:64 78:31]
  wire [3:0] _GEN_62 = _T_25 == tag_8 & valid_8 ? 4'h8 : {{1'd0}, _GEN_55}; // @[playground/src/noop/tlb.scala 73:64 79:28]
  wire [1:0] _GEN_63 = _T_25 == tag_8 & valid_8 ? pte_level_8 : _GEN_56; // @[playground/src/noop/tlb.scala 73:64 80:31]
  wire [51:0] _tlb_tag_mask_T_76 = 2'h0 == pte_level_9 ? 52'hfffffffffffff : 52'h0; // @[src/main/scala/chisel3/util/Mux.scala 81:58]
  wire [51:0] _tlb_tag_mask_T_78 = 2'h1 == pte_level_9 ? 52'hffffffffffe00 : _tlb_tag_mask_T_76; // @[src/main/scala/chisel3/util/Mux.scala 81:58]
  wire [51:0] tlb_tag_mask_9 = 2'h2 == pte_level_9 ? 52'hffffffffc0000 : _tlb_tag_mask_T_78; // @[src/main/scala/chisel3/util/Mux.scala 81:58]
  wire [51:0] _T_28 = inp_tag & tlb_tag_mask_9; // @[playground/src/noop/tlb.scala 73:24]
  wire  _GEN_64 = _T_28 == tag_9 & valid_9 | (_T_25 == tag_8 & valid_8 | (_T_22 == tag_7 & valid_7 | (_T_19 == tag_6 &
    valid_6 | (_T_16 == tag_5 & valid_5 | (_T_13 == tag_4 & valid_4 | (_T_10 == tag_3 & valid_3 | (_T_7 == tag_2 &
    valid_2 | (_T_4 == tag_1 & valid_1 | _T_1 == tag_0 & valid_0)))))))); // @[playground/src/noop/tlb.scala 73:64 74:28]
  wire [19:0] _GEN_65 = _T_28 == tag_9 & valid_9 ? paddr_9 : _GEN_58; // @[playground/src/noop/tlb.scala 73:64 75:28]
  wire [9:0] _GEN_67 = _T_28 == tag_9 & valid_9 ? info_9 : _GEN_60; // @[playground/src/noop/tlb.scala 73:64 77:28]
  wire [31:0] _GEN_68 = _T_28 == tag_9 & valid_9 ? pte_addr_9 : _GEN_61; // @[playground/src/noop/tlb.scala 73:64 78:31]
  wire [3:0] _GEN_69 = _T_28 == tag_9 & valid_9 ? 4'h9 : _GEN_62; // @[playground/src/noop/tlb.scala 73:64 79:28]
  wire [1:0] _GEN_70 = _T_28 == tag_9 & valid_9 ? pte_level_9 : _GEN_63; // @[playground/src/noop/tlb.scala 73:64 80:31]
  wire [51:0] _tlb_tag_mask_T_84 = 2'h0 == pte_level_10 ? 52'hfffffffffffff : 52'h0; // @[src/main/scala/chisel3/util/Mux.scala 81:58]
  wire [51:0] _tlb_tag_mask_T_86 = 2'h1 == pte_level_10 ? 52'hffffffffffe00 : _tlb_tag_mask_T_84; // @[src/main/scala/chisel3/util/Mux.scala 81:58]
  wire [51:0] tlb_tag_mask_10 = 2'h2 == pte_level_10 ? 52'hffffffffc0000 : _tlb_tag_mask_T_86; // @[src/main/scala/chisel3/util/Mux.scala 81:58]
  wire [51:0] _T_31 = inp_tag & tlb_tag_mask_10; // @[playground/src/noop/tlb.scala 73:24]
  wire [19:0] _GEN_72 = _T_31 == tag_10 & valid_10 ? paddr_10 : _GEN_65; // @[playground/src/noop/tlb.scala 73:64 75:28]
  wire [9:0] _GEN_74 = _T_31 == tag_10 & valid_10 ? info_10 : _GEN_67; // @[playground/src/noop/tlb.scala 73:64 77:28]
  wire [31:0] _GEN_75 = _T_31 == tag_10 & valid_10 ? pte_addr_10 : _GEN_68; // @[playground/src/noop/tlb.scala 73:64 78:31]
  wire [3:0] _GEN_76 = _T_31 == tag_10 & valid_10 ? 4'ha : _GEN_69; // @[playground/src/noop/tlb.scala 73:64 79:28]
  wire [1:0] _GEN_77 = _T_31 == tag_10 & valid_10 ? pte_level_10 : _GEN_70; // @[playground/src/noop/tlb.scala 73:64 80:31]
  wire [51:0] _tlb_tag_mask_T_92 = 2'h0 == pte_level_11 ? 52'hfffffffffffff : 52'h0; // @[src/main/scala/chisel3/util/Mux.scala 81:58]
  wire [51:0] _tlb_tag_mask_T_94 = 2'h1 == pte_level_11 ? 52'hffffffffffe00 : _tlb_tag_mask_T_92; // @[src/main/scala/chisel3/util/Mux.scala 81:58]
  wire [51:0] tlb_tag_mask_11 = 2'h2 == pte_level_11 ? 52'hffffffffc0000 : _tlb_tag_mask_T_94; // @[src/main/scala/chisel3/util/Mux.scala 81:58]
  wire [51:0] _T_34 = inp_tag & tlb_tag_mask_11; // @[playground/src/noop/tlb.scala 73:24]
  wire [19:0] _GEN_79 = _T_34 == tag_11 & valid_11 ? paddr_11 : _GEN_72; // @[playground/src/noop/tlb.scala 73:64 75:28]
  wire [9:0] _GEN_81 = _T_34 == tag_11 & valid_11 ? info_11 : _GEN_74; // @[playground/src/noop/tlb.scala 73:64 77:28]
  wire [31:0] _GEN_82 = _T_34 == tag_11 & valid_11 ? pte_addr_11 : _GEN_75; // @[playground/src/noop/tlb.scala 73:64 78:31]
  wire [3:0] _GEN_83 = _T_34 == tag_11 & valid_11 ? 4'hb : _GEN_76; // @[playground/src/noop/tlb.scala 73:64 79:28]
  wire [1:0] _GEN_84 = _T_34 == tag_11 & valid_11 ? pte_level_11 : _GEN_77; // @[playground/src/noop/tlb.scala 73:64 80:31]
  wire [51:0] _tlb_tag_mask_T_100 = 2'h0 == pte_level_12 ? 52'hfffffffffffff : 52'h0; // @[src/main/scala/chisel3/util/Mux.scala 81:58]
  wire [51:0] _tlb_tag_mask_T_102 = 2'h1 == pte_level_12 ? 52'hffffffffffe00 : _tlb_tag_mask_T_100; // @[src/main/scala/chisel3/util/Mux.scala 81:58]
  wire [51:0] tlb_tag_mask_12 = 2'h2 == pte_level_12 ? 52'hffffffffc0000 : _tlb_tag_mask_T_102; // @[src/main/scala/chisel3/util/Mux.scala 81:58]
  wire [51:0] _T_37 = inp_tag & tlb_tag_mask_12; // @[playground/src/noop/tlb.scala 73:24]
  wire [19:0] _GEN_86 = _T_37 == tag_12 & valid_12 ? paddr_12 : _GEN_79; // @[playground/src/noop/tlb.scala 73:64 75:28]
  wire [9:0] _GEN_88 = _T_37 == tag_12 & valid_12 ? info_12 : _GEN_81; // @[playground/src/noop/tlb.scala 73:64 77:28]
  wire [31:0] _GEN_89 = _T_37 == tag_12 & valid_12 ? pte_addr_12 : _GEN_82; // @[playground/src/noop/tlb.scala 73:64 78:31]
  wire [3:0] _GEN_90 = _T_37 == tag_12 & valid_12 ? 4'hc : _GEN_83; // @[playground/src/noop/tlb.scala 73:64 79:28]
  wire [1:0] _GEN_91 = _T_37 == tag_12 & valid_12 ? pte_level_12 : _GEN_84; // @[playground/src/noop/tlb.scala 73:64 80:31]
  wire [51:0] _tlb_tag_mask_T_108 = 2'h0 == pte_level_13 ? 52'hfffffffffffff : 52'h0; // @[src/main/scala/chisel3/util/Mux.scala 81:58]
  wire [51:0] _tlb_tag_mask_T_110 = 2'h1 == pte_level_13 ? 52'hffffffffffe00 : _tlb_tag_mask_T_108; // @[src/main/scala/chisel3/util/Mux.scala 81:58]
  wire [51:0] tlb_tag_mask_13 = 2'h2 == pte_level_13 ? 52'hffffffffc0000 : _tlb_tag_mask_T_110; // @[src/main/scala/chisel3/util/Mux.scala 81:58]
  wire [51:0] _T_40 = inp_tag & tlb_tag_mask_13; // @[playground/src/noop/tlb.scala 73:24]
  wire [19:0] _GEN_93 = _T_40 == tag_13 & valid_13 ? paddr_13 : _GEN_86; // @[playground/src/noop/tlb.scala 73:64 75:28]
  wire [9:0] _GEN_95 = _T_40 == tag_13 & valid_13 ? info_13 : _GEN_88; // @[playground/src/noop/tlb.scala 73:64 77:28]
  wire [31:0] _GEN_96 = _T_40 == tag_13 & valid_13 ? pte_addr_13 : _GEN_89; // @[playground/src/noop/tlb.scala 73:64 78:31]
  wire [3:0] _GEN_97 = _T_40 == tag_13 & valid_13 ? 4'hd : _GEN_90; // @[playground/src/noop/tlb.scala 73:64 79:28]
  wire [1:0] _GEN_98 = _T_40 == tag_13 & valid_13 ? pte_level_13 : _GEN_91; // @[playground/src/noop/tlb.scala 73:64 80:31]
  wire [51:0] _tlb_tag_mask_T_116 = 2'h0 == pte_level_14 ? 52'hfffffffffffff : 52'h0; // @[src/main/scala/chisel3/util/Mux.scala 81:58]
  wire [51:0] _tlb_tag_mask_T_118 = 2'h1 == pte_level_14 ? 52'hffffffffffe00 : _tlb_tag_mask_T_116; // @[src/main/scala/chisel3/util/Mux.scala 81:58]
  wire [51:0] tlb_tag_mask_14 = 2'h2 == pte_level_14 ? 52'hffffffffc0000 : _tlb_tag_mask_T_118; // @[src/main/scala/chisel3/util/Mux.scala 81:58]
  wire [51:0] _T_43 = inp_tag & tlb_tag_mask_14; // @[playground/src/noop/tlb.scala 73:24]
  wire [19:0] _GEN_100 = _T_43 == tag_14 & valid_14 ? paddr_14 : _GEN_93; // @[playground/src/noop/tlb.scala 73:64 75:28]
  wire [9:0] _GEN_102 = _T_43 == tag_14 & valid_14 ? info_14 : _GEN_95; // @[playground/src/noop/tlb.scala 73:64 77:28]
  wire [31:0] _GEN_103 = _T_43 == tag_14 & valid_14 ? pte_addr_14 : _GEN_96; // @[playground/src/noop/tlb.scala 73:64 78:31]
  wire [3:0] _GEN_104 = _T_43 == tag_14 & valid_14 ? 4'he : _GEN_97; // @[playground/src/noop/tlb.scala 73:64 79:28]
  wire [1:0] _GEN_105 = _T_43 == tag_14 & valid_14 ? pte_level_14 : _GEN_98; // @[playground/src/noop/tlb.scala 73:64 80:31]
  wire [51:0] _tlb_tag_mask_T_124 = 2'h0 == pte_level_15 ? 52'hfffffffffffff : 52'h0; // @[src/main/scala/chisel3/util/Mux.scala 81:58]
  wire [51:0] _tlb_tag_mask_T_126 = 2'h1 == pte_level_15 ? 52'hffffffffffe00 : _tlb_tag_mask_T_124; // @[src/main/scala/chisel3/util/Mux.scala 81:58]
  wire [51:0] tlb_tag_mask_15 = 2'h2 == pte_level_15 ? 52'hffffffffc0000 : _tlb_tag_mask_T_126; // @[src/main/scala/chisel3/util/Mux.scala 81:58]
  wire [51:0] _T_46 = inp_tag & tlb_tag_mask_15; // @[playground/src/noop/tlb.scala 73:24]
  wire  tlbMsg_tlbHit = _T_46 == tag_15 & valid_15 | (_T_43 == tag_14 & valid_14 | (_T_40 == tag_13 & valid_13 | (_T_37
     == tag_12 & valid_12 | (_T_34 == tag_11 & valid_11 | (_T_31 == tag_10 & valid_10 | _GEN_64))))); // @[playground/src/noop/tlb.scala 73:64 74:28]
  wire [19:0] tlbMsg_tlbPa = _T_46 == tag_15 & valid_15 ? paddr_15 : _GEN_100; // @[playground/src/noop/tlb.scala 73:64 75:28]
  wire [9:0] tlbMsg_tlbInfo = _T_46 == tag_15 & valid_15 ? info_15 : _GEN_102; // @[playground/src/noop/tlb.scala 73:64 77:28]
  wire [31:0] tlbMsg_tlbPteAddr = _T_46 == tag_15 & valid_15 ? pte_addr_15 : _GEN_103; // @[playground/src/noop/tlb.scala 73:64 78:31]
  wire [3:0] tlbMsg_tlbIdx = _T_46 == tag_15 & valid_15 ? 4'hf : _GEN_104; // @[playground/src/noop/tlb.scala 73:64 79:28]
  wire [1:0] tlbMsg_tlbLevel = _T_46 == tag_15 & valid_15 ? pte_level_15 : _GEN_105; // @[playground/src/noop/tlb.scala 73:64 80:31]
  reg [1:0] state; // @[playground/src/noop/tlb.scala 84:24]
  reg  flush_r; // @[playground/src/noop/tlb.scala 85:26]
  wire  _T_50 = state == 2'h0; // @[playground/src/noop/tlb.scala 87:20]
  wire  _GEN_113 = state == 2'h0 ? 1'h0 : valid_0; // @[playground/src/noop/tlb.scala 87:30 88:19 44:26]
  wire  _GEN_114 = state == 2'h0 ? 1'h0 : valid_1; // @[playground/src/noop/tlb.scala 87:30 88:19 44:26]
  wire  _GEN_115 = state == 2'h0 ? 1'h0 : valid_2; // @[playground/src/noop/tlb.scala 87:30 88:19 44:26]
  wire  _GEN_116 = state == 2'h0 ? 1'h0 : valid_3; // @[playground/src/noop/tlb.scala 87:30 88:19 44:26]
  wire  _GEN_117 = state == 2'h0 ? 1'h0 : valid_4; // @[playground/src/noop/tlb.scala 87:30 88:19 44:26]
  wire  _GEN_118 = state == 2'h0 ? 1'h0 : valid_5; // @[playground/src/noop/tlb.scala 87:30 88:19 44:26]
  wire  _GEN_119 = state == 2'h0 ? 1'h0 : valid_6; // @[playground/src/noop/tlb.scala 87:30 88:19 44:26]
  wire  _GEN_120 = state == 2'h0 ? 1'h0 : valid_7; // @[playground/src/noop/tlb.scala 87:30 88:19 44:26]
  wire  _GEN_121 = state == 2'h0 ? 1'h0 : valid_8; // @[playground/src/noop/tlb.scala 87:30 88:19 44:26]
  wire  _GEN_122 = state == 2'h0 ? 1'h0 : valid_9; // @[playground/src/noop/tlb.scala 87:30 88:19 44:26]
  wire  _GEN_123 = state == 2'h0 ? 1'h0 : valid_10; // @[playground/src/noop/tlb.scala 87:30 88:19 44:26]
  wire  _GEN_124 = state == 2'h0 ? 1'h0 : valid_11; // @[playground/src/noop/tlb.scala 87:30 88:19 44:26]
  wire  _GEN_125 = state == 2'h0 ? 1'h0 : valid_12; // @[playground/src/noop/tlb.scala 87:30 88:19 44:26]
  wire  _GEN_126 = state == 2'h0 ? 1'h0 : valid_13; // @[playground/src/noop/tlb.scala 87:30 88:19 44:26]
  wire  _GEN_127 = state == 2'h0 ? 1'h0 : valid_14; // @[playground/src/noop/tlb.scala 87:30 88:19 44:26]
  wire  _GEN_128 = state == 2'h0 ? 1'h0 : valid_15; // @[playground/src/noop/tlb.scala 87:30 88:19 44:26]
  wire  _GEN_130 = io_flush | flush_r ? _GEN_113 : valid_0; // @[playground/src/noop/tlb.scala 44:26 86:30]
  wire  _GEN_131 = io_flush | flush_r ? _GEN_114 : valid_1; // @[playground/src/noop/tlb.scala 44:26 86:30]
  wire  _GEN_132 = io_flush | flush_r ? _GEN_115 : valid_2; // @[playground/src/noop/tlb.scala 44:26 86:30]
  wire  _GEN_133 = io_flush | flush_r ? _GEN_116 : valid_3; // @[playground/src/noop/tlb.scala 44:26 86:30]
  wire  _GEN_134 = io_flush | flush_r ? _GEN_117 : valid_4; // @[playground/src/noop/tlb.scala 44:26 86:30]
  wire  _GEN_135 = io_flush | flush_r ? _GEN_118 : valid_5; // @[playground/src/noop/tlb.scala 44:26 86:30]
  wire  _GEN_136 = io_flush | flush_r ? _GEN_119 : valid_6; // @[playground/src/noop/tlb.scala 44:26 86:30]
  wire  _GEN_137 = io_flush | flush_r ? _GEN_120 : valid_7; // @[playground/src/noop/tlb.scala 44:26 86:30]
  wire  _GEN_138 = io_flush | flush_r ? _GEN_121 : valid_8; // @[playground/src/noop/tlb.scala 44:26 86:30]
  wire  _GEN_139 = io_flush | flush_r ? _GEN_122 : valid_9; // @[playground/src/noop/tlb.scala 44:26 86:30]
  wire  _GEN_140 = io_flush | flush_r ? _GEN_123 : valid_10; // @[playground/src/noop/tlb.scala 44:26 86:30]
  wire  _GEN_141 = io_flush | flush_r ? _GEN_124 : valid_11; // @[playground/src/noop/tlb.scala 44:26 86:30]
  wire  _GEN_142 = io_flush | flush_r ? _GEN_125 : valid_12; // @[playground/src/noop/tlb.scala 44:26 86:30]
  wire  _GEN_143 = io_flush | flush_r ? _GEN_126 : valid_13; // @[playground/src/noop/tlb.scala 44:26 86:30]
  wire  _GEN_144 = io_flush | flush_r ? _GEN_127 : valid_14; // @[playground/src/noop/tlb.scala 44:26 86:30]
  wire  _GEN_145 = io_flush | flush_r ? _GEN_128 : valid_15; // @[playground/src/noop/tlb.scala 44:26 86:30]
  wire  handshake = io_va2pa_vvalid & io_va2pa_ready; // @[playground/src/noop/tlb.scala 94:37]
  reg [1:0] m_type_r; // @[playground/src/noop/tlb.scala 95:27]
  wire [1:0] cur_m_type = handshake ? io_va2pa_m_type : m_type_r; // @[playground/src/noop/tlb.scala 96:25]
  wire  _ad_T = cur_m_type == 2'h3; // @[playground/src/noop/common.scala 243:20]
  wire [9:0] ad = cur_m_type == 2'h3 ? 10'hc0 : 10'h40; // @[playground/src/noop/common.scala 243:12]
  wire  _GEN_150 = io_va2pa_pvalid | io_va2pa_tlb_excep_en ? 1'h0 : out_valid_r; // @[playground/src/noop/tlb.scala 108:51 109:21 51:30]
  wire  _GEN_151 = io_va2pa_pvalid | io_va2pa_tlb_excep_en ? 1'h0 : out_excep_r_en; // @[playground/src/noop/tlb.scala 108:51 110:24 53:30]
  wire  dc_hand = io_dcacheRW_ready & io_dcacheRW_dc_mode != 5'h0; // @[playground/src/noop/tlb.scala 122:37]
  wire [24:0] _tlb_high_legal_T_2 = io_va2pa_vaddr[38] ? 25'h1ffffff : 25'h0; // @[playground/src/noop/tlb.scala 125:30]
  wire  tlb_high_legal = _tlb_high_legal_T_2 == io_va2pa_vaddr[63:39]; // @[playground/src/noop/tlb.scala 125:55]
  wire  _tlb_access_illegal_T_11 = cur_m_type == 2'h2 & ~(tlbMsg_tlbInfo[1] | io_mmuState_mstatus[19] & tlbMsg_tlbInfo[3
    ]); // @[playground/src/noop/tlb.scala 127:60]
  wire  _tlb_access_illegal_T_12 = cur_m_type == 2'h1 & ~tlbMsg_tlbInfo[3] | _tlb_access_illegal_T_11; // @[playground/src/noop/tlb.scala 126:89]
  wire  _tlb_access_illegal_T_16 = _ad_T & ~tlbMsg_tlbInfo[2]; // @[playground/src/noop/tlb.scala 128:57]
  wire  tlb_access_illegal = _tlb_access_illegal_T_12 | _tlb_access_illegal_T_16; // @[playground/src/noop/tlb.scala 127:152]
  wire [3:0] select = {select_prng_io_out_3,select_prng_io_out_2,select_prng_io_out_1,select_prng_io_out_0}; // @[src/main/scala/chisel3/util/random/PRNG.scala 95:17]
  reg [3:0] select_r; // @[playground/src/noop/tlb.scala 130:27]
  reg [7:0] offset; // @[playground/src/noop/tlb.scala 131:26]
  reg [1:0] level; // @[playground/src/noop/tlb.scala 132:26]
  reg  wpte_hs_r; // @[playground/src/noop/tlb.scala 134:28]
  wire [63:0] _out_excep_r_cause_T_1 = 2'h1 == io_va2pa_m_type ? 64'hc : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 81:58]
  wire [63:0] _out_excep_r_cause_T_3 = 2'h2 == io_va2pa_m_type ? 64'hd : _out_excep_r_cause_T_1; // @[src/main/scala/chisel3/util/Mux.scala 81:58]
  wire [63:0] _out_excep_r_cause_T_5 = 2'h3 == io_va2pa_m_type ? 64'hf : _out_excep_r_cause_T_3; // @[src/main/scala/chisel3/util/Mux.scala 81:58]
  wire [51:0] _paddr_mask_T_4 = 2'h0 == tlbMsg_tlbLevel ? 52'hfffffffffffff : 52'h0; // @[src/main/scala/chisel3/util/Mux.scala 81:58]
  wire [51:0] _paddr_mask_T_6 = 2'h1 == tlbMsg_tlbLevel ? 52'hffffffffffe00 : _paddr_mask_T_4; // @[src/main/scala/chisel3/util/Mux.scala 81:58]
  wire [51:0] _paddr_mask_T_8 = 2'h2 == tlbMsg_tlbLevel ? 52'hffffffffc0000 : _paddr_mask_T_6; // @[src/main/scala/chisel3/util/Mux.scala 81:58]
  wire [63:0] paddr_mask = {_paddr_mask_T_8,12'h0}; // @[playground/src/noop/tlb.scala 147:41]
  wire [31:0] _out_paddr_r_T = {tlbMsg_tlbPa, 12'h0}; // @[playground/src/noop/tlb.scala 148:93]
  wire [63:0] _out_paddr_r_T_1 = ~paddr_mask; // @[playground/src/noop/common.scala 201:19]
  wire [63:0] _out_paddr_r_T_2 = io_va2pa_vaddr & _out_paddr_r_T_1; // @[playground/src/noop/common.scala 201:17]
  wire [63:0] _GEN_3 = {{32'd0}, _out_paddr_r_T}; // @[playground/src/noop/common.scala 201:36]
  wire [63:0] _out_paddr_r_T_3 = _GEN_3 & paddr_mask; // @[playground/src/noop/common.scala 201:36]
  wire [63:0] _out_paddr_r_T_4 = _out_paddr_r_T_2 | _out_paddr_r_T_3; // @[playground/src/noop/common.scala 201:26]
  wire [9:0] _T_59 = ad & tlbMsg_tlbInfo; // @[playground/src/noop/tlb.scala 149:30]
  wire [9:0] _wpte_data_r_T = tlbMsg_tlbInfo | ad; // @[playground/src/noop/tlb.scala 153:84]
  wire [63:0] _wpte_data_r_T_1 = {34'h0,tlbMsg_tlbPa,_wpte_data_r_T}; // @[playground/src/noop/tlb.scala 153:43]
  wire [9:0] _GEN_152 = 4'h0 == tlbMsg_tlbIdx ? _wpte_data_r_T : info_0; // @[playground/src/noop/tlb.scala 154:{45,45} 41:26]
  wire [9:0] _GEN_153 = 4'h1 == tlbMsg_tlbIdx ? _wpte_data_r_T : info_1; // @[playground/src/noop/tlb.scala 154:{45,45} 41:26]
  wire [9:0] _GEN_154 = 4'h2 == tlbMsg_tlbIdx ? _wpte_data_r_T : info_2; // @[playground/src/noop/tlb.scala 154:{45,45} 41:26]
  wire [9:0] _GEN_155 = 4'h3 == tlbMsg_tlbIdx ? _wpte_data_r_T : info_3; // @[playground/src/noop/tlb.scala 154:{45,45} 41:26]
  wire [9:0] _GEN_156 = 4'h4 == tlbMsg_tlbIdx ? _wpte_data_r_T : info_4; // @[playground/src/noop/tlb.scala 154:{45,45} 41:26]
  wire [9:0] _GEN_157 = 4'h5 == tlbMsg_tlbIdx ? _wpte_data_r_T : info_5; // @[playground/src/noop/tlb.scala 154:{45,45} 41:26]
  wire [9:0] _GEN_158 = 4'h6 == tlbMsg_tlbIdx ? _wpte_data_r_T : info_6; // @[playground/src/noop/tlb.scala 154:{45,45} 41:26]
  wire [9:0] _GEN_159 = 4'h7 == tlbMsg_tlbIdx ? _wpte_data_r_T : info_7; // @[playground/src/noop/tlb.scala 154:{45,45} 41:26]
  wire [9:0] _GEN_160 = 4'h8 == tlbMsg_tlbIdx ? _wpte_data_r_T : info_8; // @[playground/src/noop/tlb.scala 154:{45,45} 41:26]
  wire [9:0] _GEN_161 = 4'h9 == tlbMsg_tlbIdx ? _wpte_data_r_T : info_9; // @[playground/src/noop/tlb.scala 154:{45,45} 41:26]
  wire [9:0] _GEN_162 = 4'ha == tlbMsg_tlbIdx ? _wpte_data_r_T : info_10; // @[playground/src/noop/tlb.scala 154:{45,45} 41:26]
  wire [9:0] _GEN_163 = 4'hb == tlbMsg_tlbIdx ? _wpte_data_r_T : info_11; // @[playground/src/noop/tlb.scala 154:{45,45} 41:26]
  wire [9:0] _GEN_164 = 4'hc == tlbMsg_tlbIdx ? _wpte_data_r_T : info_12; // @[playground/src/noop/tlb.scala 154:{45,45} 41:26]
  wire [9:0] _GEN_165 = 4'hd == tlbMsg_tlbIdx ? _wpte_data_r_T : info_13; // @[playground/src/noop/tlb.scala 154:{45,45} 41:26]
  wire [9:0] _GEN_166 = 4'he == tlbMsg_tlbIdx ? _wpte_data_r_T : info_14; // @[playground/src/noop/tlb.scala 154:{45,45} 41:26]
  wire [9:0] _GEN_167 = 4'hf == tlbMsg_tlbIdx ? _wpte_data_r_T : info_15; // @[playground/src/noop/tlb.scala 154:{45,45} 41:26]
  wire [1:0] _GEN_168 = _T_59 != ad & is_Sv39 ? 2'h3 : state; // @[playground/src/noop/tlb.scala 149:66 150:31 84:24]
  wire  _GEN_169 = _T_59 != ad & is_Sv39 ? 1'h0 : wpte_hs_r; // @[playground/src/noop/tlb.scala 134:28 149:66 151:35]
  wire [31:0] _GEN_170 = _T_59 != ad & is_Sv39 ? tlbMsg_tlbPteAddr : pte_addr_r; // @[playground/src/noop/tlb.scala 149:66 152:37 47:30]
  wire [63:0] _GEN_171 = _T_59 != ad & is_Sv39 ? _wpte_data_r_T_1 : wpte_data_r; // @[playground/src/noop/tlb.scala 149:66 153:37 48:30]
  wire [9:0] _GEN_172 = _T_59 != ad & is_Sv39 ? _GEN_152 : info_0; // @[playground/src/noop/tlb.scala 149:66 41:26]
  wire [9:0] _GEN_173 = _T_59 != ad & is_Sv39 ? _GEN_153 : info_1; // @[playground/src/noop/tlb.scala 149:66 41:26]
  wire [9:0] _GEN_174 = _T_59 != ad & is_Sv39 ? _GEN_154 : info_2; // @[playground/src/noop/tlb.scala 149:66 41:26]
  wire [9:0] _GEN_175 = _T_59 != ad & is_Sv39 ? _GEN_155 : info_3; // @[playground/src/noop/tlb.scala 149:66 41:26]
  wire [9:0] _GEN_176 = _T_59 != ad & is_Sv39 ? _GEN_156 : info_4; // @[playground/src/noop/tlb.scala 149:66 41:26]
  wire [9:0] _GEN_177 = _T_59 != ad & is_Sv39 ? _GEN_157 : info_5; // @[playground/src/noop/tlb.scala 149:66 41:26]
  wire [9:0] _GEN_178 = _T_59 != ad & is_Sv39 ? _GEN_158 : info_6; // @[playground/src/noop/tlb.scala 149:66 41:26]
  wire [9:0] _GEN_179 = _T_59 != ad & is_Sv39 ? _GEN_159 : info_7; // @[playground/src/noop/tlb.scala 149:66 41:26]
  wire [9:0] _GEN_180 = _T_59 != ad & is_Sv39 ? _GEN_160 : info_8; // @[playground/src/noop/tlb.scala 149:66 41:26]
  wire [9:0] _GEN_181 = _T_59 != ad & is_Sv39 ? _GEN_161 : info_9; // @[playground/src/noop/tlb.scala 149:66 41:26]
  wire [9:0] _GEN_182 = _T_59 != ad & is_Sv39 ? _GEN_162 : info_10; // @[playground/src/noop/tlb.scala 149:66 41:26]
  wire [9:0] _GEN_183 = _T_59 != ad & is_Sv39 ? _GEN_163 : info_11; // @[playground/src/noop/tlb.scala 149:66 41:26]
  wire [9:0] _GEN_184 = _T_59 != ad & is_Sv39 ? _GEN_164 : info_12; // @[playground/src/noop/tlb.scala 149:66 41:26]
  wire [9:0] _GEN_185 = _T_59 != ad & is_Sv39 ? _GEN_165 : info_13; // @[playground/src/noop/tlb.scala 149:66 41:26]
  wire [9:0] _GEN_186 = _T_59 != ad & is_Sv39 ? _GEN_166 : info_14; // @[playground/src/noop/tlb.scala 149:66 41:26]
  wire [9:0] _GEN_187 = _T_59 != ad & is_Sv39 ? _GEN_167 : info_15; // @[playground/src/noop/tlb.scala 149:66 41:26]
  wire [63:0] _pte_addr_r_T_1 = {{30'd0}, io_va2pa_vaddr[63:30]}; // @[playground/src/noop/tlb.scala 166:83]
  wire [55:0] _pte_addr_r_T_3 = {io_mmuState_satp[43:0],_pte_addr_r_T_1[8:0],3'h0}; // @[playground/src/noop/tlb.scala 166:42]
  wire  _GEN_188 = io_va2pa_vaddr[63:39] != _tlb_high_legal_T_2 | _GEN_151; // @[playground/src/noop/tlb.scala 162:81 164:40]
  wire [55:0] _GEN_189 = io_va2pa_vaddr[63:39] != _tlb_high_legal_T_2 ? {{24'd0}, pte_addr_r} : _pte_addr_r_T_3; // @[playground/src/noop/tlb.scala 162:81 47:30 166:36]
  wire [4:0] _GEN_190 = io_va2pa_vaddr[63:39] != _tlb_high_legal_T_2 ? 5'h0 : 5'h7; // @[playground/src/noop/tlb.scala 138:27 162:81 167:36]
  wire [7:0] _GEN_191 = io_va2pa_vaddr[63:39] != _tlb_high_legal_T_2 ? offset : 8'h1e; // @[playground/src/noop/tlb.scala 131:26 162:81 168:33]
  wire [1:0] _GEN_192 = io_va2pa_vaddr[63:39] != _tlb_high_legal_T_2 ? level : 2'h3; // @[playground/src/noop/tlb.scala 132:26 162:81 169:33]
  wire [1:0] _GEN_194 = ~tlbMsg_tlbHit ? 2'h1 : state; // @[playground/src/noop/tlb.scala 156:43 84:24]
  wire [3:0] _GEN_195 = ~tlbMsg_tlbHit ? select : select_r; // @[playground/src/noop/tlb.scala 130:27 156:43 158:32]
  wire [1:0] _GEN_196 = ~tlbMsg_tlbHit ? io_va2pa_m_type : m_type_r; // @[playground/src/noop/tlb.scala 156:43 159:32 95:27]
  wire [63:0] _GEN_197 = ~tlbMsg_tlbHit ? _out_excep_r_cause_T_5 : out_excep_r_cause; // @[playground/src/noop/tlb.scala 156:43 160:39 53:30]
  wire [63:0] _GEN_198 = ~tlbMsg_tlbHit ? io_va2pa_vaddr : out_excep_r_tval; // @[playground/src/noop/tlb.scala 156:43 161:39 53:30]
  wire  _GEN_199 = ~tlbMsg_tlbHit ? _GEN_188 : _GEN_151; // @[playground/src/noop/tlb.scala 156:43]
  wire [55:0] _GEN_200 = ~tlbMsg_tlbHit ? _GEN_189 : {{24'd0}, pte_addr_r}; // @[playground/src/noop/tlb.scala 156:43 47:30]
  wire [4:0] _GEN_201 = ~tlbMsg_tlbHit ? _GEN_190 : 5'h0; // @[playground/src/noop/tlb.scala 138:27 156:43]
  wire [7:0] _GEN_202 = ~tlbMsg_tlbHit ? _GEN_191 : offset; // @[playground/src/noop/tlb.scala 131:26 156:43]
  wire [1:0] _GEN_203 = ~tlbMsg_tlbHit ? _GEN_192 : level; // @[playground/src/noop/tlb.scala 132:26 156:43]
  wire  _GEN_204 = tlbMsg_tlbHit | _GEN_150; // @[playground/src/noop/tlb.scala 144:42 145:33]
  wire [63:0] _GEN_205 = tlbMsg_tlbHit ? _out_paddr_r_T_4 : {{32'd0}, out_paddr_r}; // @[playground/src/noop/tlb.scala 144:42 148:33 52:30]
  wire [1:0] _GEN_206 = tlbMsg_tlbHit ? _GEN_168 : _GEN_194; // @[playground/src/noop/tlb.scala 144:42]
  wire  _GEN_207 = tlbMsg_tlbHit ? _GEN_169 : wpte_hs_r; // @[playground/src/noop/tlb.scala 134:28 144:42]
  wire [55:0] _GEN_208 = tlbMsg_tlbHit ? {{24'd0}, _GEN_170} : _GEN_200; // @[playground/src/noop/tlb.scala 144:42]
  wire [63:0] _GEN_209 = tlbMsg_tlbHit ? _GEN_171 : wpte_data_r; // @[playground/src/noop/tlb.scala 144:42 48:30]
  wire [9:0] _GEN_210 = tlbMsg_tlbHit ? _GEN_172 : info_0; // @[playground/src/noop/tlb.scala 144:42 41:26]
  wire [9:0] _GEN_211 = tlbMsg_tlbHit ? _GEN_173 : info_1; // @[playground/src/noop/tlb.scala 144:42 41:26]
  wire [9:0] _GEN_212 = tlbMsg_tlbHit ? _GEN_174 : info_2; // @[playground/src/noop/tlb.scala 144:42 41:26]
  wire [9:0] _GEN_213 = tlbMsg_tlbHit ? _GEN_175 : info_3; // @[playground/src/noop/tlb.scala 144:42 41:26]
  wire [9:0] _GEN_214 = tlbMsg_tlbHit ? _GEN_176 : info_4; // @[playground/src/noop/tlb.scala 144:42 41:26]
  wire [9:0] _GEN_215 = tlbMsg_tlbHit ? _GEN_177 : info_5; // @[playground/src/noop/tlb.scala 144:42 41:26]
  wire [9:0] _GEN_216 = tlbMsg_tlbHit ? _GEN_178 : info_6; // @[playground/src/noop/tlb.scala 144:42 41:26]
  wire [9:0] _GEN_217 = tlbMsg_tlbHit ? _GEN_179 : info_7; // @[playground/src/noop/tlb.scala 144:42 41:26]
  wire [9:0] _GEN_218 = tlbMsg_tlbHit ? _GEN_180 : info_8; // @[playground/src/noop/tlb.scala 144:42 41:26]
  wire [9:0] _GEN_219 = tlbMsg_tlbHit ? _GEN_181 : info_9; // @[playground/src/noop/tlb.scala 144:42 41:26]
  wire [9:0] _GEN_220 = tlbMsg_tlbHit ? _GEN_182 : info_10; // @[playground/src/noop/tlb.scala 144:42 41:26]
  wire [9:0] _GEN_221 = tlbMsg_tlbHit ? _GEN_183 : info_11; // @[playground/src/noop/tlb.scala 144:42 41:26]
  wire [9:0] _GEN_222 = tlbMsg_tlbHit ? _GEN_184 : info_12; // @[playground/src/noop/tlb.scala 144:42 41:26]
  wire [9:0] _GEN_223 = tlbMsg_tlbHit ? _GEN_185 : info_13; // @[playground/src/noop/tlb.scala 144:42 41:26]
  wire [9:0] _GEN_224 = tlbMsg_tlbHit ? _GEN_186 : info_14; // @[playground/src/noop/tlb.scala 144:42 41:26]
  wire [9:0] _GEN_225 = tlbMsg_tlbHit ? _GEN_187 : info_15; // @[playground/src/noop/tlb.scala 144:42 41:26]
  wire [3:0] _GEN_226 = tlbMsg_tlbHit ? select_r : _GEN_195; // @[playground/src/noop/tlb.scala 130:27 144:42]
  wire [1:0] _GEN_227 = tlbMsg_tlbHit ? m_type_r : _GEN_196; // @[playground/src/noop/tlb.scala 144:42 95:27]
  wire [63:0] _GEN_228 = tlbMsg_tlbHit ? out_excep_r_cause : _GEN_197; // @[playground/src/noop/tlb.scala 144:42 53:30]
  wire [63:0] _GEN_229 = tlbMsg_tlbHit ? out_excep_r_tval : _GEN_198; // @[playground/src/noop/tlb.scala 144:42 53:30]
  wire  _GEN_230 = tlbMsg_tlbHit ? _GEN_151 : _GEN_199; // @[playground/src/noop/tlb.scala 144:42]
  wire [4:0] _GEN_231 = tlbMsg_tlbHit ? 5'h0 : _GEN_201; // @[playground/src/noop/tlb.scala 138:27 144:42]
  wire [7:0] _GEN_232 = tlbMsg_tlbHit ? offset : _GEN_202; // @[playground/src/noop/tlb.scala 131:26 144:42]
  wire [1:0] _GEN_233 = tlbMsg_tlbHit ? level : _GEN_203; // @[playground/src/noop/tlb.scala 132:26 144:42]
  wire  _GEN_234 = ~tlb_high_legal | tlbMsg_tlbHit & tlb_access_illegal | _GEN_230; // @[playground/src/noop/tlb.scala 140:85 141:36]
  wire [63:0] _GEN_235 = ~tlb_high_legal | tlbMsg_tlbHit & tlb_access_illegal ? _out_excep_r_cause_T_5 : _GEN_228; // @[playground/src/noop/tlb.scala 140:85 142:39]
  wire [63:0] _GEN_236 = ~tlb_high_legal | tlbMsg_tlbHit & tlb_access_illegal ? io_va2pa_vaddr : _GEN_229; // @[playground/src/noop/tlb.scala 140:85 143:39]
  wire  _GEN_237 = ~tlb_high_legal | tlbMsg_tlbHit & tlb_access_illegal ? _GEN_150 : _GEN_204; // @[playground/src/noop/tlb.scala 140:85]
  wire [63:0] _GEN_238 = ~tlb_high_legal | tlbMsg_tlbHit & tlb_access_illegal ? {{32'd0}, out_paddr_r} : _GEN_205; // @[playground/src/noop/tlb.scala 140:85 52:30]
  wire [1:0] _GEN_239 = ~tlb_high_legal | tlbMsg_tlbHit & tlb_access_illegal ? state : _GEN_206; // @[playground/src/noop/tlb.scala 140:85 84:24]
  wire  _GEN_240 = ~tlb_high_legal | tlbMsg_tlbHit & tlb_access_illegal ? wpte_hs_r : _GEN_207; // @[playground/src/noop/tlb.scala 134:28 140:85]
  wire [55:0] _GEN_241 = ~tlb_high_legal | tlbMsg_tlbHit & tlb_access_illegal ? {{24'd0}, pte_addr_r} : _GEN_208; // @[playground/src/noop/tlb.scala 140:85 47:30]
  wire [63:0] _GEN_242 = ~tlb_high_legal | tlbMsg_tlbHit & tlb_access_illegal ? wpte_data_r : _GEN_209; // @[playground/src/noop/tlb.scala 140:85 48:30]
  wire [9:0] _GEN_243 = ~tlb_high_legal | tlbMsg_tlbHit & tlb_access_illegal ? info_0 : _GEN_210; // @[playground/src/noop/tlb.scala 140:85 41:26]
  wire [9:0] _GEN_244 = ~tlb_high_legal | tlbMsg_tlbHit & tlb_access_illegal ? info_1 : _GEN_211; // @[playground/src/noop/tlb.scala 140:85 41:26]
  wire [9:0] _GEN_245 = ~tlb_high_legal | tlbMsg_tlbHit & tlb_access_illegal ? info_2 : _GEN_212; // @[playground/src/noop/tlb.scala 140:85 41:26]
  wire [9:0] _GEN_246 = ~tlb_high_legal | tlbMsg_tlbHit & tlb_access_illegal ? info_3 : _GEN_213; // @[playground/src/noop/tlb.scala 140:85 41:26]
  wire [9:0] _GEN_247 = ~tlb_high_legal | tlbMsg_tlbHit & tlb_access_illegal ? info_4 : _GEN_214; // @[playground/src/noop/tlb.scala 140:85 41:26]
  wire [9:0] _GEN_248 = ~tlb_high_legal | tlbMsg_tlbHit & tlb_access_illegal ? info_5 : _GEN_215; // @[playground/src/noop/tlb.scala 140:85 41:26]
  wire [9:0] _GEN_249 = ~tlb_high_legal | tlbMsg_tlbHit & tlb_access_illegal ? info_6 : _GEN_216; // @[playground/src/noop/tlb.scala 140:85 41:26]
  wire [9:0] _GEN_250 = ~tlb_high_legal | tlbMsg_tlbHit & tlb_access_illegal ? info_7 : _GEN_217; // @[playground/src/noop/tlb.scala 140:85 41:26]
  wire [9:0] _GEN_251 = ~tlb_high_legal | tlbMsg_tlbHit & tlb_access_illegal ? info_8 : _GEN_218; // @[playground/src/noop/tlb.scala 140:85 41:26]
  wire [9:0] _GEN_252 = ~tlb_high_legal | tlbMsg_tlbHit & tlb_access_illegal ? info_9 : _GEN_219; // @[playground/src/noop/tlb.scala 140:85 41:26]
  wire [9:0] _GEN_253 = ~tlb_high_legal | tlbMsg_tlbHit & tlb_access_illegal ? info_10 : _GEN_220; // @[playground/src/noop/tlb.scala 140:85 41:26]
  wire [9:0] _GEN_254 = ~tlb_high_legal | tlbMsg_tlbHit & tlb_access_illegal ? info_11 : _GEN_221; // @[playground/src/noop/tlb.scala 140:85 41:26]
  wire [9:0] _GEN_255 = ~tlb_high_legal | tlbMsg_tlbHit & tlb_access_illegal ? info_12 : _GEN_222; // @[playground/src/noop/tlb.scala 140:85 41:26]
  wire [9:0] _GEN_256 = ~tlb_high_legal | tlbMsg_tlbHit & tlb_access_illegal ? info_13 : _GEN_223; // @[playground/src/noop/tlb.scala 140:85 41:26]
  wire [9:0] _GEN_257 = ~tlb_high_legal | tlbMsg_tlbHit & tlb_access_illegal ? info_14 : _GEN_224; // @[playground/src/noop/tlb.scala 140:85 41:26]
  wire [9:0] _GEN_258 = ~tlb_high_legal | tlbMsg_tlbHit & tlb_access_illegal ? info_15 : _GEN_225; // @[playground/src/noop/tlb.scala 140:85 41:26]
  wire [3:0] _GEN_259 = ~tlb_high_legal | tlbMsg_tlbHit & tlb_access_illegal ? select_r : _GEN_226; // @[playground/src/noop/tlb.scala 130:27 140:85]
  wire [1:0] _GEN_260 = ~tlb_high_legal | tlbMsg_tlbHit & tlb_access_illegal ? m_type_r : _GEN_227; // @[playground/src/noop/tlb.scala 140:85 95:27]
  wire [4:0] _GEN_261 = ~tlb_high_legal | tlbMsg_tlbHit & tlb_access_illegal ? 5'h0 : _GEN_231; // @[playground/src/noop/tlb.scala 138:27 140:85]
  wire [7:0] _GEN_262 = ~tlb_high_legal | tlbMsg_tlbHit & tlb_access_illegal ? offset : _GEN_232; // @[playground/src/noop/tlb.scala 131:26 140:85]
  wire [1:0] _GEN_263 = ~tlb_high_legal | tlbMsg_tlbHit & tlb_access_illegal ? level : _GEN_233; // @[playground/src/noop/tlb.scala 132:26 140:85]
  wire [63:0] _GEN_268 = ~handshake ? {{32'd0}, out_paddr_r} : _GEN_238; // @[playground/src/noop/tlb.scala 139:33 52:30]
  wire [55:0] _GEN_271 = ~handshake ? {{24'd0}, pte_addr_r} : _GEN_241; // @[playground/src/noop/tlb.scala 139:33 47:30]
  wire [4:0] _dc_mode_r_T = wpte_hs_r ? 5'h0 : 5'hb; // @[playground/src/noop/tlb.scala 175:33]
  wire [4:0] _GEN_294 = io_dcacheRW_ready ? 5'h0 : _dc_mode_r_T; // @[playground/src/noop/tlb.scala 175:27 176:40 177:31]
  wire  _GEN_295 = io_dcacheRW_ready | wpte_hs_r; // @[playground/src/noop/tlb.scala 134:28 176:40 178:31]
  wire [1:0] _GEN_296 = io_dcacheRW_rvalid ? 2'h0 : state; // @[playground/src/noop/tlb.scala 180:41 181:27 84:24]
  wire [7:0] _offset_T_1 = offset - 8'h9; // @[playground/src/noop/tlb.scala 187:39]
  wire [1:0] _level_T_1 = level - 2'h1; // @[playground/src/noop/tlb.scala 188:38]
  wire [4:0] _GEN_297 = dc_hand ? 5'h0 : dc_mode_r; // @[playground/src/noop/tlb.scala 185:30 186:31 49:30]
  wire [7:0] _GEN_298 = dc_hand ? _offset_T_1 : offset; // @[playground/src/noop/tlb.scala 131:26 185:30 187:29]
  wire [1:0] _GEN_299 = dc_hand ? _level_T_1 : level; // @[playground/src/noop/tlb.scala 132:26 185:30 188:29]
  wire [63:0] _T_73 = io_dcacheRW_rdata & 64'hf; // @[playground/src/noop/tlb.scala 191:31]
  wire [63:0] _T_77 = io_dcacheRW_rdata & 64'hd0; // @[playground/src/noop/tlb.scala 192:35]
  wire [63:0] _pte_addr_r_T_5 = pre_addr >> offset; // @[playground/src/noop/tlb.scala 196:69]
  wire [55:0] _pte_addr_r_T_7 = {io_dcacheRW_rdata[53:10],_pte_addr_r_T_5[8:0],3'h0}; // @[playground/src/noop/tlb.scala 196:46]
  wire [1:0] _GEN_300 = _T_77 != 64'h0 ? 2'h0 : state; // @[playground/src/noop/tlb.scala 192:70 193:35 84:24]
  wire  _GEN_301 = _T_77 != 64'h0 | _GEN_151; // @[playground/src/noop/tlb.scala 192:70 194:44]
  wire [55:0] _GEN_302 = _T_77 != 64'h0 ? {{24'd0}, pte_addr_r} : _pte_addr_r_T_7; // @[playground/src/noop/tlb.scala 192:70 47:30 196:40]
  wire [4:0] _GEN_303 = _T_77 != 64'h0 ? _GEN_297 : 5'h7; // @[playground/src/noop/tlb.scala 192:70 197:40]
  wire  _T_83 = out_excep_r_cause == 64'hc; // @[playground/src/noop/tlb.scala 199:133]
  wire  _T_87 = io_dcacheRW_rdata[4] ? io_mmuState_priv == 2'h1 & (~io_mmuState_mstatus[18] | out_excep_r_cause == 64'hc
    ) : io_mmuState_priv == 2'h0; // @[playground/src/noop/tlb.scala 199:35]
  wire  _T_106 = out_excep_r_cause == 64'hd & ~(io_dcacheRW_rdata[1] | io_mmuState_mstatus[19] & io_dcacheRW_rdata[3]); // @[playground/src/noop/tlb.scala 208:82]
  wire  _T_107 = _T_83 & ~io_dcacheRW_rdata[3] | _T_106; // @[playground/src/noop/tlb.scala 207:102]
  wire  _T_111 = out_excep_r_cause == 64'hf & ~io_dcacheRW_rdata[2]; // @[playground/src/noop/tlb.scala 209:79]
  wire  _T_112 = _T_107 | _T_111; // @[playground/src/noop/tlb.scala 208:152]
  wire [51:0] _ppn_mask_T_4 = 2'h0 == level ? 52'hfffffffffffff : 52'h0; // @[src/main/scala/chisel3/util/Mux.scala 81:58]
  wire [51:0] _ppn_mask_T_6 = 2'h1 == level ? 52'hffffffffffe00 : _ppn_mask_T_4; // @[src/main/scala/chisel3/util/Mux.scala 81:58]
  wire [51:0] ppn_mask = 2'h2 == level ? 52'hffffffffc0000 : _ppn_mask_T_6; // @[src/main/scala/chisel3/util/Mux.scala 81:58]
  wire [51:0] _tag_T_1 = pre_addr[63:12] & ppn_mask; // @[playground/src/noop/tlb.scala 220:78]
  wire [51:0] _GEN_304 = 4'h0 == select_r ? _tag_T_1 : tag_0; // @[playground/src/noop/tlb.scala 220:{39,39} 39:26]
  wire [51:0] _GEN_305 = 4'h1 == select_r ? _tag_T_1 : tag_1; // @[playground/src/noop/tlb.scala 220:{39,39} 39:26]
  wire [51:0] _GEN_306 = 4'h2 == select_r ? _tag_T_1 : tag_2; // @[playground/src/noop/tlb.scala 220:{39,39} 39:26]
  wire [51:0] _GEN_307 = 4'h3 == select_r ? _tag_T_1 : tag_3; // @[playground/src/noop/tlb.scala 220:{39,39} 39:26]
  wire [51:0] _GEN_308 = 4'h4 == select_r ? _tag_T_1 : tag_4; // @[playground/src/noop/tlb.scala 220:{39,39} 39:26]
  wire [51:0] _GEN_309 = 4'h5 == select_r ? _tag_T_1 : tag_5; // @[playground/src/noop/tlb.scala 220:{39,39} 39:26]
  wire [51:0] _GEN_310 = 4'h6 == select_r ? _tag_T_1 : tag_6; // @[playground/src/noop/tlb.scala 220:{39,39} 39:26]
  wire [51:0] _GEN_311 = 4'h7 == select_r ? _tag_T_1 : tag_7; // @[playground/src/noop/tlb.scala 220:{39,39} 39:26]
  wire [51:0] _GEN_312 = 4'h8 == select_r ? _tag_T_1 : tag_8; // @[playground/src/noop/tlb.scala 220:{39,39} 39:26]
  wire [51:0] _GEN_313 = 4'h9 == select_r ? _tag_T_1 : tag_9; // @[playground/src/noop/tlb.scala 220:{39,39} 39:26]
  wire [51:0] _GEN_314 = 4'ha == select_r ? _tag_T_1 : tag_10; // @[playground/src/noop/tlb.scala 220:{39,39} 39:26]
  wire [51:0] _GEN_315 = 4'hb == select_r ? _tag_T_1 : tag_11; // @[playground/src/noop/tlb.scala 220:{39,39} 39:26]
  wire [51:0] _GEN_316 = 4'hc == select_r ? _tag_T_1 : tag_12; // @[playground/src/noop/tlb.scala 220:{39,39} 39:26]
  wire [51:0] _GEN_317 = 4'hd == select_r ? _tag_T_1 : tag_13; // @[playground/src/noop/tlb.scala 220:{39,39} 39:26]
  wire [51:0] _GEN_318 = 4'he == select_r ? _tag_T_1 : tag_14; // @[playground/src/noop/tlb.scala 220:{39,39} 39:26]
  wire [51:0] _GEN_319 = 4'hf == select_r ? _tag_T_1 : tag_15; // @[playground/src/noop/tlb.scala 220:{39,39} 39:26]
  wire  _GEN_320 = 4'h0 == select_r | _GEN_130; // @[playground/src/noop/tlb.scala 221:{41,41}]
  wire  _GEN_321 = 4'h1 == select_r | _GEN_131; // @[playground/src/noop/tlb.scala 221:{41,41}]
  wire  _GEN_322 = 4'h2 == select_r | _GEN_132; // @[playground/src/noop/tlb.scala 221:{41,41}]
  wire  _GEN_323 = 4'h3 == select_r | _GEN_133; // @[playground/src/noop/tlb.scala 221:{41,41}]
  wire  _GEN_324 = 4'h4 == select_r | _GEN_134; // @[playground/src/noop/tlb.scala 221:{41,41}]
  wire  _GEN_325 = 4'h5 == select_r | _GEN_135; // @[playground/src/noop/tlb.scala 221:{41,41}]
  wire  _GEN_326 = 4'h6 == select_r | _GEN_136; // @[playground/src/noop/tlb.scala 221:{41,41}]
  wire  _GEN_327 = 4'h7 == select_r | _GEN_137; // @[playground/src/noop/tlb.scala 221:{41,41}]
  wire  _GEN_328 = 4'h8 == select_r | _GEN_138; // @[playground/src/noop/tlb.scala 221:{41,41}]
  wire  _GEN_329 = 4'h9 == select_r | _GEN_139; // @[playground/src/noop/tlb.scala 221:{41,41}]
  wire  _GEN_330 = 4'ha == select_r | _GEN_140; // @[playground/src/noop/tlb.scala 221:{41,41}]
  wire  _GEN_331 = 4'hb == select_r | _GEN_141; // @[playground/src/noop/tlb.scala 221:{41,41}]
  wire  _GEN_332 = 4'hc == select_r | _GEN_142; // @[playground/src/noop/tlb.scala 221:{41,41}]
  wire  _GEN_333 = 4'hd == select_r | _GEN_143; // @[playground/src/noop/tlb.scala 221:{41,41}]
  wire  _GEN_334 = 4'he == select_r | _GEN_144; // @[playground/src/noop/tlb.scala 221:{41,41}]
  wire  _GEN_335 = 4'hf == select_r | _GEN_145; // @[playground/src/noop/tlb.scala 221:{41,41}]
  wire [51:0] _GEN_1417 = {{32'd0}, io_dcacheRW_rdata[29:10]}; // @[playground/src/noop/tlb.scala 222:53]
  wire [51:0] update_pa = _GEN_1417 & ppn_mask; // @[playground/src/noop/tlb.scala 222:53]
  wire [19:0] _GEN_336 = 4'h0 == select_r ? update_pa[19:0] : paddr_0; // @[playground/src/noop/tlb.scala 223:{41,41} 40:26]
  wire [19:0] _GEN_337 = 4'h1 == select_r ? update_pa[19:0] : paddr_1; // @[playground/src/noop/tlb.scala 223:{41,41} 40:26]
  wire [19:0] _GEN_338 = 4'h2 == select_r ? update_pa[19:0] : paddr_2; // @[playground/src/noop/tlb.scala 223:{41,41} 40:26]
  wire [19:0] _GEN_339 = 4'h3 == select_r ? update_pa[19:0] : paddr_3; // @[playground/src/noop/tlb.scala 223:{41,41} 40:26]
  wire [19:0] _GEN_340 = 4'h4 == select_r ? update_pa[19:0] : paddr_4; // @[playground/src/noop/tlb.scala 223:{41,41} 40:26]
  wire [19:0] _GEN_341 = 4'h5 == select_r ? update_pa[19:0] : paddr_5; // @[playground/src/noop/tlb.scala 223:{41,41} 40:26]
  wire [19:0] _GEN_342 = 4'h6 == select_r ? update_pa[19:0] : paddr_6; // @[playground/src/noop/tlb.scala 223:{41,41} 40:26]
  wire [19:0] _GEN_343 = 4'h7 == select_r ? update_pa[19:0] : paddr_7; // @[playground/src/noop/tlb.scala 223:{41,41} 40:26]
  wire [19:0] _GEN_344 = 4'h8 == select_r ? update_pa[19:0] : paddr_8; // @[playground/src/noop/tlb.scala 223:{41,41} 40:26]
  wire [19:0] _GEN_345 = 4'h9 == select_r ? update_pa[19:0] : paddr_9; // @[playground/src/noop/tlb.scala 223:{41,41} 40:26]
  wire [19:0] _GEN_346 = 4'ha == select_r ? update_pa[19:0] : paddr_10; // @[playground/src/noop/tlb.scala 223:{41,41} 40:26]
  wire [19:0] _GEN_347 = 4'hb == select_r ? update_pa[19:0] : paddr_11; // @[playground/src/noop/tlb.scala 223:{41,41} 40:26]
  wire [19:0] _GEN_348 = 4'hc == select_r ? update_pa[19:0] : paddr_12; // @[playground/src/noop/tlb.scala 223:{41,41} 40:26]
  wire [19:0] _GEN_349 = 4'hd == select_r ? update_pa[19:0] : paddr_13; // @[playground/src/noop/tlb.scala 223:{41,41} 40:26]
  wire [19:0] _GEN_350 = 4'he == select_r ? update_pa[19:0] : paddr_14; // @[playground/src/noop/tlb.scala 223:{41,41} 40:26]
  wire [19:0] _GEN_351 = 4'hf == select_r ? update_pa[19:0] : paddr_15; // @[playground/src/noop/tlb.scala 223:{41,41} 40:26]
  wire [31:0] _GEN_352 = 4'h0 == select_r ? pte_addr_r : pte_addr_0; // @[playground/src/noop/tlb.scala 224:{44,44} 42:30]
  wire [31:0] _GEN_353 = 4'h1 == select_r ? pte_addr_r : pte_addr_1; // @[playground/src/noop/tlb.scala 224:{44,44} 42:30]
  wire [31:0] _GEN_354 = 4'h2 == select_r ? pte_addr_r : pte_addr_2; // @[playground/src/noop/tlb.scala 224:{44,44} 42:30]
  wire [31:0] _GEN_355 = 4'h3 == select_r ? pte_addr_r : pte_addr_3; // @[playground/src/noop/tlb.scala 224:{44,44} 42:30]
  wire [31:0] _GEN_356 = 4'h4 == select_r ? pte_addr_r : pte_addr_4; // @[playground/src/noop/tlb.scala 224:{44,44} 42:30]
  wire [31:0] _GEN_357 = 4'h5 == select_r ? pte_addr_r : pte_addr_5; // @[playground/src/noop/tlb.scala 224:{44,44} 42:30]
  wire [31:0] _GEN_358 = 4'h6 == select_r ? pte_addr_r : pte_addr_6; // @[playground/src/noop/tlb.scala 224:{44,44} 42:30]
  wire [31:0] _GEN_359 = 4'h7 == select_r ? pte_addr_r : pte_addr_7; // @[playground/src/noop/tlb.scala 224:{44,44} 42:30]
  wire [31:0] _GEN_360 = 4'h8 == select_r ? pte_addr_r : pte_addr_8; // @[playground/src/noop/tlb.scala 224:{44,44} 42:30]
  wire [31:0] _GEN_361 = 4'h9 == select_r ? pte_addr_r : pte_addr_9; // @[playground/src/noop/tlb.scala 224:{44,44} 42:30]
  wire [31:0] _GEN_362 = 4'ha == select_r ? pte_addr_r : pte_addr_10; // @[playground/src/noop/tlb.scala 224:{44,44} 42:30]
  wire [31:0] _GEN_363 = 4'hb == select_r ? pte_addr_r : pte_addr_11; // @[playground/src/noop/tlb.scala 224:{44,44} 42:30]
  wire [31:0] _GEN_364 = 4'hc == select_r ? pte_addr_r : pte_addr_12; // @[playground/src/noop/tlb.scala 224:{44,44} 42:30]
  wire [31:0] _GEN_365 = 4'hd == select_r ? pte_addr_r : pte_addr_13; // @[playground/src/noop/tlb.scala 224:{44,44} 42:30]
  wire [31:0] _GEN_366 = 4'he == select_r ? pte_addr_r : pte_addr_14; // @[playground/src/noop/tlb.scala 224:{44,44} 42:30]
  wire [31:0] _GEN_367 = 4'hf == select_r ? pte_addr_r : pte_addr_15; // @[playground/src/noop/tlb.scala 224:{44,44} 42:30]
  wire [1:0] _GEN_368 = 4'h0 == select_r ? level : pte_level_0; // @[playground/src/noop/tlb.scala 225:{45,45} 43:30]
  wire [1:0] _GEN_369 = 4'h1 == select_r ? level : pte_level_1; // @[playground/src/noop/tlb.scala 225:{45,45} 43:30]
  wire [1:0] _GEN_370 = 4'h2 == select_r ? level : pte_level_2; // @[playground/src/noop/tlb.scala 225:{45,45} 43:30]
  wire [1:0] _GEN_371 = 4'h3 == select_r ? level : pte_level_3; // @[playground/src/noop/tlb.scala 225:{45,45} 43:30]
  wire [1:0] _GEN_372 = 4'h4 == select_r ? level : pte_level_4; // @[playground/src/noop/tlb.scala 225:{45,45} 43:30]
  wire [1:0] _GEN_373 = 4'h5 == select_r ? level : pte_level_5; // @[playground/src/noop/tlb.scala 225:{45,45} 43:30]
  wire [1:0] _GEN_374 = 4'h6 == select_r ? level : pte_level_6; // @[playground/src/noop/tlb.scala 225:{45,45} 43:30]
  wire [1:0] _GEN_375 = 4'h7 == select_r ? level : pte_level_7; // @[playground/src/noop/tlb.scala 225:{45,45} 43:30]
  wire [1:0] _GEN_376 = 4'h8 == select_r ? level : pte_level_8; // @[playground/src/noop/tlb.scala 225:{45,45} 43:30]
  wire [1:0] _GEN_377 = 4'h9 == select_r ? level : pte_level_9; // @[playground/src/noop/tlb.scala 225:{45,45} 43:30]
  wire [1:0] _GEN_378 = 4'ha == select_r ? level : pte_level_10; // @[playground/src/noop/tlb.scala 225:{45,45} 43:30]
  wire [1:0] _GEN_379 = 4'hb == select_r ? level : pte_level_11; // @[playground/src/noop/tlb.scala 225:{45,45} 43:30]
  wire [1:0] _GEN_380 = 4'hc == select_r ? level : pte_level_12; // @[playground/src/noop/tlb.scala 225:{45,45} 43:30]
  wire [1:0] _GEN_381 = 4'hd == select_r ? level : pte_level_13; // @[playground/src/noop/tlb.scala 225:{45,45} 43:30]
  wire [1:0] _GEN_382 = 4'he == select_r ? level : pte_level_14; // @[playground/src/noop/tlb.scala 225:{45,45} 43:30]
  wire [1:0] _GEN_383 = 4'hf == select_r ? level : pte_level_15; // @[playground/src/noop/tlb.scala 225:{45,45} 43:30]
  wire [9:0] _GEN_384 = 4'h0 == select_r ? io_dcacheRW_rdata[9:0] : info_0; // @[playground/src/noop/tlb.scala 226:{40,40} 41:26]
  wire [9:0] _GEN_385 = 4'h1 == select_r ? io_dcacheRW_rdata[9:0] : info_1; // @[playground/src/noop/tlb.scala 226:{40,40} 41:26]
  wire [9:0] _GEN_386 = 4'h2 == select_r ? io_dcacheRW_rdata[9:0] : info_2; // @[playground/src/noop/tlb.scala 226:{40,40} 41:26]
  wire [9:0] _GEN_387 = 4'h3 == select_r ? io_dcacheRW_rdata[9:0] : info_3; // @[playground/src/noop/tlb.scala 226:{40,40} 41:26]
  wire [9:0] _GEN_388 = 4'h4 == select_r ? io_dcacheRW_rdata[9:0] : info_4; // @[playground/src/noop/tlb.scala 226:{40,40} 41:26]
  wire [9:0] _GEN_389 = 4'h5 == select_r ? io_dcacheRW_rdata[9:0] : info_5; // @[playground/src/noop/tlb.scala 226:{40,40} 41:26]
  wire [9:0] _GEN_390 = 4'h6 == select_r ? io_dcacheRW_rdata[9:0] : info_6; // @[playground/src/noop/tlb.scala 226:{40,40} 41:26]
  wire [9:0] _GEN_391 = 4'h7 == select_r ? io_dcacheRW_rdata[9:0] : info_7; // @[playground/src/noop/tlb.scala 226:{40,40} 41:26]
  wire [9:0] _GEN_392 = 4'h8 == select_r ? io_dcacheRW_rdata[9:0] : info_8; // @[playground/src/noop/tlb.scala 226:{40,40} 41:26]
  wire [9:0] _GEN_393 = 4'h9 == select_r ? io_dcacheRW_rdata[9:0] : info_9; // @[playground/src/noop/tlb.scala 226:{40,40} 41:26]
  wire [9:0] _GEN_394 = 4'ha == select_r ? io_dcacheRW_rdata[9:0] : info_10; // @[playground/src/noop/tlb.scala 226:{40,40} 41:26]
  wire [9:0] _GEN_395 = 4'hb == select_r ? io_dcacheRW_rdata[9:0] : info_11; // @[playground/src/noop/tlb.scala 226:{40,40} 41:26]
  wire [9:0] _GEN_396 = 4'hc == select_r ? io_dcacheRW_rdata[9:0] : info_12; // @[playground/src/noop/tlb.scala 226:{40,40} 41:26]
  wire [9:0] _GEN_397 = 4'hd == select_r ? io_dcacheRW_rdata[9:0] : info_13; // @[playground/src/noop/tlb.scala 226:{40,40} 41:26]
  wire [9:0] _GEN_398 = 4'he == select_r ? io_dcacheRW_rdata[9:0] : info_14; // @[playground/src/noop/tlb.scala 226:{40,40} 41:26]
  wire [9:0] _GEN_399 = 4'hf == select_r ? io_dcacheRW_rdata[9:0] : info_15; // @[playground/src/noop/tlb.scala 226:{40,40} 41:26]
  wire  _GEN_401 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     | _GEN_151; // @[playground/src/noop/tlb.scala 213:117 216:40]
  wire [51:0] _GEN_402 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? tag_0 : _GEN_304; // @[playground/src/noop/tlb.scala 213:117 39:26]
  wire [51:0] _GEN_403 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? tag_1 : _GEN_305; // @[playground/src/noop/tlb.scala 213:117 39:26]
  wire [51:0] _GEN_404 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? tag_2 : _GEN_306; // @[playground/src/noop/tlb.scala 213:117 39:26]
  wire [51:0] _GEN_405 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? tag_3 : _GEN_307; // @[playground/src/noop/tlb.scala 213:117 39:26]
  wire [51:0] _GEN_406 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? tag_4 : _GEN_308; // @[playground/src/noop/tlb.scala 213:117 39:26]
  wire [51:0] _GEN_407 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? tag_5 : _GEN_309; // @[playground/src/noop/tlb.scala 213:117 39:26]
  wire [51:0] _GEN_408 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? tag_6 : _GEN_310; // @[playground/src/noop/tlb.scala 213:117 39:26]
  wire [51:0] _GEN_409 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? tag_7 : _GEN_311; // @[playground/src/noop/tlb.scala 213:117 39:26]
  wire [51:0] _GEN_410 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? tag_8 : _GEN_312; // @[playground/src/noop/tlb.scala 213:117 39:26]
  wire [51:0] _GEN_411 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? tag_9 : _GEN_313; // @[playground/src/noop/tlb.scala 213:117 39:26]
  wire [51:0] _GEN_412 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? tag_10 : _GEN_314; // @[playground/src/noop/tlb.scala 213:117 39:26]
  wire [51:0] _GEN_413 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? tag_11 : _GEN_315; // @[playground/src/noop/tlb.scala 213:117 39:26]
  wire [51:0] _GEN_414 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? tag_12 : _GEN_316; // @[playground/src/noop/tlb.scala 213:117 39:26]
  wire [51:0] _GEN_415 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? tag_13 : _GEN_317; // @[playground/src/noop/tlb.scala 213:117 39:26]
  wire [51:0] _GEN_416 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? tag_14 : _GEN_318; // @[playground/src/noop/tlb.scala 213:117 39:26]
  wire [51:0] _GEN_417 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? tag_15 : _GEN_319; // @[playground/src/noop/tlb.scala 213:117 39:26]
  wire  _GEN_418 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? _GEN_130 : _GEN_320; // @[playground/src/noop/tlb.scala 213:117]
  wire  _GEN_419 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? _GEN_131 : _GEN_321; // @[playground/src/noop/tlb.scala 213:117]
  wire  _GEN_420 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? _GEN_132 : _GEN_322; // @[playground/src/noop/tlb.scala 213:117]
  wire  _GEN_421 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? _GEN_133 : _GEN_323; // @[playground/src/noop/tlb.scala 213:117]
  wire  _GEN_422 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? _GEN_134 : _GEN_324; // @[playground/src/noop/tlb.scala 213:117]
  wire  _GEN_423 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? _GEN_135 : _GEN_325; // @[playground/src/noop/tlb.scala 213:117]
  wire  _GEN_424 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? _GEN_136 : _GEN_326; // @[playground/src/noop/tlb.scala 213:117]
  wire  _GEN_425 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? _GEN_137 : _GEN_327; // @[playground/src/noop/tlb.scala 213:117]
  wire  _GEN_426 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? _GEN_138 : _GEN_328; // @[playground/src/noop/tlb.scala 213:117]
  wire  _GEN_427 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? _GEN_139 : _GEN_329; // @[playground/src/noop/tlb.scala 213:117]
  wire  _GEN_428 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? _GEN_140 : _GEN_330; // @[playground/src/noop/tlb.scala 213:117]
  wire  _GEN_429 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? _GEN_141 : _GEN_331; // @[playground/src/noop/tlb.scala 213:117]
  wire  _GEN_430 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? _GEN_142 : _GEN_332; // @[playground/src/noop/tlb.scala 213:117]
  wire  _GEN_431 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? _GEN_143 : _GEN_333; // @[playground/src/noop/tlb.scala 213:117]
  wire  _GEN_432 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? _GEN_144 : _GEN_334; // @[playground/src/noop/tlb.scala 213:117]
  wire  _GEN_433 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? _GEN_145 : _GEN_335; // @[playground/src/noop/tlb.scala 213:117]
  wire [19:0] _GEN_434 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? paddr_0 : _GEN_336; // @[playground/src/noop/tlb.scala 213:117 40:26]
  wire [19:0] _GEN_435 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? paddr_1 : _GEN_337; // @[playground/src/noop/tlb.scala 213:117 40:26]
  wire [19:0] _GEN_436 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? paddr_2 : _GEN_338; // @[playground/src/noop/tlb.scala 213:117 40:26]
  wire [19:0] _GEN_437 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? paddr_3 : _GEN_339; // @[playground/src/noop/tlb.scala 213:117 40:26]
  wire [19:0] _GEN_438 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? paddr_4 : _GEN_340; // @[playground/src/noop/tlb.scala 213:117 40:26]
  wire [19:0] _GEN_439 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? paddr_5 : _GEN_341; // @[playground/src/noop/tlb.scala 213:117 40:26]
  wire [19:0] _GEN_440 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? paddr_6 : _GEN_342; // @[playground/src/noop/tlb.scala 213:117 40:26]
  wire [19:0] _GEN_441 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? paddr_7 : _GEN_343; // @[playground/src/noop/tlb.scala 213:117 40:26]
  wire [19:0] _GEN_442 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? paddr_8 : _GEN_344; // @[playground/src/noop/tlb.scala 213:117 40:26]
  wire [19:0] _GEN_443 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? paddr_9 : _GEN_345; // @[playground/src/noop/tlb.scala 213:117 40:26]
  wire [19:0] _GEN_444 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? paddr_10 : _GEN_346; // @[playground/src/noop/tlb.scala 213:117 40:26]
  wire [19:0] _GEN_445 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? paddr_11 : _GEN_347; // @[playground/src/noop/tlb.scala 213:117 40:26]
  wire [19:0] _GEN_446 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? paddr_12 : _GEN_348; // @[playground/src/noop/tlb.scala 213:117 40:26]
  wire [19:0] _GEN_447 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? paddr_13 : _GEN_349; // @[playground/src/noop/tlb.scala 213:117 40:26]
  wire [19:0] _GEN_448 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? paddr_14 : _GEN_350; // @[playground/src/noop/tlb.scala 213:117 40:26]
  wire [19:0] _GEN_449 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? paddr_15 : _GEN_351; // @[playground/src/noop/tlb.scala 213:117 40:26]
  wire [31:0] _GEN_450 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? pte_addr_0 : _GEN_352; // @[playground/src/noop/tlb.scala 213:117 42:30]
  wire [31:0] _GEN_451 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? pte_addr_1 : _GEN_353; // @[playground/src/noop/tlb.scala 213:117 42:30]
  wire [31:0] _GEN_452 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? pte_addr_2 : _GEN_354; // @[playground/src/noop/tlb.scala 213:117 42:30]
  wire [31:0] _GEN_453 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? pte_addr_3 : _GEN_355; // @[playground/src/noop/tlb.scala 213:117 42:30]
  wire [31:0] _GEN_454 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? pte_addr_4 : _GEN_356; // @[playground/src/noop/tlb.scala 213:117 42:30]
  wire [31:0] _GEN_455 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? pte_addr_5 : _GEN_357; // @[playground/src/noop/tlb.scala 213:117 42:30]
  wire [31:0] _GEN_456 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? pte_addr_6 : _GEN_358; // @[playground/src/noop/tlb.scala 213:117 42:30]
  wire [31:0] _GEN_457 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? pte_addr_7 : _GEN_359; // @[playground/src/noop/tlb.scala 213:117 42:30]
  wire [31:0] _GEN_458 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? pte_addr_8 : _GEN_360; // @[playground/src/noop/tlb.scala 213:117 42:30]
  wire [31:0] _GEN_459 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? pte_addr_9 : _GEN_361; // @[playground/src/noop/tlb.scala 213:117 42:30]
  wire [31:0] _GEN_460 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? pte_addr_10 : _GEN_362; // @[playground/src/noop/tlb.scala 213:117 42:30]
  wire [31:0] _GEN_461 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? pte_addr_11 : _GEN_363; // @[playground/src/noop/tlb.scala 213:117 42:30]
  wire [31:0] _GEN_462 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? pte_addr_12 : _GEN_364; // @[playground/src/noop/tlb.scala 213:117 42:30]
  wire [31:0] _GEN_463 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? pte_addr_13 : _GEN_365; // @[playground/src/noop/tlb.scala 213:117 42:30]
  wire [31:0] _GEN_464 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? pte_addr_14 : _GEN_366; // @[playground/src/noop/tlb.scala 213:117 42:30]
  wire [31:0] _GEN_465 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? pte_addr_15 : _GEN_367; // @[playground/src/noop/tlb.scala 213:117 42:30]
  wire [1:0] _GEN_466 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? pte_level_0 : _GEN_368; // @[playground/src/noop/tlb.scala 213:117 43:30]
  wire [1:0] _GEN_467 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? pte_level_1 : _GEN_369; // @[playground/src/noop/tlb.scala 213:117 43:30]
  wire [1:0] _GEN_468 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? pte_level_2 : _GEN_370; // @[playground/src/noop/tlb.scala 213:117 43:30]
  wire [1:0] _GEN_469 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? pte_level_3 : _GEN_371; // @[playground/src/noop/tlb.scala 213:117 43:30]
  wire [1:0] _GEN_470 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? pte_level_4 : _GEN_372; // @[playground/src/noop/tlb.scala 213:117 43:30]
  wire [1:0] _GEN_471 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? pte_level_5 : _GEN_373; // @[playground/src/noop/tlb.scala 213:117 43:30]
  wire [1:0] _GEN_472 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? pte_level_6 : _GEN_374; // @[playground/src/noop/tlb.scala 213:117 43:30]
  wire [1:0] _GEN_473 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? pte_level_7 : _GEN_375; // @[playground/src/noop/tlb.scala 213:117 43:30]
  wire [1:0] _GEN_474 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? pte_level_8 : _GEN_376; // @[playground/src/noop/tlb.scala 213:117 43:30]
  wire [1:0] _GEN_475 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? pte_level_9 : _GEN_377; // @[playground/src/noop/tlb.scala 213:117 43:30]
  wire [1:0] _GEN_476 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? pte_level_10 : _GEN_378; // @[playground/src/noop/tlb.scala 213:117 43:30]
  wire [1:0] _GEN_477 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? pte_level_11 : _GEN_379; // @[playground/src/noop/tlb.scala 213:117 43:30]
  wire [1:0] _GEN_478 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? pte_level_12 : _GEN_380; // @[playground/src/noop/tlb.scala 213:117 43:30]
  wire [1:0] _GEN_479 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? pte_level_13 : _GEN_381; // @[playground/src/noop/tlb.scala 213:117 43:30]
  wire [1:0] _GEN_480 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? pte_level_14 : _GEN_382; // @[playground/src/noop/tlb.scala 213:117 43:30]
  wire [1:0] _GEN_481 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? pte_level_15 : _GEN_383; // @[playground/src/noop/tlb.scala 213:117 43:30]
  wire [9:0] _GEN_482 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? info_0 : _GEN_384; // @[playground/src/noop/tlb.scala 213:117 41:26]
  wire [9:0] _GEN_483 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? info_1 : _GEN_385; // @[playground/src/noop/tlb.scala 213:117 41:26]
  wire [9:0] _GEN_484 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? info_2 : _GEN_386; // @[playground/src/noop/tlb.scala 213:117 41:26]
  wire [9:0] _GEN_485 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? info_3 : _GEN_387; // @[playground/src/noop/tlb.scala 213:117 41:26]
  wire [9:0] _GEN_486 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? info_4 : _GEN_388; // @[playground/src/noop/tlb.scala 213:117 41:26]
  wire [9:0] _GEN_487 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? info_5 : _GEN_389; // @[playground/src/noop/tlb.scala 213:117 41:26]
  wire [9:0] _GEN_488 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? info_6 : _GEN_390; // @[playground/src/noop/tlb.scala 213:117 41:26]
  wire [9:0] _GEN_489 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? info_7 : _GEN_391; // @[playground/src/noop/tlb.scala 213:117 41:26]
  wire [9:0] _GEN_490 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? info_8 : _GEN_392; // @[playground/src/noop/tlb.scala 213:117 41:26]
  wire [9:0] _GEN_491 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? info_9 : _GEN_393; // @[playground/src/noop/tlb.scala 213:117 41:26]
  wire [9:0] _GEN_492 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? info_10 : _GEN_394; // @[playground/src/noop/tlb.scala 213:117 41:26]
  wire [9:0] _GEN_493 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? info_11 : _GEN_395; // @[playground/src/noop/tlb.scala 213:117 41:26]
  wire [9:0] _GEN_494 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? info_12 : _GEN_396; // @[playground/src/noop/tlb.scala 213:117 41:26]
  wire [9:0] _GEN_495 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? info_13 : _GEN_397; // @[playground/src/noop/tlb.scala 213:117 41:26]
  wire [9:0] _GEN_496 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? info_14 : _GEN_398; // @[playground/src/noop/tlb.scala 213:117 41:26]
  wire [9:0] _GEN_497 = level == 2'h1 & io_dcacheRW_rdata[18:10] != 9'h0 | level == 2'h2 & io_dcacheRW_rdata[27:10] != 18'h0
     ? info_15 : _GEN_399; // @[playground/src/noop/tlb.scala 213:117 41:26]
  wire  _GEN_499 = _T_112 | _GEN_401; // @[playground/src/noop/tlb.scala 209:99 212:40]
  wire [51:0] _GEN_500 = _T_112 ? tag_0 : _GEN_402; // @[playground/src/noop/tlb.scala 209:99 39:26]
  wire [51:0] _GEN_501 = _T_112 ? tag_1 : _GEN_403; // @[playground/src/noop/tlb.scala 209:99 39:26]
  wire [51:0] _GEN_502 = _T_112 ? tag_2 : _GEN_404; // @[playground/src/noop/tlb.scala 209:99 39:26]
  wire [51:0] _GEN_503 = _T_112 ? tag_3 : _GEN_405; // @[playground/src/noop/tlb.scala 209:99 39:26]
  wire [51:0] _GEN_504 = _T_112 ? tag_4 : _GEN_406; // @[playground/src/noop/tlb.scala 209:99 39:26]
  wire [51:0] _GEN_505 = _T_112 ? tag_5 : _GEN_407; // @[playground/src/noop/tlb.scala 209:99 39:26]
  wire [51:0] _GEN_506 = _T_112 ? tag_6 : _GEN_408; // @[playground/src/noop/tlb.scala 209:99 39:26]
  wire [51:0] _GEN_507 = _T_112 ? tag_7 : _GEN_409; // @[playground/src/noop/tlb.scala 209:99 39:26]
  wire [51:0] _GEN_508 = _T_112 ? tag_8 : _GEN_410; // @[playground/src/noop/tlb.scala 209:99 39:26]
  wire [51:0] _GEN_509 = _T_112 ? tag_9 : _GEN_411; // @[playground/src/noop/tlb.scala 209:99 39:26]
  wire [51:0] _GEN_510 = _T_112 ? tag_10 : _GEN_412; // @[playground/src/noop/tlb.scala 209:99 39:26]
  wire [51:0] _GEN_511 = _T_112 ? tag_11 : _GEN_413; // @[playground/src/noop/tlb.scala 209:99 39:26]
  wire [51:0] _GEN_512 = _T_112 ? tag_12 : _GEN_414; // @[playground/src/noop/tlb.scala 209:99 39:26]
  wire [51:0] _GEN_513 = _T_112 ? tag_13 : _GEN_415; // @[playground/src/noop/tlb.scala 209:99 39:26]
  wire [51:0] _GEN_514 = _T_112 ? tag_14 : _GEN_416; // @[playground/src/noop/tlb.scala 209:99 39:26]
  wire [51:0] _GEN_515 = _T_112 ? tag_15 : _GEN_417; // @[playground/src/noop/tlb.scala 209:99 39:26]
  wire  _GEN_516 = _T_112 ? _GEN_130 : _GEN_418; // @[playground/src/noop/tlb.scala 209:99]
  wire  _GEN_517 = _T_112 ? _GEN_131 : _GEN_419; // @[playground/src/noop/tlb.scala 209:99]
  wire  _GEN_518 = _T_112 ? _GEN_132 : _GEN_420; // @[playground/src/noop/tlb.scala 209:99]
  wire  _GEN_519 = _T_112 ? _GEN_133 : _GEN_421; // @[playground/src/noop/tlb.scala 209:99]
  wire  _GEN_520 = _T_112 ? _GEN_134 : _GEN_422; // @[playground/src/noop/tlb.scala 209:99]
  wire  _GEN_521 = _T_112 ? _GEN_135 : _GEN_423; // @[playground/src/noop/tlb.scala 209:99]
  wire  _GEN_522 = _T_112 ? _GEN_136 : _GEN_424; // @[playground/src/noop/tlb.scala 209:99]
  wire  _GEN_523 = _T_112 ? _GEN_137 : _GEN_425; // @[playground/src/noop/tlb.scala 209:99]
  wire  _GEN_524 = _T_112 ? _GEN_138 : _GEN_426; // @[playground/src/noop/tlb.scala 209:99]
  wire  _GEN_525 = _T_112 ? _GEN_139 : _GEN_427; // @[playground/src/noop/tlb.scala 209:99]
  wire  _GEN_526 = _T_112 ? _GEN_140 : _GEN_428; // @[playground/src/noop/tlb.scala 209:99]
  wire  _GEN_527 = _T_112 ? _GEN_141 : _GEN_429; // @[playground/src/noop/tlb.scala 209:99]
  wire  _GEN_528 = _T_112 ? _GEN_142 : _GEN_430; // @[playground/src/noop/tlb.scala 209:99]
  wire  _GEN_529 = _T_112 ? _GEN_143 : _GEN_431; // @[playground/src/noop/tlb.scala 209:99]
  wire  _GEN_530 = _T_112 ? _GEN_144 : _GEN_432; // @[playground/src/noop/tlb.scala 209:99]
  wire  _GEN_531 = _T_112 ? _GEN_145 : _GEN_433; // @[playground/src/noop/tlb.scala 209:99]
  wire [19:0] _GEN_532 = _T_112 ? paddr_0 : _GEN_434; // @[playground/src/noop/tlb.scala 209:99 40:26]
  wire [19:0] _GEN_533 = _T_112 ? paddr_1 : _GEN_435; // @[playground/src/noop/tlb.scala 209:99 40:26]
  wire [19:0] _GEN_534 = _T_112 ? paddr_2 : _GEN_436; // @[playground/src/noop/tlb.scala 209:99 40:26]
  wire [19:0] _GEN_535 = _T_112 ? paddr_3 : _GEN_437; // @[playground/src/noop/tlb.scala 209:99 40:26]
  wire [19:0] _GEN_536 = _T_112 ? paddr_4 : _GEN_438; // @[playground/src/noop/tlb.scala 209:99 40:26]
  wire [19:0] _GEN_537 = _T_112 ? paddr_5 : _GEN_439; // @[playground/src/noop/tlb.scala 209:99 40:26]
  wire [19:0] _GEN_538 = _T_112 ? paddr_6 : _GEN_440; // @[playground/src/noop/tlb.scala 209:99 40:26]
  wire [19:0] _GEN_539 = _T_112 ? paddr_7 : _GEN_441; // @[playground/src/noop/tlb.scala 209:99 40:26]
  wire [19:0] _GEN_540 = _T_112 ? paddr_8 : _GEN_442; // @[playground/src/noop/tlb.scala 209:99 40:26]
  wire [19:0] _GEN_541 = _T_112 ? paddr_9 : _GEN_443; // @[playground/src/noop/tlb.scala 209:99 40:26]
  wire [19:0] _GEN_542 = _T_112 ? paddr_10 : _GEN_444; // @[playground/src/noop/tlb.scala 209:99 40:26]
  wire [19:0] _GEN_543 = _T_112 ? paddr_11 : _GEN_445; // @[playground/src/noop/tlb.scala 209:99 40:26]
  wire [19:0] _GEN_544 = _T_112 ? paddr_12 : _GEN_446; // @[playground/src/noop/tlb.scala 209:99 40:26]
  wire [19:0] _GEN_545 = _T_112 ? paddr_13 : _GEN_447; // @[playground/src/noop/tlb.scala 209:99 40:26]
  wire [19:0] _GEN_546 = _T_112 ? paddr_14 : _GEN_448; // @[playground/src/noop/tlb.scala 209:99 40:26]
  wire [19:0] _GEN_547 = _T_112 ? paddr_15 : _GEN_449; // @[playground/src/noop/tlb.scala 209:99 40:26]
  wire [31:0] _GEN_548 = _T_112 ? pte_addr_0 : _GEN_450; // @[playground/src/noop/tlb.scala 209:99 42:30]
  wire [31:0] _GEN_549 = _T_112 ? pte_addr_1 : _GEN_451; // @[playground/src/noop/tlb.scala 209:99 42:30]
  wire [31:0] _GEN_550 = _T_112 ? pte_addr_2 : _GEN_452; // @[playground/src/noop/tlb.scala 209:99 42:30]
  wire [31:0] _GEN_551 = _T_112 ? pte_addr_3 : _GEN_453; // @[playground/src/noop/tlb.scala 209:99 42:30]
  wire [31:0] _GEN_552 = _T_112 ? pte_addr_4 : _GEN_454; // @[playground/src/noop/tlb.scala 209:99 42:30]
  wire [31:0] _GEN_553 = _T_112 ? pte_addr_5 : _GEN_455; // @[playground/src/noop/tlb.scala 209:99 42:30]
  wire [31:0] _GEN_554 = _T_112 ? pte_addr_6 : _GEN_456; // @[playground/src/noop/tlb.scala 209:99 42:30]
  wire [31:0] _GEN_555 = _T_112 ? pte_addr_7 : _GEN_457; // @[playground/src/noop/tlb.scala 209:99 42:30]
  wire [31:0] _GEN_556 = _T_112 ? pte_addr_8 : _GEN_458; // @[playground/src/noop/tlb.scala 209:99 42:30]
  wire [31:0] _GEN_557 = _T_112 ? pte_addr_9 : _GEN_459; // @[playground/src/noop/tlb.scala 209:99 42:30]
  wire [31:0] _GEN_558 = _T_112 ? pte_addr_10 : _GEN_460; // @[playground/src/noop/tlb.scala 209:99 42:30]
  wire [31:0] _GEN_559 = _T_112 ? pte_addr_11 : _GEN_461; // @[playground/src/noop/tlb.scala 209:99 42:30]
  wire [31:0] _GEN_560 = _T_112 ? pte_addr_12 : _GEN_462; // @[playground/src/noop/tlb.scala 209:99 42:30]
  wire [31:0] _GEN_561 = _T_112 ? pte_addr_13 : _GEN_463; // @[playground/src/noop/tlb.scala 209:99 42:30]
  wire [31:0] _GEN_562 = _T_112 ? pte_addr_14 : _GEN_464; // @[playground/src/noop/tlb.scala 209:99 42:30]
  wire [31:0] _GEN_563 = _T_112 ? pte_addr_15 : _GEN_465; // @[playground/src/noop/tlb.scala 209:99 42:30]
  wire [1:0] _GEN_564 = _T_112 ? pte_level_0 : _GEN_466; // @[playground/src/noop/tlb.scala 209:99 43:30]
  wire [1:0] _GEN_565 = _T_112 ? pte_level_1 : _GEN_467; // @[playground/src/noop/tlb.scala 209:99 43:30]
  wire [1:0] _GEN_566 = _T_112 ? pte_level_2 : _GEN_468; // @[playground/src/noop/tlb.scala 209:99 43:30]
  wire [1:0] _GEN_567 = _T_112 ? pte_level_3 : _GEN_469; // @[playground/src/noop/tlb.scala 209:99 43:30]
  wire [1:0] _GEN_568 = _T_112 ? pte_level_4 : _GEN_470; // @[playground/src/noop/tlb.scala 209:99 43:30]
  wire [1:0] _GEN_569 = _T_112 ? pte_level_5 : _GEN_471; // @[playground/src/noop/tlb.scala 209:99 43:30]
  wire [1:0] _GEN_570 = _T_112 ? pte_level_6 : _GEN_472; // @[playground/src/noop/tlb.scala 209:99 43:30]
  wire [1:0] _GEN_571 = _T_112 ? pte_level_7 : _GEN_473; // @[playground/src/noop/tlb.scala 209:99 43:30]
  wire [1:0] _GEN_572 = _T_112 ? pte_level_8 : _GEN_474; // @[playground/src/noop/tlb.scala 209:99 43:30]
  wire [1:0] _GEN_573 = _T_112 ? pte_level_9 : _GEN_475; // @[playground/src/noop/tlb.scala 209:99 43:30]
  wire [1:0] _GEN_574 = _T_112 ? pte_level_10 : _GEN_476; // @[playground/src/noop/tlb.scala 209:99 43:30]
  wire [1:0] _GEN_575 = _T_112 ? pte_level_11 : _GEN_477; // @[playground/src/noop/tlb.scala 209:99 43:30]
  wire [1:0] _GEN_576 = _T_112 ? pte_level_12 : _GEN_478; // @[playground/src/noop/tlb.scala 209:99 43:30]
  wire [1:0] _GEN_577 = _T_112 ? pte_level_13 : _GEN_479; // @[playground/src/noop/tlb.scala 209:99 43:30]
  wire [1:0] _GEN_578 = _T_112 ? pte_level_14 : _GEN_480; // @[playground/src/noop/tlb.scala 209:99 43:30]
  wire [1:0] _GEN_579 = _T_112 ? pte_level_15 : _GEN_481; // @[playground/src/noop/tlb.scala 209:99 43:30]
  wire [9:0] _GEN_580 = _T_112 ? info_0 : _GEN_482; // @[playground/src/noop/tlb.scala 209:99 41:26]
  wire [9:0] _GEN_581 = _T_112 ? info_1 : _GEN_483; // @[playground/src/noop/tlb.scala 209:99 41:26]
  wire [9:0] _GEN_582 = _T_112 ? info_2 : _GEN_484; // @[playground/src/noop/tlb.scala 209:99 41:26]
  wire [9:0] _GEN_583 = _T_112 ? info_3 : _GEN_485; // @[playground/src/noop/tlb.scala 209:99 41:26]
  wire [9:0] _GEN_584 = _T_112 ? info_4 : _GEN_486; // @[playground/src/noop/tlb.scala 209:99 41:26]
  wire [9:0] _GEN_585 = _T_112 ? info_5 : _GEN_487; // @[playground/src/noop/tlb.scala 209:99 41:26]
  wire [9:0] _GEN_586 = _T_112 ? info_6 : _GEN_488; // @[playground/src/noop/tlb.scala 209:99 41:26]
  wire [9:0] _GEN_587 = _T_112 ? info_7 : _GEN_489; // @[playground/src/noop/tlb.scala 209:99 41:26]
  wire [9:0] _GEN_588 = _T_112 ? info_8 : _GEN_490; // @[playground/src/noop/tlb.scala 209:99 41:26]
  wire [9:0] _GEN_589 = _T_112 ? info_9 : _GEN_491; // @[playground/src/noop/tlb.scala 209:99 41:26]
  wire [9:0] _GEN_590 = _T_112 ? info_10 : _GEN_492; // @[playground/src/noop/tlb.scala 209:99 41:26]
  wire [9:0] _GEN_591 = _T_112 ? info_11 : _GEN_493; // @[playground/src/noop/tlb.scala 209:99 41:26]
  wire [9:0] _GEN_592 = _T_112 ? info_12 : _GEN_494; // @[playground/src/noop/tlb.scala 209:99 41:26]
  wire [9:0] _GEN_593 = _T_112 ? info_13 : _GEN_495; // @[playground/src/noop/tlb.scala 209:99 41:26]
  wire [9:0] _GEN_594 = _T_112 ? info_14 : _GEN_496; // @[playground/src/noop/tlb.scala 209:99 41:26]
  wire [9:0] _GEN_595 = _T_112 ? info_15 : _GEN_497; // @[playground/src/noop/tlb.scala 209:99 41:26]
  wire  _GEN_597 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] | _GEN_499; // @[playground/src/noop/tlb.scala 203:87 206:40]
  wire [51:0] _GEN_598 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? tag_0 : _GEN_500; // @[playground/src/noop/tlb.scala 203:87 39:26]
  wire [51:0] _GEN_599 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? tag_1 : _GEN_501; // @[playground/src/noop/tlb.scala 203:87 39:26]
  wire [51:0] _GEN_600 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? tag_2 : _GEN_502; // @[playground/src/noop/tlb.scala 203:87 39:26]
  wire [51:0] _GEN_601 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? tag_3 : _GEN_503; // @[playground/src/noop/tlb.scala 203:87 39:26]
  wire [51:0] _GEN_602 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? tag_4 : _GEN_504; // @[playground/src/noop/tlb.scala 203:87 39:26]
  wire [51:0] _GEN_603 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? tag_5 : _GEN_505; // @[playground/src/noop/tlb.scala 203:87 39:26]
  wire [51:0] _GEN_604 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? tag_6 : _GEN_506; // @[playground/src/noop/tlb.scala 203:87 39:26]
  wire [51:0] _GEN_605 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? tag_7 : _GEN_507; // @[playground/src/noop/tlb.scala 203:87 39:26]
  wire [51:0] _GEN_606 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? tag_8 : _GEN_508; // @[playground/src/noop/tlb.scala 203:87 39:26]
  wire [51:0] _GEN_607 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? tag_9 : _GEN_509; // @[playground/src/noop/tlb.scala 203:87 39:26]
  wire [51:0] _GEN_608 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? tag_10 : _GEN_510; // @[playground/src/noop/tlb.scala 203:87 39:26]
  wire [51:0] _GEN_609 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? tag_11 : _GEN_511; // @[playground/src/noop/tlb.scala 203:87 39:26]
  wire [51:0] _GEN_610 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? tag_12 : _GEN_512; // @[playground/src/noop/tlb.scala 203:87 39:26]
  wire [51:0] _GEN_611 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? tag_13 : _GEN_513; // @[playground/src/noop/tlb.scala 203:87 39:26]
  wire [51:0] _GEN_612 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? tag_14 : _GEN_514; // @[playground/src/noop/tlb.scala 203:87 39:26]
  wire [51:0] _GEN_613 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? tag_15 : _GEN_515; // @[playground/src/noop/tlb.scala 203:87 39:26]
  wire  _GEN_614 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? _GEN_130 : _GEN_516; // @[playground/src/noop/tlb.scala 203:87]
  wire  _GEN_615 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? _GEN_131 : _GEN_517; // @[playground/src/noop/tlb.scala 203:87]
  wire  _GEN_616 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? _GEN_132 : _GEN_518; // @[playground/src/noop/tlb.scala 203:87]
  wire  _GEN_617 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? _GEN_133 : _GEN_519; // @[playground/src/noop/tlb.scala 203:87]
  wire  _GEN_618 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? _GEN_134 : _GEN_520; // @[playground/src/noop/tlb.scala 203:87]
  wire  _GEN_619 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? _GEN_135 : _GEN_521; // @[playground/src/noop/tlb.scala 203:87]
  wire  _GEN_620 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? _GEN_136 : _GEN_522; // @[playground/src/noop/tlb.scala 203:87]
  wire  _GEN_621 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? _GEN_137 : _GEN_523; // @[playground/src/noop/tlb.scala 203:87]
  wire  _GEN_622 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? _GEN_138 : _GEN_524; // @[playground/src/noop/tlb.scala 203:87]
  wire  _GEN_623 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? _GEN_139 : _GEN_525; // @[playground/src/noop/tlb.scala 203:87]
  wire  _GEN_624 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? _GEN_140 : _GEN_526; // @[playground/src/noop/tlb.scala 203:87]
  wire  _GEN_625 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? _GEN_141 : _GEN_527; // @[playground/src/noop/tlb.scala 203:87]
  wire  _GEN_626 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? _GEN_142 : _GEN_528; // @[playground/src/noop/tlb.scala 203:87]
  wire  _GEN_627 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? _GEN_143 : _GEN_529; // @[playground/src/noop/tlb.scala 203:87]
  wire  _GEN_628 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? _GEN_144 : _GEN_530; // @[playground/src/noop/tlb.scala 203:87]
  wire  _GEN_629 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? _GEN_145 : _GEN_531; // @[playground/src/noop/tlb.scala 203:87]
  wire [19:0] _GEN_630 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? paddr_0 : _GEN_532; // @[playground/src/noop/tlb.scala 203:87 40:26]
  wire [19:0] _GEN_631 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? paddr_1 : _GEN_533; // @[playground/src/noop/tlb.scala 203:87 40:26]
  wire [19:0] _GEN_632 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? paddr_2 : _GEN_534; // @[playground/src/noop/tlb.scala 203:87 40:26]
  wire [19:0] _GEN_633 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? paddr_3 : _GEN_535; // @[playground/src/noop/tlb.scala 203:87 40:26]
  wire [19:0] _GEN_634 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? paddr_4 : _GEN_536; // @[playground/src/noop/tlb.scala 203:87 40:26]
  wire [19:0] _GEN_635 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? paddr_5 : _GEN_537; // @[playground/src/noop/tlb.scala 203:87 40:26]
  wire [19:0] _GEN_636 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? paddr_6 : _GEN_538; // @[playground/src/noop/tlb.scala 203:87 40:26]
  wire [19:0] _GEN_637 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? paddr_7 : _GEN_539; // @[playground/src/noop/tlb.scala 203:87 40:26]
  wire [19:0] _GEN_638 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? paddr_8 : _GEN_540; // @[playground/src/noop/tlb.scala 203:87 40:26]
  wire [19:0] _GEN_639 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? paddr_9 : _GEN_541; // @[playground/src/noop/tlb.scala 203:87 40:26]
  wire [19:0] _GEN_640 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? paddr_10 : _GEN_542; // @[playground/src/noop/tlb.scala 203:87 40:26]
  wire [19:0] _GEN_641 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? paddr_11 : _GEN_543; // @[playground/src/noop/tlb.scala 203:87 40:26]
  wire [19:0] _GEN_642 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? paddr_12 : _GEN_544; // @[playground/src/noop/tlb.scala 203:87 40:26]
  wire [19:0] _GEN_643 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? paddr_13 : _GEN_545; // @[playground/src/noop/tlb.scala 203:87 40:26]
  wire [19:0] _GEN_644 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? paddr_14 : _GEN_546; // @[playground/src/noop/tlb.scala 203:87 40:26]
  wire [19:0] _GEN_645 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? paddr_15 : _GEN_547; // @[playground/src/noop/tlb.scala 203:87 40:26]
  wire [31:0] _GEN_646 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? pte_addr_0 : _GEN_548; // @[playground/src/noop/tlb.scala 203:87 42:30]
  wire [31:0] _GEN_647 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? pte_addr_1 : _GEN_549; // @[playground/src/noop/tlb.scala 203:87 42:30]
  wire [31:0] _GEN_648 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? pte_addr_2 : _GEN_550; // @[playground/src/noop/tlb.scala 203:87 42:30]
  wire [31:0] _GEN_649 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? pte_addr_3 : _GEN_551; // @[playground/src/noop/tlb.scala 203:87 42:30]
  wire [31:0] _GEN_650 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? pte_addr_4 : _GEN_552; // @[playground/src/noop/tlb.scala 203:87 42:30]
  wire [31:0] _GEN_651 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? pte_addr_5 : _GEN_553; // @[playground/src/noop/tlb.scala 203:87 42:30]
  wire [31:0] _GEN_652 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? pte_addr_6 : _GEN_554; // @[playground/src/noop/tlb.scala 203:87 42:30]
  wire [31:0] _GEN_653 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? pte_addr_7 : _GEN_555; // @[playground/src/noop/tlb.scala 203:87 42:30]
  wire [31:0] _GEN_654 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? pte_addr_8 : _GEN_556; // @[playground/src/noop/tlb.scala 203:87 42:30]
  wire [31:0] _GEN_655 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? pte_addr_9 : _GEN_557; // @[playground/src/noop/tlb.scala 203:87 42:30]
  wire [31:0] _GEN_656 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? pte_addr_10 : _GEN_558; // @[playground/src/noop/tlb.scala 203:87 42:30]
  wire [31:0] _GEN_657 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? pte_addr_11 : _GEN_559; // @[playground/src/noop/tlb.scala 203:87 42:30]
  wire [31:0] _GEN_658 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? pte_addr_12 : _GEN_560; // @[playground/src/noop/tlb.scala 203:87 42:30]
  wire [31:0] _GEN_659 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? pte_addr_13 : _GEN_561; // @[playground/src/noop/tlb.scala 203:87 42:30]
  wire [31:0] _GEN_660 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? pte_addr_14 : _GEN_562; // @[playground/src/noop/tlb.scala 203:87 42:30]
  wire [31:0] _GEN_661 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? pte_addr_15 : _GEN_563; // @[playground/src/noop/tlb.scala 203:87 42:30]
  wire [1:0] _GEN_662 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? pte_level_0 : _GEN_564; // @[playground/src/noop/tlb.scala 203:87 43:30]
  wire [1:0] _GEN_663 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? pte_level_1 : _GEN_565; // @[playground/src/noop/tlb.scala 203:87 43:30]
  wire [1:0] _GEN_664 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? pte_level_2 : _GEN_566; // @[playground/src/noop/tlb.scala 203:87 43:30]
  wire [1:0] _GEN_665 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? pte_level_3 : _GEN_567; // @[playground/src/noop/tlb.scala 203:87 43:30]
  wire [1:0] _GEN_666 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? pte_level_4 : _GEN_568; // @[playground/src/noop/tlb.scala 203:87 43:30]
  wire [1:0] _GEN_667 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? pte_level_5 : _GEN_569; // @[playground/src/noop/tlb.scala 203:87 43:30]
  wire [1:0] _GEN_668 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? pte_level_6 : _GEN_570; // @[playground/src/noop/tlb.scala 203:87 43:30]
  wire [1:0] _GEN_669 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? pte_level_7 : _GEN_571; // @[playground/src/noop/tlb.scala 203:87 43:30]
  wire [1:0] _GEN_670 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? pte_level_8 : _GEN_572; // @[playground/src/noop/tlb.scala 203:87 43:30]
  wire [1:0] _GEN_671 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? pte_level_9 : _GEN_573; // @[playground/src/noop/tlb.scala 203:87 43:30]
  wire [1:0] _GEN_672 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? pte_level_10 : _GEN_574; // @[playground/src/noop/tlb.scala 203:87 43:30]
  wire [1:0] _GEN_673 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? pte_level_11 : _GEN_575; // @[playground/src/noop/tlb.scala 203:87 43:30]
  wire [1:0] _GEN_674 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? pte_level_12 : _GEN_576; // @[playground/src/noop/tlb.scala 203:87 43:30]
  wire [1:0] _GEN_675 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? pte_level_13 : _GEN_577; // @[playground/src/noop/tlb.scala 203:87 43:30]
  wire [1:0] _GEN_676 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? pte_level_14 : _GEN_578; // @[playground/src/noop/tlb.scala 203:87 43:30]
  wire [1:0] _GEN_677 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? pte_level_15 : _GEN_579; // @[playground/src/noop/tlb.scala 203:87 43:30]
  wire [9:0] _GEN_678 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? info_0 : _GEN_580; // @[playground/src/noop/tlb.scala 203:87 41:26]
  wire [9:0] _GEN_679 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? info_1 : _GEN_581; // @[playground/src/noop/tlb.scala 203:87 41:26]
  wire [9:0] _GEN_680 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? info_2 : _GEN_582; // @[playground/src/noop/tlb.scala 203:87 41:26]
  wire [9:0] _GEN_681 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? info_3 : _GEN_583; // @[playground/src/noop/tlb.scala 203:87 41:26]
  wire [9:0] _GEN_682 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? info_4 : _GEN_584; // @[playground/src/noop/tlb.scala 203:87 41:26]
  wire [9:0] _GEN_683 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? info_5 : _GEN_585; // @[playground/src/noop/tlb.scala 203:87 41:26]
  wire [9:0] _GEN_684 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? info_6 : _GEN_586; // @[playground/src/noop/tlb.scala 203:87 41:26]
  wire [9:0] _GEN_685 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? info_7 : _GEN_587; // @[playground/src/noop/tlb.scala 203:87 41:26]
  wire [9:0] _GEN_686 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? info_8 : _GEN_588; // @[playground/src/noop/tlb.scala 203:87 41:26]
  wire [9:0] _GEN_687 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? info_9 : _GEN_589; // @[playground/src/noop/tlb.scala 203:87 41:26]
  wire [9:0] _GEN_688 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? info_10 : _GEN_590; // @[playground/src/noop/tlb.scala 203:87 41:26]
  wire [9:0] _GEN_689 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? info_11 : _GEN_591; // @[playground/src/noop/tlb.scala 203:87 41:26]
  wire [9:0] _GEN_690 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? info_12 : _GEN_592; // @[playground/src/noop/tlb.scala 203:87 41:26]
  wire [9:0] _GEN_691 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? info_13 : _GEN_593; // @[playground/src/noop/tlb.scala 203:87 41:26]
  wire [9:0] _GEN_692 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? info_14 : _GEN_594; // @[playground/src/noop/tlb.scala 203:87 41:26]
  wire [9:0] _GEN_693 = ~io_dcacheRW_rdata[0] | ~io_dcacheRW_rdata[1] & io_dcacheRW_rdata[2] ? info_15 : _GEN_595; // @[playground/src/noop/tlb.scala 203:87 41:26]
  wire  _GEN_695 = _T_87 | _GEN_597; // @[playground/src/noop/tlb.scala 199:193 202:40]
  wire [51:0] _GEN_696 = _T_87 ? tag_0 : _GEN_598; // @[playground/src/noop/tlb.scala 199:193 39:26]
  wire [51:0] _GEN_697 = _T_87 ? tag_1 : _GEN_599; // @[playground/src/noop/tlb.scala 199:193 39:26]
  wire [51:0] _GEN_698 = _T_87 ? tag_2 : _GEN_600; // @[playground/src/noop/tlb.scala 199:193 39:26]
  wire [51:0] _GEN_699 = _T_87 ? tag_3 : _GEN_601; // @[playground/src/noop/tlb.scala 199:193 39:26]
  wire [51:0] _GEN_700 = _T_87 ? tag_4 : _GEN_602; // @[playground/src/noop/tlb.scala 199:193 39:26]
  wire [51:0] _GEN_701 = _T_87 ? tag_5 : _GEN_603; // @[playground/src/noop/tlb.scala 199:193 39:26]
  wire [51:0] _GEN_702 = _T_87 ? tag_6 : _GEN_604; // @[playground/src/noop/tlb.scala 199:193 39:26]
  wire [51:0] _GEN_703 = _T_87 ? tag_7 : _GEN_605; // @[playground/src/noop/tlb.scala 199:193 39:26]
  wire [51:0] _GEN_704 = _T_87 ? tag_8 : _GEN_606; // @[playground/src/noop/tlb.scala 199:193 39:26]
  wire [51:0] _GEN_705 = _T_87 ? tag_9 : _GEN_607; // @[playground/src/noop/tlb.scala 199:193 39:26]
  wire [51:0] _GEN_706 = _T_87 ? tag_10 : _GEN_608; // @[playground/src/noop/tlb.scala 199:193 39:26]
  wire [51:0] _GEN_707 = _T_87 ? tag_11 : _GEN_609; // @[playground/src/noop/tlb.scala 199:193 39:26]
  wire [51:0] _GEN_708 = _T_87 ? tag_12 : _GEN_610; // @[playground/src/noop/tlb.scala 199:193 39:26]
  wire [51:0] _GEN_709 = _T_87 ? tag_13 : _GEN_611; // @[playground/src/noop/tlb.scala 199:193 39:26]
  wire [51:0] _GEN_710 = _T_87 ? tag_14 : _GEN_612; // @[playground/src/noop/tlb.scala 199:193 39:26]
  wire [51:0] _GEN_711 = _T_87 ? tag_15 : _GEN_613; // @[playground/src/noop/tlb.scala 199:193 39:26]
  wire  _GEN_712 = _T_87 ? _GEN_130 : _GEN_614; // @[playground/src/noop/tlb.scala 199:193]
  wire  _GEN_713 = _T_87 ? _GEN_131 : _GEN_615; // @[playground/src/noop/tlb.scala 199:193]
  wire  _GEN_714 = _T_87 ? _GEN_132 : _GEN_616; // @[playground/src/noop/tlb.scala 199:193]
  wire  _GEN_715 = _T_87 ? _GEN_133 : _GEN_617; // @[playground/src/noop/tlb.scala 199:193]
  wire  _GEN_716 = _T_87 ? _GEN_134 : _GEN_618; // @[playground/src/noop/tlb.scala 199:193]
  wire  _GEN_717 = _T_87 ? _GEN_135 : _GEN_619; // @[playground/src/noop/tlb.scala 199:193]
  wire  _GEN_718 = _T_87 ? _GEN_136 : _GEN_620; // @[playground/src/noop/tlb.scala 199:193]
  wire  _GEN_719 = _T_87 ? _GEN_137 : _GEN_621; // @[playground/src/noop/tlb.scala 199:193]
  wire  _GEN_720 = _T_87 ? _GEN_138 : _GEN_622; // @[playground/src/noop/tlb.scala 199:193]
  wire  _GEN_721 = _T_87 ? _GEN_139 : _GEN_623; // @[playground/src/noop/tlb.scala 199:193]
  wire  _GEN_722 = _T_87 ? _GEN_140 : _GEN_624; // @[playground/src/noop/tlb.scala 199:193]
  wire  _GEN_723 = _T_87 ? _GEN_141 : _GEN_625; // @[playground/src/noop/tlb.scala 199:193]
  wire  _GEN_724 = _T_87 ? _GEN_142 : _GEN_626; // @[playground/src/noop/tlb.scala 199:193]
  wire  _GEN_725 = _T_87 ? _GEN_143 : _GEN_627; // @[playground/src/noop/tlb.scala 199:193]
  wire  _GEN_726 = _T_87 ? _GEN_144 : _GEN_628; // @[playground/src/noop/tlb.scala 199:193]
  wire  _GEN_727 = _T_87 ? _GEN_145 : _GEN_629; // @[playground/src/noop/tlb.scala 199:193]
  wire [19:0] _GEN_728 = _T_87 ? paddr_0 : _GEN_630; // @[playground/src/noop/tlb.scala 199:193 40:26]
  wire [19:0] _GEN_729 = _T_87 ? paddr_1 : _GEN_631; // @[playground/src/noop/tlb.scala 199:193 40:26]
  wire [19:0] _GEN_730 = _T_87 ? paddr_2 : _GEN_632; // @[playground/src/noop/tlb.scala 199:193 40:26]
  wire [19:0] _GEN_731 = _T_87 ? paddr_3 : _GEN_633; // @[playground/src/noop/tlb.scala 199:193 40:26]
  wire [19:0] _GEN_732 = _T_87 ? paddr_4 : _GEN_634; // @[playground/src/noop/tlb.scala 199:193 40:26]
  wire [19:0] _GEN_733 = _T_87 ? paddr_5 : _GEN_635; // @[playground/src/noop/tlb.scala 199:193 40:26]
  wire [19:0] _GEN_734 = _T_87 ? paddr_6 : _GEN_636; // @[playground/src/noop/tlb.scala 199:193 40:26]
  wire [19:0] _GEN_735 = _T_87 ? paddr_7 : _GEN_637; // @[playground/src/noop/tlb.scala 199:193 40:26]
  wire [19:0] _GEN_736 = _T_87 ? paddr_8 : _GEN_638; // @[playground/src/noop/tlb.scala 199:193 40:26]
  wire [19:0] _GEN_737 = _T_87 ? paddr_9 : _GEN_639; // @[playground/src/noop/tlb.scala 199:193 40:26]
  wire [19:0] _GEN_738 = _T_87 ? paddr_10 : _GEN_640; // @[playground/src/noop/tlb.scala 199:193 40:26]
  wire [19:0] _GEN_739 = _T_87 ? paddr_11 : _GEN_641; // @[playground/src/noop/tlb.scala 199:193 40:26]
  wire [19:0] _GEN_740 = _T_87 ? paddr_12 : _GEN_642; // @[playground/src/noop/tlb.scala 199:193 40:26]
  wire [19:0] _GEN_741 = _T_87 ? paddr_13 : _GEN_643; // @[playground/src/noop/tlb.scala 199:193 40:26]
  wire [19:0] _GEN_742 = _T_87 ? paddr_14 : _GEN_644; // @[playground/src/noop/tlb.scala 199:193 40:26]
  wire [19:0] _GEN_743 = _T_87 ? paddr_15 : _GEN_645; // @[playground/src/noop/tlb.scala 199:193 40:26]
  wire [31:0] _GEN_744 = _T_87 ? pte_addr_0 : _GEN_646; // @[playground/src/noop/tlb.scala 199:193 42:30]
  wire [31:0] _GEN_745 = _T_87 ? pte_addr_1 : _GEN_647; // @[playground/src/noop/tlb.scala 199:193 42:30]
  wire [31:0] _GEN_746 = _T_87 ? pte_addr_2 : _GEN_648; // @[playground/src/noop/tlb.scala 199:193 42:30]
  wire [31:0] _GEN_747 = _T_87 ? pte_addr_3 : _GEN_649; // @[playground/src/noop/tlb.scala 199:193 42:30]
  wire [31:0] _GEN_748 = _T_87 ? pte_addr_4 : _GEN_650; // @[playground/src/noop/tlb.scala 199:193 42:30]
  wire [31:0] _GEN_749 = _T_87 ? pte_addr_5 : _GEN_651; // @[playground/src/noop/tlb.scala 199:193 42:30]
  wire [31:0] _GEN_750 = _T_87 ? pte_addr_6 : _GEN_652; // @[playground/src/noop/tlb.scala 199:193 42:30]
  wire [31:0] _GEN_751 = _T_87 ? pte_addr_7 : _GEN_653; // @[playground/src/noop/tlb.scala 199:193 42:30]
  wire [31:0] _GEN_752 = _T_87 ? pte_addr_8 : _GEN_654; // @[playground/src/noop/tlb.scala 199:193 42:30]
  wire [31:0] _GEN_753 = _T_87 ? pte_addr_9 : _GEN_655; // @[playground/src/noop/tlb.scala 199:193 42:30]
  wire [31:0] _GEN_754 = _T_87 ? pte_addr_10 : _GEN_656; // @[playground/src/noop/tlb.scala 199:193 42:30]
  wire [31:0] _GEN_755 = _T_87 ? pte_addr_11 : _GEN_657; // @[playground/src/noop/tlb.scala 199:193 42:30]
  wire [31:0] _GEN_756 = _T_87 ? pte_addr_12 : _GEN_658; // @[playground/src/noop/tlb.scala 199:193 42:30]
  wire [31:0] _GEN_757 = _T_87 ? pte_addr_13 : _GEN_659; // @[playground/src/noop/tlb.scala 199:193 42:30]
  wire [31:0] _GEN_758 = _T_87 ? pte_addr_14 : _GEN_660; // @[playground/src/noop/tlb.scala 199:193 42:30]
  wire [31:0] _GEN_759 = _T_87 ? pte_addr_15 : _GEN_661; // @[playground/src/noop/tlb.scala 199:193 42:30]
  wire [1:0] _GEN_760 = _T_87 ? pte_level_0 : _GEN_662; // @[playground/src/noop/tlb.scala 199:193 43:30]
  wire [1:0] _GEN_761 = _T_87 ? pte_level_1 : _GEN_663; // @[playground/src/noop/tlb.scala 199:193 43:30]
  wire [1:0] _GEN_762 = _T_87 ? pte_level_2 : _GEN_664; // @[playground/src/noop/tlb.scala 199:193 43:30]
  wire [1:0] _GEN_763 = _T_87 ? pte_level_3 : _GEN_665; // @[playground/src/noop/tlb.scala 199:193 43:30]
  wire [1:0] _GEN_764 = _T_87 ? pte_level_4 : _GEN_666; // @[playground/src/noop/tlb.scala 199:193 43:30]
  wire [1:0] _GEN_765 = _T_87 ? pte_level_5 : _GEN_667; // @[playground/src/noop/tlb.scala 199:193 43:30]
  wire [1:0] _GEN_766 = _T_87 ? pte_level_6 : _GEN_668; // @[playground/src/noop/tlb.scala 199:193 43:30]
  wire [1:0] _GEN_767 = _T_87 ? pte_level_7 : _GEN_669; // @[playground/src/noop/tlb.scala 199:193 43:30]
  wire [1:0] _GEN_768 = _T_87 ? pte_level_8 : _GEN_670; // @[playground/src/noop/tlb.scala 199:193 43:30]
  wire [1:0] _GEN_769 = _T_87 ? pte_level_9 : _GEN_671; // @[playground/src/noop/tlb.scala 199:193 43:30]
  wire [1:0] _GEN_770 = _T_87 ? pte_level_10 : _GEN_672; // @[playground/src/noop/tlb.scala 199:193 43:30]
  wire [1:0] _GEN_771 = _T_87 ? pte_level_11 : _GEN_673; // @[playground/src/noop/tlb.scala 199:193 43:30]
  wire [1:0] _GEN_772 = _T_87 ? pte_level_12 : _GEN_674; // @[playground/src/noop/tlb.scala 199:193 43:30]
  wire [1:0] _GEN_773 = _T_87 ? pte_level_13 : _GEN_675; // @[playground/src/noop/tlb.scala 199:193 43:30]
  wire [1:0] _GEN_774 = _T_87 ? pte_level_14 : _GEN_676; // @[playground/src/noop/tlb.scala 199:193 43:30]
  wire [1:0] _GEN_775 = _T_87 ? pte_level_15 : _GEN_677; // @[playground/src/noop/tlb.scala 199:193 43:30]
  wire [9:0] _GEN_776 = _T_87 ? info_0 : _GEN_678; // @[playground/src/noop/tlb.scala 199:193 41:26]
  wire [9:0] _GEN_777 = _T_87 ? info_1 : _GEN_679; // @[playground/src/noop/tlb.scala 199:193 41:26]
  wire [9:0] _GEN_778 = _T_87 ? info_2 : _GEN_680; // @[playground/src/noop/tlb.scala 199:193 41:26]
  wire [9:0] _GEN_779 = _T_87 ? info_3 : _GEN_681; // @[playground/src/noop/tlb.scala 199:193 41:26]
  wire [9:0] _GEN_780 = _T_87 ? info_4 : _GEN_682; // @[playground/src/noop/tlb.scala 199:193 41:26]
  wire [9:0] _GEN_781 = _T_87 ? info_5 : _GEN_683; // @[playground/src/noop/tlb.scala 199:193 41:26]
  wire [9:0] _GEN_782 = _T_87 ? info_6 : _GEN_684; // @[playground/src/noop/tlb.scala 199:193 41:26]
  wire [9:0] _GEN_783 = _T_87 ? info_7 : _GEN_685; // @[playground/src/noop/tlb.scala 199:193 41:26]
  wire [9:0] _GEN_784 = _T_87 ? info_8 : _GEN_686; // @[playground/src/noop/tlb.scala 199:193 41:26]
  wire [9:0] _GEN_785 = _T_87 ? info_9 : _GEN_687; // @[playground/src/noop/tlb.scala 199:193 41:26]
  wire [9:0] _GEN_786 = _T_87 ? info_10 : _GEN_688; // @[playground/src/noop/tlb.scala 199:193 41:26]
  wire [9:0] _GEN_787 = _T_87 ? info_11 : _GEN_689; // @[playground/src/noop/tlb.scala 199:193 41:26]
  wire [9:0] _GEN_788 = _T_87 ? info_12 : _GEN_690; // @[playground/src/noop/tlb.scala 199:193 41:26]
  wire [9:0] _GEN_789 = _T_87 ? info_13 : _GEN_691; // @[playground/src/noop/tlb.scala 199:193 41:26]
  wire [9:0] _GEN_790 = _T_87 ? info_14 : _GEN_692; // @[playground/src/noop/tlb.scala 199:193 41:26]
  wire [9:0] _GEN_791 = _T_87 ? info_15 : _GEN_693; // @[playground/src/noop/tlb.scala 199:193 41:26]
  wire [1:0] _GEN_792 = _T_73 == 64'h1 ? _GEN_300 : 2'h0; // @[playground/src/noop/tlb.scala 191:76]
  wire  _GEN_793 = _T_73 == 64'h1 ? _GEN_301 : _GEN_695; // @[playground/src/noop/tlb.scala 191:76]
  wire [55:0] _GEN_794 = _T_73 == 64'h1 ? _GEN_302 : {{24'd0}, pte_addr_r}; // @[playground/src/noop/tlb.scala 191:76 47:30]
  wire [4:0] _GEN_795 = _T_73 == 64'h1 ? _GEN_303 : _GEN_297; // @[playground/src/noop/tlb.scala 191:76]
  wire [51:0] _GEN_796 = _T_73 == 64'h1 ? tag_0 : _GEN_696; // @[playground/src/noop/tlb.scala 191:76 39:26]
  wire [51:0] _GEN_797 = _T_73 == 64'h1 ? tag_1 : _GEN_697; // @[playground/src/noop/tlb.scala 191:76 39:26]
  wire [51:0] _GEN_798 = _T_73 == 64'h1 ? tag_2 : _GEN_698; // @[playground/src/noop/tlb.scala 191:76 39:26]
  wire [51:0] _GEN_799 = _T_73 == 64'h1 ? tag_3 : _GEN_699; // @[playground/src/noop/tlb.scala 191:76 39:26]
  wire [51:0] _GEN_800 = _T_73 == 64'h1 ? tag_4 : _GEN_700; // @[playground/src/noop/tlb.scala 191:76 39:26]
  wire [51:0] _GEN_801 = _T_73 == 64'h1 ? tag_5 : _GEN_701; // @[playground/src/noop/tlb.scala 191:76 39:26]
  wire [51:0] _GEN_802 = _T_73 == 64'h1 ? tag_6 : _GEN_702; // @[playground/src/noop/tlb.scala 191:76 39:26]
  wire [51:0] _GEN_803 = _T_73 == 64'h1 ? tag_7 : _GEN_703; // @[playground/src/noop/tlb.scala 191:76 39:26]
  wire [51:0] _GEN_804 = _T_73 == 64'h1 ? tag_8 : _GEN_704; // @[playground/src/noop/tlb.scala 191:76 39:26]
  wire [51:0] _GEN_805 = _T_73 == 64'h1 ? tag_9 : _GEN_705; // @[playground/src/noop/tlb.scala 191:76 39:26]
  wire [51:0] _GEN_806 = _T_73 == 64'h1 ? tag_10 : _GEN_706; // @[playground/src/noop/tlb.scala 191:76 39:26]
  wire [51:0] _GEN_807 = _T_73 == 64'h1 ? tag_11 : _GEN_707; // @[playground/src/noop/tlb.scala 191:76 39:26]
  wire [51:0] _GEN_808 = _T_73 == 64'h1 ? tag_12 : _GEN_708; // @[playground/src/noop/tlb.scala 191:76 39:26]
  wire [51:0] _GEN_809 = _T_73 == 64'h1 ? tag_13 : _GEN_709; // @[playground/src/noop/tlb.scala 191:76 39:26]
  wire [51:0] _GEN_810 = _T_73 == 64'h1 ? tag_14 : _GEN_710; // @[playground/src/noop/tlb.scala 191:76 39:26]
  wire [51:0] _GEN_811 = _T_73 == 64'h1 ? tag_15 : _GEN_711; // @[playground/src/noop/tlb.scala 191:76 39:26]
  wire  _GEN_812 = _T_73 == 64'h1 ? _GEN_130 : _GEN_712; // @[playground/src/noop/tlb.scala 191:76]
  wire  _GEN_813 = _T_73 == 64'h1 ? _GEN_131 : _GEN_713; // @[playground/src/noop/tlb.scala 191:76]
  wire  _GEN_814 = _T_73 == 64'h1 ? _GEN_132 : _GEN_714; // @[playground/src/noop/tlb.scala 191:76]
  wire  _GEN_815 = _T_73 == 64'h1 ? _GEN_133 : _GEN_715; // @[playground/src/noop/tlb.scala 191:76]
  wire  _GEN_816 = _T_73 == 64'h1 ? _GEN_134 : _GEN_716; // @[playground/src/noop/tlb.scala 191:76]
  wire  _GEN_817 = _T_73 == 64'h1 ? _GEN_135 : _GEN_717; // @[playground/src/noop/tlb.scala 191:76]
  wire  _GEN_818 = _T_73 == 64'h1 ? _GEN_136 : _GEN_718; // @[playground/src/noop/tlb.scala 191:76]
  wire  _GEN_819 = _T_73 == 64'h1 ? _GEN_137 : _GEN_719; // @[playground/src/noop/tlb.scala 191:76]
  wire  _GEN_820 = _T_73 == 64'h1 ? _GEN_138 : _GEN_720; // @[playground/src/noop/tlb.scala 191:76]
  wire  _GEN_821 = _T_73 == 64'h1 ? _GEN_139 : _GEN_721; // @[playground/src/noop/tlb.scala 191:76]
  wire  _GEN_822 = _T_73 == 64'h1 ? _GEN_140 : _GEN_722; // @[playground/src/noop/tlb.scala 191:76]
  wire  _GEN_823 = _T_73 == 64'h1 ? _GEN_141 : _GEN_723; // @[playground/src/noop/tlb.scala 191:76]
  wire  _GEN_824 = _T_73 == 64'h1 ? _GEN_142 : _GEN_724; // @[playground/src/noop/tlb.scala 191:76]
  wire  _GEN_825 = _T_73 == 64'h1 ? _GEN_143 : _GEN_725; // @[playground/src/noop/tlb.scala 191:76]
  wire  _GEN_826 = _T_73 == 64'h1 ? _GEN_144 : _GEN_726; // @[playground/src/noop/tlb.scala 191:76]
  wire  _GEN_827 = _T_73 == 64'h1 ? _GEN_145 : _GEN_727; // @[playground/src/noop/tlb.scala 191:76]
  wire [19:0] _GEN_828 = _T_73 == 64'h1 ? paddr_0 : _GEN_728; // @[playground/src/noop/tlb.scala 191:76 40:26]
  wire [19:0] _GEN_829 = _T_73 == 64'h1 ? paddr_1 : _GEN_729; // @[playground/src/noop/tlb.scala 191:76 40:26]
  wire [19:0] _GEN_830 = _T_73 == 64'h1 ? paddr_2 : _GEN_730; // @[playground/src/noop/tlb.scala 191:76 40:26]
  wire [19:0] _GEN_831 = _T_73 == 64'h1 ? paddr_3 : _GEN_731; // @[playground/src/noop/tlb.scala 191:76 40:26]
  wire [19:0] _GEN_832 = _T_73 == 64'h1 ? paddr_4 : _GEN_732; // @[playground/src/noop/tlb.scala 191:76 40:26]
  wire [19:0] _GEN_833 = _T_73 == 64'h1 ? paddr_5 : _GEN_733; // @[playground/src/noop/tlb.scala 191:76 40:26]
  wire [19:0] _GEN_834 = _T_73 == 64'h1 ? paddr_6 : _GEN_734; // @[playground/src/noop/tlb.scala 191:76 40:26]
  wire [19:0] _GEN_835 = _T_73 == 64'h1 ? paddr_7 : _GEN_735; // @[playground/src/noop/tlb.scala 191:76 40:26]
  wire [19:0] _GEN_836 = _T_73 == 64'h1 ? paddr_8 : _GEN_736; // @[playground/src/noop/tlb.scala 191:76 40:26]
  wire [19:0] _GEN_837 = _T_73 == 64'h1 ? paddr_9 : _GEN_737; // @[playground/src/noop/tlb.scala 191:76 40:26]
  wire [19:0] _GEN_838 = _T_73 == 64'h1 ? paddr_10 : _GEN_738; // @[playground/src/noop/tlb.scala 191:76 40:26]
  wire [19:0] _GEN_839 = _T_73 == 64'h1 ? paddr_11 : _GEN_739; // @[playground/src/noop/tlb.scala 191:76 40:26]
  wire [19:0] _GEN_840 = _T_73 == 64'h1 ? paddr_12 : _GEN_740; // @[playground/src/noop/tlb.scala 191:76 40:26]
  wire [19:0] _GEN_841 = _T_73 == 64'h1 ? paddr_13 : _GEN_741; // @[playground/src/noop/tlb.scala 191:76 40:26]
  wire [19:0] _GEN_842 = _T_73 == 64'h1 ? paddr_14 : _GEN_742; // @[playground/src/noop/tlb.scala 191:76 40:26]
  wire [19:0] _GEN_843 = _T_73 == 64'h1 ? paddr_15 : _GEN_743; // @[playground/src/noop/tlb.scala 191:76 40:26]
  wire [31:0] _GEN_844 = _T_73 == 64'h1 ? pte_addr_0 : _GEN_744; // @[playground/src/noop/tlb.scala 191:76 42:30]
  wire [31:0] _GEN_845 = _T_73 == 64'h1 ? pte_addr_1 : _GEN_745; // @[playground/src/noop/tlb.scala 191:76 42:30]
  wire [31:0] _GEN_846 = _T_73 == 64'h1 ? pte_addr_2 : _GEN_746; // @[playground/src/noop/tlb.scala 191:76 42:30]
  wire [31:0] _GEN_847 = _T_73 == 64'h1 ? pte_addr_3 : _GEN_747; // @[playground/src/noop/tlb.scala 191:76 42:30]
  wire [31:0] _GEN_848 = _T_73 == 64'h1 ? pte_addr_4 : _GEN_748; // @[playground/src/noop/tlb.scala 191:76 42:30]
  wire [31:0] _GEN_849 = _T_73 == 64'h1 ? pte_addr_5 : _GEN_749; // @[playground/src/noop/tlb.scala 191:76 42:30]
  wire [31:0] _GEN_850 = _T_73 == 64'h1 ? pte_addr_6 : _GEN_750; // @[playground/src/noop/tlb.scala 191:76 42:30]
  wire [31:0] _GEN_851 = _T_73 == 64'h1 ? pte_addr_7 : _GEN_751; // @[playground/src/noop/tlb.scala 191:76 42:30]
  wire [31:0] _GEN_852 = _T_73 == 64'h1 ? pte_addr_8 : _GEN_752; // @[playground/src/noop/tlb.scala 191:76 42:30]
  wire [31:0] _GEN_853 = _T_73 == 64'h1 ? pte_addr_9 : _GEN_753; // @[playground/src/noop/tlb.scala 191:76 42:30]
  wire [31:0] _GEN_854 = _T_73 == 64'h1 ? pte_addr_10 : _GEN_754; // @[playground/src/noop/tlb.scala 191:76 42:30]
  wire [31:0] _GEN_855 = _T_73 == 64'h1 ? pte_addr_11 : _GEN_755; // @[playground/src/noop/tlb.scala 191:76 42:30]
  wire [31:0] _GEN_856 = _T_73 == 64'h1 ? pte_addr_12 : _GEN_756; // @[playground/src/noop/tlb.scala 191:76 42:30]
  wire [31:0] _GEN_857 = _T_73 == 64'h1 ? pte_addr_13 : _GEN_757; // @[playground/src/noop/tlb.scala 191:76 42:30]
  wire [31:0] _GEN_858 = _T_73 == 64'h1 ? pte_addr_14 : _GEN_758; // @[playground/src/noop/tlb.scala 191:76 42:30]
  wire [31:0] _GEN_859 = _T_73 == 64'h1 ? pte_addr_15 : _GEN_759; // @[playground/src/noop/tlb.scala 191:76 42:30]
  wire [1:0] _GEN_860 = _T_73 == 64'h1 ? pte_level_0 : _GEN_760; // @[playground/src/noop/tlb.scala 191:76 43:30]
  wire [1:0] _GEN_861 = _T_73 == 64'h1 ? pte_level_1 : _GEN_761; // @[playground/src/noop/tlb.scala 191:76 43:30]
  wire [1:0] _GEN_862 = _T_73 == 64'h1 ? pte_level_2 : _GEN_762; // @[playground/src/noop/tlb.scala 191:76 43:30]
  wire [1:0] _GEN_863 = _T_73 == 64'h1 ? pte_level_3 : _GEN_763; // @[playground/src/noop/tlb.scala 191:76 43:30]
  wire [1:0] _GEN_864 = _T_73 == 64'h1 ? pte_level_4 : _GEN_764; // @[playground/src/noop/tlb.scala 191:76 43:30]
  wire [1:0] _GEN_865 = _T_73 == 64'h1 ? pte_level_5 : _GEN_765; // @[playground/src/noop/tlb.scala 191:76 43:30]
  wire [1:0] _GEN_866 = _T_73 == 64'h1 ? pte_level_6 : _GEN_766; // @[playground/src/noop/tlb.scala 191:76 43:30]
  wire [1:0] _GEN_867 = _T_73 == 64'h1 ? pte_level_7 : _GEN_767; // @[playground/src/noop/tlb.scala 191:76 43:30]
  wire [1:0] _GEN_868 = _T_73 == 64'h1 ? pte_level_8 : _GEN_768; // @[playground/src/noop/tlb.scala 191:76 43:30]
  wire [1:0] _GEN_869 = _T_73 == 64'h1 ? pte_level_9 : _GEN_769; // @[playground/src/noop/tlb.scala 191:76 43:30]
  wire [1:0] _GEN_870 = _T_73 == 64'h1 ? pte_level_10 : _GEN_770; // @[playground/src/noop/tlb.scala 191:76 43:30]
  wire [1:0] _GEN_871 = _T_73 == 64'h1 ? pte_level_11 : _GEN_771; // @[playground/src/noop/tlb.scala 191:76 43:30]
  wire [1:0] _GEN_872 = _T_73 == 64'h1 ? pte_level_12 : _GEN_772; // @[playground/src/noop/tlb.scala 191:76 43:30]
  wire [1:0] _GEN_873 = _T_73 == 64'h1 ? pte_level_13 : _GEN_773; // @[playground/src/noop/tlb.scala 191:76 43:30]
  wire [1:0] _GEN_874 = _T_73 == 64'h1 ? pte_level_14 : _GEN_774; // @[playground/src/noop/tlb.scala 191:76 43:30]
  wire [1:0] _GEN_875 = _T_73 == 64'h1 ? pte_level_15 : _GEN_775; // @[playground/src/noop/tlb.scala 191:76 43:30]
  wire [9:0] _GEN_876 = _T_73 == 64'h1 ? info_0 : _GEN_776; // @[playground/src/noop/tlb.scala 191:76 41:26]
  wire [9:0] _GEN_877 = _T_73 == 64'h1 ? info_1 : _GEN_777; // @[playground/src/noop/tlb.scala 191:76 41:26]
  wire [9:0] _GEN_878 = _T_73 == 64'h1 ? info_2 : _GEN_778; // @[playground/src/noop/tlb.scala 191:76 41:26]
  wire [9:0] _GEN_879 = _T_73 == 64'h1 ? info_3 : _GEN_779; // @[playground/src/noop/tlb.scala 191:76 41:26]
  wire [9:0] _GEN_880 = _T_73 == 64'h1 ? info_4 : _GEN_780; // @[playground/src/noop/tlb.scala 191:76 41:26]
  wire [9:0] _GEN_881 = _T_73 == 64'h1 ? info_5 : _GEN_781; // @[playground/src/noop/tlb.scala 191:76 41:26]
  wire [9:0] _GEN_882 = _T_73 == 64'h1 ? info_6 : _GEN_782; // @[playground/src/noop/tlb.scala 191:76 41:26]
  wire [9:0] _GEN_883 = _T_73 == 64'h1 ? info_7 : _GEN_783; // @[playground/src/noop/tlb.scala 191:76 41:26]
  wire [9:0] _GEN_884 = _T_73 == 64'h1 ? info_8 : _GEN_784; // @[playground/src/noop/tlb.scala 191:76 41:26]
  wire [9:0] _GEN_885 = _T_73 == 64'h1 ? info_9 : _GEN_785; // @[playground/src/noop/tlb.scala 191:76 41:26]
  wire [9:0] _GEN_886 = _T_73 == 64'h1 ? info_10 : _GEN_786; // @[playground/src/noop/tlb.scala 191:76 41:26]
  wire [9:0] _GEN_887 = _T_73 == 64'h1 ? info_11 : _GEN_787; // @[playground/src/noop/tlb.scala 191:76 41:26]
  wire [9:0] _GEN_888 = _T_73 == 64'h1 ? info_12 : _GEN_788; // @[playground/src/noop/tlb.scala 191:76 41:26]
  wire [9:0] _GEN_889 = _T_73 == 64'h1 ? info_13 : _GEN_789; // @[playground/src/noop/tlb.scala 191:76 41:26]
  wire [9:0] _GEN_890 = _T_73 == 64'h1 ? info_14 : _GEN_790; // @[playground/src/noop/tlb.scala 191:76 41:26]
  wire [9:0] _GEN_891 = _T_73 == 64'h1 ? info_15 : _GEN_791; // @[playground/src/noop/tlb.scala 191:76 41:26]
  wire [1:0] _GEN_892 = io_dcacheRW_rvalid ? _GEN_792 : state; // @[playground/src/noop/tlb.scala 190:41 84:24]
  wire  _GEN_893 = io_dcacheRW_rvalid ? _GEN_793 : _GEN_151; // @[playground/src/noop/tlb.scala 190:41]
  wire [55:0] _GEN_894 = io_dcacheRW_rvalid ? _GEN_794 : {{24'd0}, pte_addr_r}; // @[playground/src/noop/tlb.scala 190:41 47:30]
  wire [4:0] _GEN_895 = io_dcacheRW_rvalid ? _GEN_795 : _GEN_297; // @[playground/src/noop/tlb.scala 190:41]
  wire [51:0] _GEN_896 = io_dcacheRW_rvalid ? _GEN_796 : tag_0; // @[playground/src/noop/tlb.scala 190:41 39:26]
  wire [51:0] _GEN_897 = io_dcacheRW_rvalid ? _GEN_797 : tag_1; // @[playground/src/noop/tlb.scala 190:41 39:26]
  wire [51:0] _GEN_898 = io_dcacheRW_rvalid ? _GEN_798 : tag_2; // @[playground/src/noop/tlb.scala 190:41 39:26]
  wire [51:0] _GEN_899 = io_dcacheRW_rvalid ? _GEN_799 : tag_3; // @[playground/src/noop/tlb.scala 190:41 39:26]
  wire [51:0] _GEN_900 = io_dcacheRW_rvalid ? _GEN_800 : tag_4; // @[playground/src/noop/tlb.scala 190:41 39:26]
  wire [51:0] _GEN_901 = io_dcacheRW_rvalid ? _GEN_801 : tag_5; // @[playground/src/noop/tlb.scala 190:41 39:26]
  wire [51:0] _GEN_902 = io_dcacheRW_rvalid ? _GEN_802 : tag_6; // @[playground/src/noop/tlb.scala 190:41 39:26]
  wire [51:0] _GEN_903 = io_dcacheRW_rvalid ? _GEN_803 : tag_7; // @[playground/src/noop/tlb.scala 190:41 39:26]
  wire [51:0] _GEN_904 = io_dcacheRW_rvalid ? _GEN_804 : tag_8; // @[playground/src/noop/tlb.scala 190:41 39:26]
  wire [51:0] _GEN_905 = io_dcacheRW_rvalid ? _GEN_805 : tag_9; // @[playground/src/noop/tlb.scala 190:41 39:26]
  wire [51:0] _GEN_906 = io_dcacheRW_rvalid ? _GEN_806 : tag_10; // @[playground/src/noop/tlb.scala 190:41 39:26]
  wire [51:0] _GEN_907 = io_dcacheRW_rvalid ? _GEN_807 : tag_11; // @[playground/src/noop/tlb.scala 190:41 39:26]
  wire [51:0] _GEN_908 = io_dcacheRW_rvalid ? _GEN_808 : tag_12; // @[playground/src/noop/tlb.scala 190:41 39:26]
  wire [51:0] _GEN_909 = io_dcacheRW_rvalid ? _GEN_809 : tag_13; // @[playground/src/noop/tlb.scala 190:41 39:26]
  wire [51:0] _GEN_910 = io_dcacheRW_rvalid ? _GEN_810 : tag_14; // @[playground/src/noop/tlb.scala 190:41 39:26]
  wire [51:0] _GEN_911 = io_dcacheRW_rvalid ? _GEN_811 : tag_15; // @[playground/src/noop/tlb.scala 190:41 39:26]
  wire  _GEN_912 = io_dcacheRW_rvalid ? _GEN_812 : _GEN_130; // @[playground/src/noop/tlb.scala 190:41]
  wire  _GEN_913 = io_dcacheRW_rvalid ? _GEN_813 : _GEN_131; // @[playground/src/noop/tlb.scala 190:41]
  wire  _GEN_914 = io_dcacheRW_rvalid ? _GEN_814 : _GEN_132; // @[playground/src/noop/tlb.scala 190:41]
  wire  _GEN_915 = io_dcacheRW_rvalid ? _GEN_815 : _GEN_133; // @[playground/src/noop/tlb.scala 190:41]
  wire  _GEN_916 = io_dcacheRW_rvalid ? _GEN_816 : _GEN_134; // @[playground/src/noop/tlb.scala 190:41]
  wire  _GEN_917 = io_dcacheRW_rvalid ? _GEN_817 : _GEN_135; // @[playground/src/noop/tlb.scala 190:41]
  wire  _GEN_918 = io_dcacheRW_rvalid ? _GEN_818 : _GEN_136; // @[playground/src/noop/tlb.scala 190:41]
  wire  _GEN_919 = io_dcacheRW_rvalid ? _GEN_819 : _GEN_137; // @[playground/src/noop/tlb.scala 190:41]
  wire  _GEN_920 = io_dcacheRW_rvalid ? _GEN_820 : _GEN_138; // @[playground/src/noop/tlb.scala 190:41]
  wire  _GEN_921 = io_dcacheRW_rvalid ? _GEN_821 : _GEN_139; // @[playground/src/noop/tlb.scala 190:41]
  wire  _GEN_922 = io_dcacheRW_rvalid ? _GEN_822 : _GEN_140; // @[playground/src/noop/tlb.scala 190:41]
  wire  _GEN_923 = io_dcacheRW_rvalid ? _GEN_823 : _GEN_141; // @[playground/src/noop/tlb.scala 190:41]
  wire  _GEN_924 = io_dcacheRW_rvalid ? _GEN_824 : _GEN_142; // @[playground/src/noop/tlb.scala 190:41]
  wire  _GEN_925 = io_dcacheRW_rvalid ? _GEN_825 : _GEN_143; // @[playground/src/noop/tlb.scala 190:41]
  wire  _GEN_926 = io_dcacheRW_rvalid ? _GEN_826 : _GEN_144; // @[playground/src/noop/tlb.scala 190:41]
  wire  _GEN_927 = io_dcacheRW_rvalid ? _GEN_827 : _GEN_145; // @[playground/src/noop/tlb.scala 190:41]
  wire [19:0] _GEN_928 = io_dcacheRW_rvalid ? _GEN_828 : paddr_0; // @[playground/src/noop/tlb.scala 190:41 40:26]
  wire [19:0] _GEN_929 = io_dcacheRW_rvalid ? _GEN_829 : paddr_1; // @[playground/src/noop/tlb.scala 190:41 40:26]
  wire [19:0] _GEN_930 = io_dcacheRW_rvalid ? _GEN_830 : paddr_2; // @[playground/src/noop/tlb.scala 190:41 40:26]
  wire [19:0] _GEN_931 = io_dcacheRW_rvalid ? _GEN_831 : paddr_3; // @[playground/src/noop/tlb.scala 190:41 40:26]
  wire [19:0] _GEN_932 = io_dcacheRW_rvalid ? _GEN_832 : paddr_4; // @[playground/src/noop/tlb.scala 190:41 40:26]
  wire [19:0] _GEN_933 = io_dcacheRW_rvalid ? _GEN_833 : paddr_5; // @[playground/src/noop/tlb.scala 190:41 40:26]
  wire [19:0] _GEN_934 = io_dcacheRW_rvalid ? _GEN_834 : paddr_6; // @[playground/src/noop/tlb.scala 190:41 40:26]
  wire [19:0] _GEN_935 = io_dcacheRW_rvalid ? _GEN_835 : paddr_7; // @[playground/src/noop/tlb.scala 190:41 40:26]
  wire [19:0] _GEN_936 = io_dcacheRW_rvalid ? _GEN_836 : paddr_8; // @[playground/src/noop/tlb.scala 190:41 40:26]
  wire [19:0] _GEN_937 = io_dcacheRW_rvalid ? _GEN_837 : paddr_9; // @[playground/src/noop/tlb.scala 190:41 40:26]
  wire [19:0] _GEN_938 = io_dcacheRW_rvalid ? _GEN_838 : paddr_10; // @[playground/src/noop/tlb.scala 190:41 40:26]
  wire [19:0] _GEN_939 = io_dcacheRW_rvalid ? _GEN_839 : paddr_11; // @[playground/src/noop/tlb.scala 190:41 40:26]
  wire [19:0] _GEN_940 = io_dcacheRW_rvalid ? _GEN_840 : paddr_12; // @[playground/src/noop/tlb.scala 190:41 40:26]
  wire [19:0] _GEN_941 = io_dcacheRW_rvalid ? _GEN_841 : paddr_13; // @[playground/src/noop/tlb.scala 190:41 40:26]
  wire [19:0] _GEN_942 = io_dcacheRW_rvalid ? _GEN_842 : paddr_14; // @[playground/src/noop/tlb.scala 190:41 40:26]
  wire [19:0] _GEN_943 = io_dcacheRW_rvalid ? _GEN_843 : paddr_15; // @[playground/src/noop/tlb.scala 190:41 40:26]
  wire [31:0] _GEN_944 = io_dcacheRW_rvalid ? _GEN_844 : pte_addr_0; // @[playground/src/noop/tlb.scala 190:41 42:30]
  wire [31:0] _GEN_945 = io_dcacheRW_rvalid ? _GEN_845 : pte_addr_1; // @[playground/src/noop/tlb.scala 190:41 42:30]
  wire [31:0] _GEN_946 = io_dcacheRW_rvalid ? _GEN_846 : pte_addr_2; // @[playground/src/noop/tlb.scala 190:41 42:30]
  wire [31:0] _GEN_947 = io_dcacheRW_rvalid ? _GEN_847 : pte_addr_3; // @[playground/src/noop/tlb.scala 190:41 42:30]
  wire [31:0] _GEN_948 = io_dcacheRW_rvalid ? _GEN_848 : pte_addr_4; // @[playground/src/noop/tlb.scala 190:41 42:30]
  wire [31:0] _GEN_949 = io_dcacheRW_rvalid ? _GEN_849 : pte_addr_5; // @[playground/src/noop/tlb.scala 190:41 42:30]
  wire [31:0] _GEN_950 = io_dcacheRW_rvalid ? _GEN_850 : pte_addr_6; // @[playground/src/noop/tlb.scala 190:41 42:30]
  wire [31:0] _GEN_951 = io_dcacheRW_rvalid ? _GEN_851 : pte_addr_7; // @[playground/src/noop/tlb.scala 190:41 42:30]
  wire [31:0] _GEN_952 = io_dcacheRW_rvalid ? _GEN_852 : pte_addr_8; // @[playground/src/noop/tlb.scala 190:41 42:30]
  wire [31:0] _GEN_953 = io_dcacheRW_rvalid ? _GEN_853 : pte_addr_9; // @[playground/src/noop/tlb.scala 190:41 42:30]
  wire [31:0] _GEN_954 = io_dcacheRW_rvalid ? _GEN_854 : pte_addr_10; // @[playground/src/noop/tlb.scala 190:41 42:30]
  wire [31:0] _GEN_955 = io_dcacheRW_rvalid ? _GEN_855 : pte_addr_11; // @[playground/src/noop/tlb.scala 190:41 42:30]
  wire [31:0] _GEN_956 = io_dcacheRW_rvalid ? _GEN_856 : pte_addr_12; // @[playground/src/noop/tlb.scala 190:41 42:30]
  wire [31:0] _GEN_957 = io_dcacheRW_rvalid ? _GEN_857 : pte_addr_13; // @[playground/src/noop/tlb.scala 190:41 42:30]
  wire [31:0] _GEN_958 = io_dcacheRW_rvalid ? _GEN_858 : pte_addr_14; // @[playground/src/noop/tlb.scala 190:41 42:30]
  wire [31:0] _GEN_959 = io_dcacheRW_rvalid ? _GEN_859 : pte_addr_15; // @[playground/src/noop/tlb.scala 190:41 42:30]
  wire [1:0] _GEN_960 = io_dcacheRW_rvalid ? _GEN_860 : pte_level_0; // @[playground/src/noop/tlb.scala 190:41 43:30]
  wire [1:0] _GEN_961 = io_dcacheRW_rvalid ? _GEN_861 : pte_level_1; // @[playground/src/noop/tlb.scala 190:41 43:30]
  wire [1:0] _GEN_962 = io_dcacheRW_rvalid ? _GEN_862 : pte_level_2; // @[playground/src/noop/tlb.scala 190:41 43:30]
  wire [1:0] _GEN_963 = io_dcacheRW_rvalid ? _GEN_863 : pte_level_3; // @[playground/src/noop/tlb.scala 190:41 43:30]
  wire [1:0] _GEN_964 = io_dcacheRW_rvalid ? _GEN_864 : pte_level_4; // @[playground/src/noop/tlb.scala 190:41 43:30]
  wire [1:0] _GEN_965 = io_dcacheRW_rvalid ? _GEN_865 : pte_level_5; // @[playground/src/noop/tlb.scala 190:41 43:30]
  wire [1:0] _GEN_966 = io_dcacheRW_rvalid ? _GEN_866 : pte_level_6; // @[playground/src/noop/tlb.scala 190:41 43:30]
  wire [1:0] _GEN_967 = io_dcacheRW_rvalid ? _GEN_867 : pte_level_7; // @[playground/src/noop/tlb.scala 190:41 43:30]
  wire [1:0] _GEN_968 = io_dcacheRW_rvalid ? _GEN_868 : pte_level_8; // @[playground/src/noop/tlb.scala 190:41 43:30]
  wire [1:0] _GEN_969 = io_dcacheRW_rvalid ? _GEN_869 : pte_level_9; // @[playground/src/noop/tlb.scala 190:41 43:30]
  wire [1:0] _GEN_970 = io_dcacheRW_rvalid ? _GEN_870 : pte_level_10; // @[playground/src/noop/tlb.scala 190:41 43:30]
  wire [1:0] _GEN_971 = io_dcacheRW_rvalid ? _GEN_871 : pte_level_11; // @[playground/src/noop/tlb.scala 190:41 43:30]
  wire [1:0] _GEN_972 = io_dcacheRW_rvalid ? _GEN_872 : pte_level_12; // @[playground/src/noop/tlb.scala 190:41 43:30]
  wire [1:0] _GEN_973 = io_dcacheRW_rvalid ? _GEN_873 : pte_level_13; // @[playground/src/noop/tlb.scala 190:41 43:30]
  wire [1:0] _GEN_974 = io_dcacheRW_rvalid ? _GEN_874 : pte_level_14; // @[playground/src/noop/tlb.scala 190:41 43:30]
  wire [1:0] _GEN_975 = io_dcacheRW_rvalid ? _GEN_875 : pte_level_15; // @[playground/src/noop/tlb.scala 190:41 43:30]
  wire [9:0] _GEN_976 = io_dcacheRW_rvalid ? _GEN_876 : info_0; // @[playground/src/noop/tlb.scala 190:41 41:26]
  wire [9:0] _GEN_977 = io_dcacheRW_rvalid ? _GEN_877 : info_1; // @[playground/src/noop/tlb.scala 190:41 41:26]
  wire [9:0] _GEN_978 = io_dcacheRW_rvalid ? _GEN_878 : info_2; // @[playground/src/noop/tlb.scala 190:41 41:26]
  wire [9:0] _GEN_979 = io_dcacheRW_rvalid ? _GEN_879 : info_3; // @[playground/src/noop/tlb.scala 190:41 41:26]
  wire [9:0] _GEN_980 = io_dcacheRW_rvalid ? _GEN_880 : info_4; // @[playground/src/noop/tlb.scala 190:41 41:26]
  wire [9:0] _GEN_981 = io_dcacheRW_rvalid ? _GEN_881 : info_5; // @[playground/src/noop/tlb.scala 190:41 41:26]
  wire [9:0] _GEN_982 = io_dcacheRW_rvalid ? _GEN_882 : info_6; // @[playground/src/noop/tlb.scala 190:41 41:26]
  wire [9:0] _GEN_983 = io_dcacheRW_rvalid ? _GEN_883 : info_7; // @[playground/src/noop/tlb.scala 190:41 41:26]
  wire [9:0] _GEN_984 = io_dcacheRW_rvalid ? _GEN_884 : info_8; // @[playground/src/noop/tlb.scala 190:41 41:26]
  wire [9:0] _GEN_985 = io_dcacheRW_rvalid ? _GEN_885 : info_9; // @[playground/src/noop/tlb.scala 190:41 41:26]
  wire [9:0] _GEN_986 = io_dcacheRW_rvalid ? _GEN_886 : info_10; // @[playground/src/noop/tlb.scala 190:41 41:26]
  wire [9:0] _GEN_987 = io_dcacheRW_rvalid ? _GEN_887 : info_11; // @[playground/src/noop/tlb.scala 190:41 41:26]
  wire [9:0] _GEN_988 = io_dcacheRW_rvalid ? _GEN_888 : info_12; // @[playground/src/noop/tlb.scala 190:41 41:26]
  wire [9:0] _GEN_989 = io_dcacheRW_rvalid ? _GEN_889 : info_13; // @[playground/src/noop/tlb.scala 190:41 41:26]
  wire [9:0] _GEN_990 = io_dcacheRW_rvalid ? _GEN_890 : info_14; // @[playground/src/noop/tlb.scala 190:41 41:26]
  wire [9:0] _GEN_991 = io_dcacheRW_rvalid ? _GEN_891 : info_15; // @[playground/src/noop/tlb.scala 190:41 41:26]
  wire [4:0] _GEN_992 = 2'h1 == state ? _GEN_895 : dc_mode_r; // @[playground/src/noop/tlb.scala 136:22 49:30]
  wire [7:0] _GEN_993 = 2'h1 == state ? _GEN_298 : offset; // @[playground/src/noop/tlb.scala 136:22 131:26]
  wire [1:0] _GEN_994 = 2'h1 == state ? _GEN_299 : level; // @[playground/src/noop/tlb.scala 136:22 132:26]
  wire [1:0] _GEN_995 = 2'h1 == state ? _GEN_892 : state; // @[playground/src/noop/tlb.scala 136:22 84:24]
  wire  _GEN_996 = 2'h1 == state ? _GEN_893 : _GEN_151; // @[playground/src/noop/tlb.scala 136:22]
  wire [55:0] _GEN_997 = 2'h1 == state ? _GEN_894 : {{24'd0}, pte_addr_r}; // @[playground/src/noop/tlb.scala 136:22 47:30]
  wire [51:0] _GEN_998 = 2'h1 == state ? _GEN_896 : tag_0; // @[playground/src/noop/tlb.scala 136:22 39:26]
  wire [51:0] _GEN_999 = 2'h1 == state ? _GEN_897 : tag_1; // @[playground/src/noop/tlb.scala 136:22 39:26]
  wire [51:0] _GEN_1000 = 2'h1 == state ? _GEN_898 : tag_2; // @[playground/src/noop/tlb.scala 136:22 39:26]
  wire [51:0] _GEN_1001 = 2'h1 == state ? _GEN_899 : tag_3; // @[playground/src/noop/tlb.scala 136:22 39:26]
  wire [51:0] _GEN_1002 = 2'h1 == state ? _GEN_900 : tag_4; // @[playground/src/noop/tlb.scala 136:22 39:26]
  wire [51:0] _GEN_1003 = 2'h1 == state ? _GEN_901 : tag_5; // @[playground/src/noop/tlb.scala 136:22 39:26]
  wire [51:0] _GEN_1004 = 2'h1 == state ? _GEN_902 : tag_6; // @[playground/src/noop/tlb.scala 136:22 39:26]
  wire [51:0] _GEN_1005 = 2'h1 == state ? _GEN_903 : tag_7; // @[playground/src/noop/tlb.scala 136:22 39:26]
  wire [51:0] _GEN_1006 = 2'h1 == state ? _GEN_904 : tag_8; // @[playground/src/noop/tlb.scala 136:22 39:26]
  wire [51:0] _GEN_1007 = 2'h1 == state ? _GEN_905 : tag_9; // @[playground/src/noop/tlb.scala 136:22 39:26]
  wire [51:0] _GEN_1008 = 2'h1 == state ? _GEN_906 : tag_10; // @[playground/src/noop/tlb.scala 136:22 39:26]
  wire [51:0] _GEN_1009 = 2'h1 == state ? _GEN_907 : tag_11; // @[playground/src/noop/tlb.scala 136:22 39:26]
  wire [51:0] _GEN_1010 = 2'h1 == state ? _GEN_908 : tag_12; // @[playground/src/noop/tlb.scala 136:22 39:26]
  wire [51:0] _GEN_1011 = 2'h1 == state ? _GEN_909 : tag_13; // @[playground/src/noop/tlb.scala 136:22 39:26]
  wire [51:0] _GEN_1012 = 2'h1 == state ? _GEN_910 : tag_14; // @[playground/src/noop/tlb.scala 136:22 39:26]
  wire [51:0] _GEN_1013 = 2'h1 == state ? _GEN_911 : tag_15; // @[playground/src/noop/tlb.scala 136:22 39:26]
  wire  _GEN_1014 = 2'h1 == state ? _GEN_912 : _GEN_130; // @[playground/src/noop/tlb.scala 136:22]
  wire  _GEN_1015 = 2'h1 == state ? _GEN_913 : _GEN_131; // @[playground/src/noop/tlb.scala 136:22]
  wire  _GEN_1016 = 2'h1 == state ? _GEN_914 : _GEN_132; // @[playground/src/noop/tlb.scala 136:22]
  wire  _GEN_1017 = 2'h1 == state ? _GEN_915 : _GEN_133; // @[playground/src/noop/tlb.scala 136:22]
  wire  _GEN_1018 = 2'h1 == state ? _GEN_916 : _GEN_134; // @[playground/src/noop/tlb.scala 136:22]
  wire  _GEN_1019 = 2'h1 == state ? _GEN_917 : _GEN_135; // @[playground/src/noop/tlb.scala 136:22]
  wire  _GEN_1020 = 2'h1 == state ? _GEN_918 : _GEN_136; // @[playground/src/noop/tlb.scala 136:22]
  wire  _GEN_1021 = 2'h1 == state ? _GEN_919 : _GEN_137; // @[playground/src/noop/tlb.scala 136:22]
  wire  _GEN_1022 = 2'h1 == state ? _GEN_920 : _GEN_138; // @[playground/src/noop/tlb.scala 136:22]
  wire  _GEN_1023 = 2'h1 == state ? _GEN_921 : _GEN_139; // @[playground/src/noop/tlb.scala 136:22]
  wire  _GEN_1024 = 2'h1 == state ? _GEN_922 : _GEN_140; // @[playground/src/noop/tlb.scala 136:22]
  wire  _GEN_1025 = 2'h1 == state ? _GEN_923 : _GEN_141; // @[playground/src/noop/tlb.scala 136:22]
  wire  _GEN_1026 = 2'h1 == state ? _GEN_924 : _GEN_142; // @[playground/src/noop/tlb.scala 136:22]
  wire  _GEN_1027 = 2'h1 == state ? _GEN_925 : _GEN_143; // @[playground/src/noop/tlb.scala 136:22]
  wire  _GEN_1028 = 2'h1 == state ? _GEN_926 : _GEN_144; // @[playground/src/noop/tlb.scala 136:22]
  wire  _GEN_1029 = 2'h1 == state ? _GEN_927 : _GEN_145; // @[playground/src/noop/tlb.scala 136:22]
  wire [19:0] _GEN_1030 = 2'h1 == state ? _GEN_928 : paddr_0; // @[playground/src/noop/tlb.scala 136:22 40:26]
  wire [19:0] _GEN_1031 = 2'h1 == state ? _GEN_929 : paddr_1; // @[playground/src/noop/tlb.scala 136:22 40:26]
  wire [19:0] _GEN_1032 = 2'h1 == state ? _GEN_930 : paddr_2; // @[playground/src/noop/tlb.scala 136:22 40:26]
  wire [19:0] _GEN_1033 = 2'h1 == state ? _GEN_931 : paddr_3; // @[playground/src/noop/tlb.scala 136:22 40:26]
  wire [19:0] _GEN_1034 = 2'h1 == state ? _GEN_932 : paddr_4; // @[playground/src/noop/tlb.scala 136:22 40:26]
  wire [19:0] _GEN_1035 = 2'h1 == state ? _GEN_933 : paddr_5; // @[playground/src/noop/tlb.scala 136:22 40:26]
  wire [19:0] _GEN_1036 = 2'h1 == state ? _GEN_934 : paddr_6; // @[playground/src/noop/tlb.scala 136:22 40:26]
  wire [19:0] _GEN_1037 = 2'h1 == state ? _GEN_935 : paddr_7; // @[playground/src/noop/tlb.scala 136:22 40:26]
  wire [19:0] _GEN_1038 = 2'h1 == state ? _GEN_936 : paddr_8; // @[playground/src/noop/tlb.scala 136:22 40:26]
  wire [19:0] _GEN_1039 = 2'h1 == state ? _GEN_937 : paddr_9; // @[playground/src/noop/tlb.scala 136:22 40:26]
  wire [19:0] _GEN_1040 = 2'h1 == state ? _GEN_938 : paddr_10; // @[playground/src/noop/tlb.scala 136:22 40:26]
  wire [19:0] _GEN_1041 = 2'h1 == state ? _GEN_939 : paddr_11; // @[playground/src/noop/tlb.scala 136:22 40:26]
  wire [19:0] _GEN_1042 = 2'h1 == state ? _GEN_940 : paddr_12; // @[playground/src/noop/tlb.scala 136:22 40:26]
  wire [19:0] _GEN_1043 = 2'h1 == state ? _GEN_941 : paddr_13; // @[playground/src/noop/tlb.scala 136:22 40:26]
  wire [19:0] _GEN_1044 = 2'h1 == state ? _GEN_942 : paddr_14; // @[playground/src/noop/tlb.scala 136:22 40:26]
  wire [19:0] _GEN_1045 = 2'h1 == state ? _GEN_943 : paddr_15; // @[playground/src/noop/tlb.scala 136:22 40:26]
  wire [31:0] _GEN_1046 = 2'h1 == state ? _GEN_944 : pte_addr_0; // @[playground/src/noop/tlb.scala 136:22 42:30]
  wire [31:0] _GEN_1047 = 2'h1 == state ? _GEN_945 : pte_addr_1; // @[playground/src/noop/tlb.scala 136:22 42:30]
  wire [31:0] _GEN_1048 = 2'h1 == state ? _GEN_946 : pte_addr_2; // @[playground/src/noop/tlb.scala 136:22 42:30]
  wire [31:0] _GEN_1049 = 2'h1 == state ? _GEN_947 : pte_addr_3; // @[playground/src/noop/tlb.scala 136:22 42:30]
  wire [31:0] _GEN_1050 = 2'h1 == state ? _GEN_948 : pte_addr_4; // @[playground/src/noop/tlb.scala 136:22 42:30]
  wire [31:0] _GEN_1051 = 2'h1 == state ? _GEN_949 : pte_addr_5; // @[playground/src/noop/tlb.scala 136:22 42:30]
  wire [31:0] _GEN_1052 = 2'h1 == state ? _GEN_950 : pte_addr_6; // @[playground/src/noop/tlb.scala 136:22 42:30]
  wire [31:0] _GEN_1053 = 2'h1 == state ? _GEN_951 : pte_addr_7; // @[playground/src/noop/tlb.scala 136:22 42:30]
  wire [31:0] _GEN_1054 = 2'h1 == state ? _GEN_952 : pte_addr_8; // @[playground/src/noop/tlb.scala 136:22 42:30]
  wire [31:0] _GEN_1055 = 2'h1 == state ? _GEN_953 : pte_addr_9; // @[playground/src/noop/tlb.scala 136:22 42:30]
  wire [31:0] _GEN_1056 = 2'h1 == state ? _GEN_954 : pte_addr_10; // @[playground/src/noop/tlb.scala 136:22 42:30]
  wire [31:0] _GEN_1057 = 2'h1 == state ? _GEN_955 : pte_addr_11; // @[playground/src/noop/tlb.scala 136:22 42:30]
  wire [31:0] _GEN_1058 = 2'h1 == state ? _GEN_956 : pte_addr_12; // @[playground/src/noop/tlb.scala 136:22 42:30]
  wire [31:0] _GEN_1059 = 2'h1 == state ? _GEN_957 : pte_addr_13; // @[playground/src/noop/tlb.scala 136:22 42:30]
  wire [31:0] _GEN_1060 = 2'h1 == state ? _GEN_958 : pte_addr_14; // @[playground/src/noop/tlb.scala 136:22 42:30]
  wire [31:0] _GEN_1061 = 2'h1 == state ? _GEN_959 : pte_addr_15; // @[playground/src/noop/tlb.scala 136:22 42:30]
  wire [1:0] _GEN_1062 = 2'h1 == state ? _GEN_960 : pte_level_0; // @[playground/src/noop/tlb.scala 136:22 43:30]
  wire [1:0] _GEN_1063 = 2'h1 == state ? _GEN_961 : pte_level_1; // @[playground/src/noop/tlb.scala 136:22 43:30]
  wire [1:0] _GEN_1064 = 2'h1 == state ? _GEN_962 : pte_level_2; // @[playground/src/noop/tlb.scala 136:22 43:30]
  wire [1:0] _GEN_1065 = 2'h1 == state ? _GEN_963 : pte_level_3; // @[playground/src/noop/tlb.scala 136:22 43:30]
  wire [1:0] _GEN_1066 = 2'h1 == state ? _GEN_964 : pte_level_4; // @[playground/src/noop/tlb.scala 136:22 43:30]
  wire [1:0] _GEN_1067 = 2'h1 == state ? _GEN_965 : pte_level_5; // @[playground/src/noop/tlb.scala 136:22 43:30]
  wire [1:0] _GEN_1068 = 2'h1 == state ? _GEN_966 : pte_level_6; // @[playground/src/noop/tlb.scala 136:22 43:30]
  wire [1:0] _GEN_1069 = 2'h1 == state ? _GEN_967 : pte_level_7; // @[playground/src/noop/tlb.scala 136:22 43:30]
  wire [1:0] _GEN_1070 = 2'h1 == state ? _GEN_968 : pte_level_8; // @[playground/src/noop/tlb.scala 136:22 43:30]
  wire [1:0] _GEN_1071 = 2'h1 == state ? _GEN_969 : pte_level_9; // @[playground/src/noop/tlb.scala 136:22 43:30]
  wire [1:0] _GEN_1072 = 2'h1 == state ? _GEN_970 : pte_level_10; // @[playground/src/noop/tlb.scala 136:22 43:30]
  wire [1:0] _GEN_1073 = 2'h1 == state ? _GEN_971 : pte_level_11; // @[playground/src/noop/tlb.scala 136:22 43:30]
  wire [1:0] _GEN_1074 = 2'h1 == state ? _GEN_972 : pte_level_12; // @[playground/src/noop/tlb.scala 136:22 43:30]
  wire [1:0] _GEN_1075 = 2'h1 == state ? _GEN_973 : pte_level_13; // @[playground/src/noop/tlb.scala 136:22 43:30]
  wire [1:0] _GEN_1076 = 2'h1 == state ? _GEN_974 : pte_level_14; // @[playground/src/noop/tlb.scala 136:22 43:30]
  wire [1:0] _GEN_1077 = 2'h1 == state ? _GEN_975 : pte_level_15; // @[playground/src/noop/tlb.scala 136:22 43:30]
  wire [9:0] _GEN_1078 = 2'h1 == state ? _GEN_976 : info_0; // @[playground/src/noop/tlb.scala 136:22 41:26]
  wire [9:0] _GEN_1079 = 2'h1 == state ? _GEN_977 : info_1; // @[playground/src/noop/tlb.scala 136:22 41:26]
  wire [9:0] _GEN_1080 = 2'h1 == state ? _GEN_978 : info_2; // @[playground/src/noop/tlb.scala 136:22 41:26]
  wire [9:0] _GEN_1081 = 2'h1 == state ? _GEN_979 : info_3; // @[playground/src/noop/tlb.scala 136:22 41:26]
  wire [9:0] _GEN_1082 = 2'h1 == state ? _GEN_980 : info_4; // @[playground/src/noop/tlb.scala 136:22 41:26]
  wire [9:0] _GEN_1083 = 2'h1 == state ? _GEN_981 : info_5; // @[playground/src/noop/tlb.scala 136:22 41:26]
  wire [9:0] _GEN_1084 = 2'h1 == state ? _GEN_982 : info_6; // @[playground/src/noop/tlb.scala 136:22 41:26]
  wire [9:0] _GEN_1085 = 2'h1 == state ? _GEN_983 : info_7; // @[playground/src/noop/tlb.scala 136:22 41:26]
  wire [9:0] _GEN_1086 = 2'h1 == state ? _GEN_984 : info_8; // @[playground/src/noop/tlb.scala 136:22 41:26]
  wire [9:0] _GEN_1087 = 2'h1 == state ? _GEN_985 : info_9; // @[playground/src/noop/tlb.scala 136:22 41:26]
  wire [9:0] _GEN_1088 = 2'h1 == state ? _GEN_986 : info_10; // @[playground/src/noop/tlb.scala 136:22 41:26]
  wire [9:0] _GEN_1089 = 2'h1 == state ? _GEN_987 : info_11; // @[playground/src/noop/tlb.scala 136:22 41:26]
  wire [9:0] _GEN_1090 = 2'h1 == state ? _GEN_988 : info_12; // @[playground/src/noop/tlb.scala 136:22 41:26]
  wire [9:0] _GEN_1091 = 2'h1 == state ? _GEN_989 : info_13; // @[playground/src/noop/tlb.scala 136:22 41:26]
  wire [9:0] _GEN_1092 = 2'h1 == state ? _GEN_990 : info_14; // @[playground/src/noop/tlb.scala 136:22 41:26]
  wire [9:0] _GEN_1093 = 2'h1 == state ? _GEN_991 : info_15; // @[playground/src/noop/tlb.scala 136:22 41:26]
  wire [55:0] _GEN_1100 = 2'h3 == state ? {{24'd0}, pte_addr_r} : _GEN_997; // @[playground/src/noop/tlb.scala 136:22 47:30]
  wire [63:0] _GEN_1202 = 2'h0 == state ? _GEN_268 : {{32'd0}, out_paddr_r}; // @[playground/src/noop/tlb.scala 136:22 52:30]
  wire [55:0] _GEN_1205 = 2'h0 == state ? _GEN_271 : _GEN_1100; // @[playground/src/noop/tlb.scala 136:22]
  wire [63:0] _GEN_1312 = is_Sv39 | state != 2'h0 ? _GEN_1202 : io_va2pa_vaddr; // @[playground/src/noop/tlb.scala 135:37 233:21]
  wire [55:0] _GEN_1315 = is_Sv39 | state != 2'h0 ? _GEN_1205 : {{24'd0}, pte_addr_r}; // @[playground/src/noop/tlb.scala 135:37 47:30]
  wire [55:0] _GEN_1418 = reset ? 56'h0 : _GEN_1315; // @[playground/src/noop/tlb.scala 47:{30,30}]
  wire [63:0] _GEN_1419 = reset ? 64'h0 : _GEN_1312; // @[playground/src/noop/tlb.scala 52:{30,30}]
  MaxPeriodFibonacciLFSR_2 select_prng ( // @[src/main/scala/chisel3/util/random/PRNG.scala 91:22]
    .clock(select_prng_clock),
    .reset(select_prng_reset),
    .io_out_0(select_prng_io_out_0),
    .io_out_1(select_prng_io_out_1),
    .io_out_2(select_prng_io_out_2),
    .io_out_3(select_prng_io_out_3)
  );
  assign io_va2pa_ready = io_va2pa_vvalid & _T_50 & ~io_flush & ~flush_r; // @[playground/src/noop/tlb.scala 98:74]
  assign io_va2pa_paddr = out_paddr_r; // @[playground/src/noop/tlb.scala 113:20]
  assign io_va2pa_pvalid = out_valid_r; // @[playground/src/noop/tlb.scala 114:21]
  assign io_va2pa_tlb_excep_cause = out_excep_r_cause; // @[playground/src/noop/tlb.scala 115:24]
  assign io_va2pa_tlb_excep_tval = out_excep_r_tval; // @[playground/src/noop/tlb.scala 115:24]
  assign io_va2pa_tlb_excep_en = out_excep_r_en; // @[playground/src/noop/tlb.scala 115:24]
  assign io_dcacheRW_addr = pte_addr_r; // @[playground/src/noop/tlb.scala 117:22]
  assign io_dcacheRW_wdata = wpte_data_r; // @[playground/src/noop/tlb.scala 118:23]
  assign io_dcacheRW_dc_mode = dc_mode_r; // @[playground/src/noop/tlb.scala 119:25]
  assign select_prng_clock = clock;
  assign select_prng_reset = reset;
  always @(posedge clock) begin
    if (reset) begin // @[playground/src/noop/tlb.scala 39:26]
      tag_0 <= 52'h0; // @[playground/src/noop/tlb.scala 39:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (!(2'h0 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
        if (!(2'h3 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
          tag_0 <= _GEN_998;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 39:26]
      tag_1 <= 52'h0; // @[playground/src/noop/tlb.scala 39:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (!(2'h0 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
        if (!(2'h3 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
          tag_1 <= _GEN_999;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 39:26]
      tag_2 <= 52'h0; // @[playground/src/noop/tlb.scala 39:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (!(2'h0 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
        if (!(2'h3 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
          tag_2 <= _GEN_1000;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 39:26]
      tag_3 <= 52'h0; // @[playground/src/noop/tlb.scala 39:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (!(2'h0 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
        if (!(2'h3 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
          tag_3 <= _GEN_1001;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 39:26]
      tag_4 <= 52'h0; // @[playground/src/noop/tlb.scala 39:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (!(2'h0 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
        if (!(2'h3 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
          tag_4 <= _GEN_1002;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 39:26]
      tag_5 <= 52'h0; // @[playground/src/noop/tlb.scala 39:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (!(2'h0 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
        if (!(2'h3 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
          tag_5 <= _GEN_1003;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 39:26]
      tag_6 <= 52'h0; // @[playground/src/noop/tlb.scala 39:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (!(2'h0 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
        if (!(2'h3 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
          tag_6 <= _GEN_1004;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 39:26]
      tag_7 <= 52'h0; // @[playground/src/noop/tlb.scala 39:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (!(2'h0 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
        if (!(2'h3 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
          tag_7 <= _GEN_1005;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 39:26]
      tag_8 <= 52'h0; // @[playground/src/noop/tlb.scala 39:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (!(2'h0 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
        if (!(2'h3 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
          tag_8 <= _GEN_1006;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 39:26]
      tag_9 <= 52'h0; // @[playground/src/noop/tlb.scala 39:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (!(2'h0 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
        if (!(2'h3 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
          tag_9 <= _GEN_1007;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 39:26]
      tag_10 <= 52'h0; // @[playground/src/noop/tlb.scala 39:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (!(2'h0 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
        if (!(2'h3 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
          tag_10 <= _GEN_1008;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 39:26]
      tag_11 <= 52'h0; // @[playground/src/noop/tlb.scala 39:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (!(2'h0 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
        if (!(2'h3 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
          tag_11 <= _GEN_1009;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 39:26]
      tag_12 <= 52'h0; // @[playground/src/noop/tlb.scala 39:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (!(2'h0 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
        if (!(2'h3 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
          tag_12 <= _GEN_1010;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 39:26]
      tag_13 <= 52'h0; // @[playground/src/noop/tlb.scala 39:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (!(2'h0 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
        if (!(2'h3 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
          tag_13 <= _GEN_1011;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 39:26]
      tag_14 <= 52'h0; // @[playground/src/noop/tlb.scala 39:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (!(2'h0 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
        if (!(2'h3 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
          tag_14 <= _GEN_1012;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 39:26]
      tag_15 <= 52'h0; // @[playground/src/noop/tlb.scala 39:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (!(2'h0 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
        if (!(2'h3 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
          tag_15 <= _GEN_1013;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 40:26]
      paddr_0 <= 20'h0; // @[playground/src/noop/tlb.scala 40:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (!(2'h0 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
        if (!(2'h3 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
          paddr_0 <= _GEN_1030;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 40:26]
      paddr_1 <= 20'h0; // @[playground/src/noop/tlb.scala 40:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (!(2'h0 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
        if (!(2'h3 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
          paddr_1 <= _GEN_1031;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 40:26]
      paddr_2 <= 20'h0; // @[playground/src/noop/tlb.scala 40:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (!(2'h0 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
        if (!(2'h3 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
          paddr_2 <= _GEN_1032;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 40:26]
      paddr_3 <= 20'h0; // @[playground/src/noop/tlb.scala 40:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (!(2'h0 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
        if (!(2'h3 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
          paddr_3 <= _GEN_1033;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 40:26]
      paddr_4 <= 20'h0; // @[playground/src/noop/tlb.scala 40:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (!(2'h0 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
        if (!(2'h3 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
          paddr_4 <= _GEN_1034;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 40:26]
      paddr_5 <= 20'h0; // @[playground/src/noop/tlb.scala 40:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (!(2'h0 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
        if (!(2'h3 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
          paddr_5 <= _GEN_1035;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 40:26]
      paddr_6 <= 20'h0; // @[playground/src/noop/tlb.scala 40:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (!(2'h0 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
        if (!(2'h3 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
          paddr_6 <= _GEN_1036;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 40:26]
      paddr_7 <= 20'h0; // @[playground/src/noop/tlb.scala 40:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (!(2'h0 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
        if (!(2'h3 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
          paddr_7 <= _GEN_1037;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 40:26]
      paddr_8 <= 20'h0; // @[playground/src/noop/tlb.scala 40:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (!(2'h0 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
        if (!(2'h3 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
          paddr_8 <= _GEN_1038;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 40:26]
      paddr_9 <= 20'h0; // @[playground/src/noop/tlb.scala 40:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (!(2'h0 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
        if (!(2'h3 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
          paddr_9 <= _GEN_1039;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 40:26]
      paddr_10 <= 20'h0; // @[playground/src/noop/tlb.scala 40:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (!(2'h0 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
        if (!(2'h3 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
          paddr_10 <= _GEN_1040;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 40:26]
      paddr_11 <= 20'h0; // @[playground/src/noop/tlb.scala 40:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (!(2'h0 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
        if (!(2'h3 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
          paddr_11 <= _GEN_1041;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 40:26]
      paddr_12 <= 20'h0; // @[playground/src/noop/tlb.scala 40:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (!(2'h0 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
        if (!(2'h3 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
          paddr_12 <= _GEN_1042;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 40:26]
      paddr_13 <= 20'h0; // @[playground/src/noop/tlb.scala 40:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (!(2'h0 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
        if (!(2'h3 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
          paddr_13 <= _GEN_1043;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 40:26]
      paddr_14 <= 20'h0; // @[playground/src/noop/tlb.scala 40:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (!(2'h0 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
        if (!(2'h3 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
          paddr_14 <= _GEN_1044;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 40:26]
      paddr_15 <= 20'h0; // @[playground/src/noop/tlb.scala 40:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (!(2'h0 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
        if (!(2'h3 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
          paddr_15 <= _GEN_1045;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 41:26]
      info_0 <= 10'h0; // @[playground/src/noop/tlb.scala 41:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (2'h0 == state) begin // @[playground/src/noop/tlb.scala 136:22]
        if (!(~handshake)) begin // @[playground/src/noop/tlb.scala 139:33]
          info_0 <= _GEN_243;
        end
      end else if (!(2'h3 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
        info_0 <= _GEN_1078;
      end
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 41:26]
      info_1 <= 10'h0; // @[playground/src/noop/tlb.scala 41:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (2'h0 == state) begin // @[playground/src/noop/tlb.scala 136:22]
        if (!(~handshake)) begin // @[playground/src/noop/tlb.scala 139:33]
          info_1 <= _GEN_244;
        end
      end else if (!(2'h3 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
        info_1 <= _GEN_1079;
      end
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 41:26]
      info_2 <= 10'h0; // @[playground/src/noop/tlb.scala 41:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (2'h0 == state) begin // @[playground/src/noop/tlb.scala 136:22]
        if (!(~handshake)) begin // @[playground/src/noop/tlb.scala 139:33]
          info_2 <= _GEN_245;
        end
      end else if (!(2'h3 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
        info_2 <= _GEN_1080;
      end
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 41:26]
      info_3 <= 10'h0; // @[playground/src/noop/tlb.scala 41:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (2'h0 == state) begin // @[playground/src/noop/tlb.scala 136:22]
        if (!(~handshake)) begin // @[playground/src/noop/tlb.scala 139:33]
          info_3 <= _GEN_246;
        end
      end else if (!(2'h3 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
        info_3 <= _GEN_1081;
      end
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 41:26]
      info_4 <= 10'h0; // @[playground/src/noop/tlb.scala 41:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (2'h0 == state) begin // @[playground/src/noop/tlb.scala 136:22]
        if (!(~handshake)) begin // @[playground/src/noop/tlb.scala 139:33]
          info_4 <= _GEN_247;
        end
      end else if (!(2'h3 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
        info_4 <= _GEN_1082;
      end
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 41:26]
      info_5 <= 10'h0; // @[playground/src/noop/tlb.scala 41:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (2'h0 == state) begin // @[playground/src/noop/tlb.scala 136:22]
        if (!(~handshake)) begin // @[playground/src/noop/tlb.scala 139:33]
          info_5 <= _GEN_248;
        end
      end else if (!(2'h3 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
        info_5 <= _GEN_1083;
      end
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 41:26]
      info_6 <= 10'h0; // @[playground/src/noop/tlb.scala 41:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (2'h0 == state) begin // @[playground/src/noop/tlb.scala 136:22]
        if (!(~handshake)) begin // @[playground/src/noop/tlb.scala 139:33]
          info_6 <= _GEN_249;
        end
      end else if (!(2'h3 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
        info_6 <= _GEN_1084;
      end
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 41:26]
      info_7 <= 10'h0; // @[playground/src/noop/tlb.scala 41:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (2'h0 == state) begin // @[playground/src/noop/tlb.scala 136:22]
        if (!(~handshake)) begin // @[playground/src/noop/tlb.scala 139:33]
          info_7 <= _GEN_250;
        end
      end else if (!(2'h3 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
        info_7 <= _GEN_1085;
      end
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 41:26]
      info_8 <= 10'h0; // @[playground/src/noop/tlb.scala 41:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (2'h0 == state) begin // @[playground/src/noop/tlb.scala 136:22]
        if (!(~handshake)) begin // @[playground/src/noop/tlb.scala 139:33]
          info_8 <= _GEN_251;
        end
      end else if (!(2'h3 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
        info_8 <= _GEN_1086;
      end
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 41:26]
      info_9 <= 10'h0; // @[playground/src/noop/tlb.scala 41:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (2'h0 == state) begin // @[playground/src/noop/tlb.scala 136:22]
        if (!(~handshake)) begin // @[playground/src/noop/tlb.scala 139:33]
          info_9 <= _GEN_252;
        end
      end else if (!(2'h3 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
        info_9 <= _GEN_1087;
      end
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 41:26]
      info_10 <= 10'h0; // @[playground/src/noop/tlb.scala 41:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (2'h0 == state) begin // @[playground/src/noop/tlb.scala 136:22]
        if (!(~handshake)) begin // @[playground/src/noop/tlb.scala 139:33]
          info_10 <= _GEN_253;
        end
      end else if (!(2'h3 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
        info_10 <= _GEN_1088;
      end
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 41:26]
      info_11 <= 10'h0; // @[playground/src/noop/tlb.scala 41:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (2'h0 == state) begin // @[playground/src/noop/tlb.scala 136:22]
        if (!(~handshake)) begin // @[playground/src/noop/tlb.scala 139:33]
          info_11 <= _GEN_254;
        end
      end else if (!(2'h3 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
        info_11 <= _GEN_1089;
      end
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 41:26]
      info_12 <= 10'h0; // @[playground/src/noop/tlb.scala 41:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (2'h0 == state) begin // @[playground/src/noop/tlb.scala 136:22]
        if (!(~handshake)) begin // @[playground/src/noop/tlb.scala 139:33]
          info_12 <= _GEN_255;
        end
      end else if (!(2'h3 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
        info_12 <= _GEN_1090;
      end
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 41:26]
      info_13 <= 10'h0; // @[playground/src/noop/tlb.scala 41:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (2'h0 == state) begin // @[playground/src/noop/tlb.scala 136:22]
        if (!(~handshake)) begin // @[playground/src/noop/tlb.scala 139:33]
          info_13 <= _GEN_256;
        end
      end else if (!(2'h3 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
        info_13 <= _GEN_1091;
      end
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 41:26]
      info_14 <= 10'h0; // @[playground/src/noop/tlb.scala 41:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (2'h0 == state) begin // @[playground/src/noop/tlb.scala 136:22]
        if (!(~handshake)) begin // @[playground/src/noop/tlb.scala 139:33]
          info_14 <= _GEN_257;
        end
      end else if (!(2'h3 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
        info_14 <= _GEN_1092;
      end
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 41:26]
      info_15 <= 10'h0; // @[playground/src/noop/tlb.scala 41:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (2'h0 == state) begin // @[playground/src/noop/tlb.scala 136:22]
        if (!(~handshake)) begin // @[playground/src/noop/tlb.scala 139:33]
          info_15 <= _GEN_258;
        end
      end else if (!(2'h3 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
        info_15 <= _GEN_1093;
      end
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 42:30]
      pte_addr_0 <= 32'h0; // @[playground/src/noop/tlb.scala 42:30]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (!(2'h0 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
        if (!(2'h3 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
          pte_addr_0 <= _GEN_1046;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 42:30]
      pte_addr_1 <= 32'h0; // @[playground/src/noop/tlb.scala 42:30]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (!(2'h0 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
        if (!(2'h3 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
          pte_addr_1 <= _GEN_1047;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 42:30]
      pte_addr_2 <= 32'h0; // @[playground/src/noop/tlb.scala 42:30]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (!(2'h0 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
        if (!(2'h3 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
          pte_addr_2 <= _GEN_1048;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 42:30]
      pte_addr_3 <= 32'h0; // @[playground/src/noop/tlb.scala 42:30]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (!(2'h0 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
        if (!(2'h3 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
          pte_addr_3 <= _GEN_1049;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 42:30]
      pte_addr_4 <= 32'h0; // @[playground/src/noop/tlb.scala 42:30]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (!(2'h0 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
        if (!(2'h3 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
          pte_addr_4 <= _GEN_1050;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 42:30]
      pte_addr_5 <= 32'h0; // @[playground/src/noop/tlb.scala 42:30]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (!(2'h0 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
        if (!(2'h3 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
          pte_addr_5 <= _GEN_1051;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 42:30]
      pte_addr_6 <= 32'h0; // @[playground/src/noop/tlb.scala 42:30]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (!(2'h0 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
        if (!(2'h3 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
          pte_addr_6 <= _GEN_1052;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 42:30]
      pte_addr_7 <= 32'h0; // @[playground/src/noop/tlb.scala 42:30]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (!(2'h0 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
        if (!(2'h3 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
          pte_addr_7 <= _GEN_1053;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 42:30]
      pte_addr_8 <= 32'h0; // @[playground/src/noop/tlb.scala 42:30]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (!(2'h0 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
        if (!(2'h3 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
          pte_addr_8 <= _GEN_1054;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 42:30]
      pte_addr_9 <= 32'h0; // @[playground/src/noop/tlb.scala 42:30]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (!(2'h0 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
        if (!(2'h3 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
          pte_addr_9 <= _GEN_1055;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 42:30]
      pte_addr_10 <= 32'h0; // @[playground/src/noop/tlb.scala 42:30]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (!(2'h0 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
        if (!(2'h3 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
          pte_addr_10 <= _GEN_1056;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 42:30]
      pte_addr_11 <= 32'h0; // @[playground/src/noop/tlb.scala 42:30]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (!(2'h0 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
        if (!(2'h3 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
          pte_addr_11 <= _GEN_1057;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 42:30]
      pte_addr_12 <= 32'h0; // @[playground/src/noop/tlb.scala 42:30]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (!(2'h0 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
        if (!(2'h3 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
          pte_addr_12 <= _GEN_1058;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 42:30]
      pte_addr_13 <= 32'h0; // @[playground/src/noop/tlb.scala 42:30]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (!(2'h0 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
        if (!(2'h3 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
          pte_addr_13 <= _GEN_1059;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 42:30]
      pte_addr_14 <= 32'h0; // @[playground/src/noop/tlb.scala 42:30]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (!(2'h0 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
        if (!(2'h3 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
          pte_addr_14 <= _GEN_1060;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 42:30]
      pte_addr_15 <= 32'h0; // @[playground/src/noop/tlb.scala 42:30]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (!(2'h0 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
        if (!(2'h3 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
          pte_addr_15 <= _GEN_1061;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 43:30]
      pte_level_0 <= 2'h0; // @[playground/src/noop/tlb.scala 43:30]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (!(2'h0 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
        if (!(2'h3 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
          pte_level_0 <= _GEN_1062;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 43:30]
      pte_level_1 <= 2'h0; // @[playground/src/noop/tlb.scala 43:30]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (!(2'h0 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
        if (!(2'h3 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
          pte_level_1 <= _GEN_1063;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 43:30]
      pte_level_2 <= 2'h0; // @[playground/src/noop/tlb.scala 43:30]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (!(2'h0 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
        if (!(2'h3 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
          pte_level_2 <= _GEN_1064;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 43:30]
      pte_level_3 <= 2'h0; // @[playground/src/noop/tlb.scala 43:30]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (!(2'h0 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
        if (!(2'h3 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
          pte_level_3 <= _GEN_1065;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 43:30]
      pte_level_4 <= 2'h0; // @[playground/src/noop/tlb.scala 43:30]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (!(2'h0 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
        if (!(2'h3 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
          pte_level_4 <= _GEN_1066;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 43:30]
      pte_level_5 <= 2'h0; // @[playground/src/noop/tlb.scala 43:30]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (!(2'h0 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
        if (!(2'h3 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
          pte_level_5 <= _GEN_1067;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 43:30]
      pte_level_6 <= 2'h0; // @[playground/src/noop/tlb.scala 43:30]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (!(2'h0 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
        if (!(2'h3 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
          pte_level_6 <= _GEN_1068;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 43:30]
      pte_level_7 <= 2'h0; // @[playground/src/noop/tlb.scala 43:30]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (!(2'h0 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
        if (!(2'h3 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
          pte_level_7 <= _GEN_1069;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 43:30]
      pte_level_8 <= 2'h0; // @[playground/src/noop/tlb.scala 43:30]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (!(2'h0 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
        if (!(2'h3 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
          pte_level_8 <= _GEN_1070;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 43:30]
      pte_level_9 <= 2'h0; // @[playground/src/noop/tlb.scala 43:30]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (!(2'h0 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
        if (!(2'h3 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
          pte_level_9 <= _GEN_1071;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 43:30]
      pte_level_10 <= 2'h0; // @[playground/src/noop/tlb.scala 43:30]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (!(2'h0 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
        if (!(2'h3 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
          pte_level_10 <= _GEN_1072;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 43:30]
      pte_level_11 <= 2'h0; // @[playground/src/noop/tlb.scala 43:30]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (!(2'h0 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
        if (!(2'h3 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
          pte_level_11 <= _GEN_1073;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 43:30]
      pte_level_12 <= 2'h0; // @[playground/src/noop/tlb.scala 43:30]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (!(2'h0 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
        if (!(2'h3 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
          pte_level_12 <= _GEN_1074;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 43:30]
      pte_level_13 <= 2'h0; // @[playground/src/noop/tlb.scala 43:30]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (!(2'h0 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
        if (!(2'h3 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
          pte_level_13 <= _GEN_1075;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 43:30]
      pte_level_14 <= 2'h0; // @[playground/src/noop/tlb.scala 43:30]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (!(2'h0 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
        if (!(2'h3 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
          pte_level_14 <= _GEN_1076;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 43:30]
      pte_level_15 <= 2'h0; // @[playground/src/noop/tlb.scala 43:30]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (!(2'h0 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
        if (!(2'h3 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
          pte_level_15 <= _GEN_1077;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 44:26]
      valid_0 <= 1'h0; // @[playground/src/noop/tlb.scala 44:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (2'h0 == state) begin // @[playground/src/noop/tlb.scala 136:22]
        valid_0 <= _GEN_130;
      end else if (2'h3 == state) begin // @[playground/src/noop/tlb.scala 136:22]
        valid_0 <= _GEN_130;
      end else begin
        valid_0 <= _GEN_1014;
      end
    end else begin
      valid_0 <= _GEN_130;
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 44:26]
      valid_1 <= 1'h0; // @[playground/src/noop/tlb.scala 44:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (2'h0 == state) begin // @[playground/src/noop/tlb.scala 136:22]
        valid_1 <= _GEN_131;
      end else if (2'h3 == state) begin // @[playground/src/noop/tlb.scala 136:22]
        valid_1 <= _GEN_131;
      end else begin
        valid_1 <= _GEN_1015;
      end
    end else begin
      valid_1 <= _GEN_131;
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 44:26]
      valid_2 <= 1'h0; // @[playground/src/noop/tlb.scala 44:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (2'h0 == state) begin // @[playground/src/noop/tlb.scala 136:22]
        valid_2 <= _GEN_132;
      end else if (2'h3 == state) begin // @[playground/src/noop/tlb.scala 136:22]
        valid_2 <= _GEN_132;
      end else begin
        valid_2 <= _GEN_1016;
      end
    end else begin
      valid_2 <= _GEN_132;
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 44:26]
      valid_3 <= 1'h0; // @[playground/src/noop/tlb.scala 44:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (2'h0 == state) begin // @[playground/src/noop/tlb.scala 136:22]
        valid_3 <= _GEN_133;
      end else if (2'h3 == state) begin // @[playground/src/noop/tlb.scala 136:22]
        valid_3 <= _GEN_133;
      end else begin
        valid_3 <= _GEN_1017;
      end
    end else begin
      valid_3 <= _GEN_133;
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 44:26]
      valid_4 <= 1'h0; // @[playground/src/noop/tlb.scala 44:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (2'h0 == state) begin // @[playground/src/noop/tlb.scala 136:22]
        valid_4 <= _GEN_134;
      end else if (2'h3 == state) begin // @[playground/src/noop/tlb.scala 136:22]
        valid_4 <= _GEN_134;
      end else begin
        valid_4 <= _GEN_1018;
      end
    end else begin
      valid_4 <= _GEN_134;
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 44:26]
      valid_5 <= 1'h0; // @[playground/src/noop/tlb.scala 44:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (2'h0 == state) begin // @[playground/src/noop/tlb.scala 136:22]
        valid_5 <= _GEN_135;
      end else if (2'h3 == state) begin // @[playground/src/noop/tlb.scala 136:22]
        valid_5 <= _GEN_135;
      end else begin
        valid_5 <= _GEN_1019;
      end
    end else begin
      valid_5 <= _GEN_135;
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 44:26]
      valid_6 <= 1'h0; // @[playground/src/noop/tlb.scala 44:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (2'h0 == state) begin // @[playground/src/noop/tlb.scala 136:22]
        valid_6 <= _GEN_136;
      end else if (2'h3 == state) begin // @[playground/src/noop/tlb.scala 136:22]
        valid_6 <= _GEN_136;
      end else begin
        valid_6 <= _GEN_1020;
      end
    end else begin
      valid_6 <= _GEN_136;
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 44:26]
      valid_7 <= 1'h0; // @[playground/src/noop/tlb.scala 44:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (2'h0 == state) begin // @[playground/src/noop/tlb.scala 136:22]
        valid_7 <= _GEN_137;
      end else if (2'h3 == state) begin // @[playground/src/noop/tlb.scala 136:22]
        valid_7 <= _GEN_137;
      end else begin
        valid_7 <= _GEN_1021;
      end
    end else begin
      valid_7 <= _GEN_137;
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 44:26]
      valid_8 <= 1'h0; // @[playground/src/noop/tlb.scala 44:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (2'h0 == state) begin // @[playground/src/noop/tlb.scala 136:22]
        valid_8 <= _GEN_138;
      end else if (2'h3 == state) begin // @[playground/src/noop/tlb.scala 136:22]
        valid_8 <= _GEN_138;
      end else begin
        valid_8 <= _GEN_1022;
      end
    end else begin
      valid_8 <= _GEN_138;
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 44:26]
      valid_9 <= 1'h0; // @[playground/src/noop/tlb.scala 44:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (2'h0 == state) begin // @[playground/src/noop/tlb.scala 136:22]
        valid_9 <= _GEN_139;
      end else if (2'h3 == state) begin // @[playground/src/noop/tlb.scala 136:22]
        valid_9 <= _GEN_139;
      end else begin
        valid_9 <= _GEN_1023;
      end
    end else begin
      valid_9 <= _GEN_139;
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 44:26]
      valid_10 <= 1'h0; // @[playground/src/noop/tlb.scala 44:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (2'h0 == state) begin // @[playground/src/noop/tlb.scala 136:22]
        valid_10 <= _GEN_140;
      end else if (2'h3 == state) begin // @[playground/src/noop/tlb.scala 136:22]
        valid_10 <= _GEN_140;
      end else begin
        valid_10 <= _GEN_1024;
      end
    end else begin
      valid_10 <= _GEN_140;
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 44:26]
      valid_11 <= 1'h0; // @[playground/src/noop/tlb.scala 44:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (2'h0 == state) begin // @[playground/src/noop/tlb.scala 136:22]
        valid_11 <= _GEN_141;
      end else if (2'h3 == state) begin // @[playground/src/noop/tlb.scala 136:22]
        valid_11 <= _GEN_141;
      end else begin
        valid_11 <= _GEN_1025;
      end
    end else begin
      valid_11 <= _GEN_141;
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 44:26]
      valid_12 <= 1'h0; // @[playground/src/noop/tlb.scala 44:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (2'h0 == state) begin // @[playground/src/noop/tlb.scala 136:22]
        valid_12 <= _GEN_142;
      end else if (2'h3 == state) begin // @[playground/src/noop/tlb.scala 136:22]
        valid_12 <= _GEN_142;
      end else begin
        valid_12 <= _GEN_1026;
      end
    end else begin
      valid_12 <= _GEN_142;
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 44:26]
      valid_13 <= 1'h0; // @[playground/src/noop/tlb.scala 44:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (2'h0 == state) begin // @[playground/src/noop/tlb.scala 136:22]
        valid_13 <= _GEN_143;
      end else if (2'h3 == state) begin // @[playground/src/noop/tlb.scala 136:22]
        valid_13 <= _GEN_143;
      end else begin
        valid_13 <= _GEN_1027;
      end
    end else begin
      valid_13 <= _GEN_143;
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 44:26]
      valid_14 <= 1'h0; // @[playground/src/noop/tlb.scala 44:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (2'h0 == state) begin // @[playground/src/noop/tlb.scala 136:22]
        valid_14 <= _GEN_144;
      end else if (2'h3 == state) begin // @[playground/src/noop/tlb.scala 136:22]
        valid_14 <= _GEN_144;
      end else begin
        valid_14 <= _GEN_1028;
      end
    end else begin
      valid_14 <= _GEN_144;
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 44:26]
      valid_15 <= 1'h0; // @[playground/src/noop/tlb.scala 44:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (2'h0 == state) begin // @[playground/src/noop/tlb.scala 136:22]
        valid_15 <= _GEN_145;
      end else if (2'h3 == state) begin // @[playground/src/noop/tlb.scala 136:22]
        valid_15 <= _GEN_145;
      end else begin
        valid_15 <= _GEN_1029;
      end
    end else begin
      valid_15 <= _GEN_145;
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 46:30]
      pre_addr <= 64'h0; // @[playground/src/noop/tlb.scala 46:30]
    end else if (handshake) begin // @[playground/src/noop/tlb.scala 101:20]
      pre_addr <= io_va2pa_vaddr; // @[playground/src/noop/tlb.scala 103:18]
    end else if (io_va2pa_ready & io_va2pa_vvalid) begin // @[playground/src/noop/tlb.scala 54:44]
      pre_addr <= io_va2pa_vaddr; // @[playground/src/noop/tlb.scala 55:18]
    end
    pte_addr_r <= _GEN_1418[31:0]; // @[playground/src/noop/tlb.scala 47:{30,30}]
    if (reset) begin // @[playground/src/noop/tlb.scala 48:30]
      wpte_data_r <= 64'h0; // @[playground/src/noop/tlb.scala 48:30]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (2'h0 == state) begin // @[playground/src/noop/tlb.scala 136:22]
        if (!(~handshake)) begin // @[playground/src/noop/tlb.scala 139:33]
          wpte_data_r <= _GEN_242;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 49:30]
      dc_mode_r <= 5'h0; // @[playground/src/noop/tlb.scala 49:30]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (2'h0 == state) begin // @[playground/src/noop/tlb.scala 136:22]
        if (~handshake) begin // @[playground/src/noop/tlb.scala 139:33]
          dc_mode_r <= 5'h0; // @[playground/src/noop/tlb.scala 138:27]
        end else begin
          dc_mode_r <= _GEN_261;
        end
      end else if (2'h3 == state) begin // @[playground/src/noop/tlb.scala 136:22]
        dc_mode_r <= _GEN_294;
      end else begin
        dc_mode_r <= _GEN_992;
      end
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 51:30]
      out_valid_r <= 1'h0; // @[playground/src/noop/tlb.scala 51:30]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (2'h0 == state) begin // @[playground/src/noop/tlb.scala 136:22]
        if (~handshake) begin // @[playground/src/noop/tlb.scala 139:33]
          out_valid_r <= _GEN_150;
        end else begin
          out_valid_r <= _GEN_237;
        end
      end else begin
        out_valid_r <= _GEN_150;
      end
    end else begin
      out_valid_r <= io_va2pa_vvalid; // @[playground/src/noop/tlb.scala 232:21]
    end
    out_paddr_r <= _GEN_1419[31:0]; // @[playground/src/noop/tlb.scala 52:{30,30}]
    if (reset) begin // @[playground/src/noop/tlb.scala 53:30]
      out_excep_r_cause <= 64'h0; // @[playground/src/noop/tlb.scala 53:30]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (2'h0 == state) begin // @[playground/src/noop/tlb.scala 136:22]
        if (!(~handshake)) begin // @[playground/src/noop/tlb.scala 139:33]
          out_excep_r_cause <= _GEN_235;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 53:30]
      out_excep_r_tval <= 64'h0; // @[playground/src/noop/tlb.scala 53:30]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (2'h0 == state) begin // @[playground/src/noop/tlb.scala 136:22]
        if (!(~handshake)) begin // @[playground/src/noop/tlb.scala 139:33]
          out_excep_r_tval <= _GEN_236;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 53:30]
      out_excep_r_en <= 1'h0; // @[playground/src/noop/tlb.scala 53:30]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (2'h0 == state) begin // @[playground/src/noop/tlb.scala 136:22]
        if (~handshake) begin // @[playground/src/noop/tlb.scala 139:33]
          out_excep_r_en <= _GEN_151;
        end else begin
          out_excep_r_en <= _GEN_234;
        end
      end else if (2'h3 == state) begin // @[playground/src/noop/tlb.scala 136:22]
        out_excep_r_en <= _GEN_151;
      end else begin
        out_excep_r_en <= _GEN_996;
      end
    end else begin
      out_excep_r_en <= _GEN_151;
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 84:24]
      state <= 2'h0; // @[playground/src/noop/tlb.scala 84:24]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (2'h0 == state) begin // @[playground/src/noop/tlb.scala 136:22]
        if (!(~handshake)) begin // @[playground/src/noop/tlb.scala 139:33]
          state <= _GEN_239;
        end
      end else if (2'h3 == state) begin // @[playground/src/noop/tlb.scala 136:22]
        state <= _GEN_296;
      end else begin
        state <= _GEN_995;
      end
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 85:26]
      flush_r <= 1'h0; // @[playground/src/noop/tlb.scala 85:26]
    end else if (io_flush | flush_r) begin // @[playground/src/noop/tlb.scala 86:30]
      if (state == 2'h0) begin // @[playground/src/noop/tlb.scala 87:30]
        flush_r <= 1'h0; // @[playground/src/noop/tlb.scala 89:21]
      end else begin
        flush_r <= 1'h1; // @[playground/src/noop/tlb.scala 91:21]
      end
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 95:27]
      m_type_r <= 2'h0; // @[playground/src/noop/tlb.scala 95:27]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (2'h0 == state) begin // @[playground/src/noop/tlb.scala 136:22]
        if (!(~handshake)) begin // @[playground/src/noop/tlb.scala 139:33]
          m_type_r <= _GEN_260;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 130:27]
      select_r <= 4'h0; // @[playground/src/noop/tlb.scala 130:27]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (2'h0 == state) begin // @[playground/src/noop/tlb.scala 136:22]
        if (!(~handshake)) begin // @[playground/src/noop/tlb.scala 139:33]
          select_r <= _GEN_259;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 131:26]
      offset <= 8'h0; // @[playground/src/noop/tlb.scala 131:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (2'h0 == state) begin // @[playground/src/noop/tlb.scala 136:22]
        if (!(~handshake)) begin // @[playground/src/noop/tlb.scala 139:33]
          offset <= _GEN_262;
        end
      end else if (!(2'h3 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
        offset <= _GEN_993;
      end
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 132:26]
      level <= 2'h0; // @[playground/src/noop/tlb.scala 132:26]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (2'h0 == state) begin // @[playground/src/noop/tlb.scala 136:22]
        if (!(~handshake)) begin // @[playground/src/noop/tlb.scala 139:33]
          level <= _GEN_263;
        end
      end else if (!(2'h3 == state)) begin // @[playground/src/noop/tlb.scala 136:22]
        level <= _GEN_994;
      end
    end
    if (reset) begin // @[playground/src/noop/tlb.scala 134:28]
      wpte_hs_r <= 1'h0; // @[playground/src/noop/tlb.scala 134:28]
    end else if (is_Sv39 | state != 2'h0) begin // @[playground/src/noop/tlb.scala 135:37]
      if (2'h0 == state) begin // @[playground/src/noop/tlb.scala 136:22]
        if (!(~handshake)) begin // @[playground/src/noop/tlb.scala 139:33]
          wpte_hs_r <= _GEN_240;
        end
      end else if (2'h3 == state) begin // @[playground/src/noop/tlb.scala 136:22]
        wpte_hs_r <= _GEN_295;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  tag_0 = _RAND_0[51:0];
  _RAND_1 = {2{`RANDOM}};
  tag_1 = _RAND_1[51:0];
  _RAND_2 = {2{`RANDOM}};
  tag_2 = _RAND_2[51:0];
  _RAND_3 = {2{`RANDOM}};
  tag_3 = _RAND_3[51:0];
  _RAND_4 = {2{`RANDOM}};
  tag_4 = _RAND_4[51:0];
  _RAND_5 = {2{`RANDOM}};
  tag_5 = _RAND_5[51:0];
  _RAND_6 = {2{`RANDOM}};
  tag_6 = _RAND_6[51:0];
  _RAND_7 = {2{`RANDOM}};
  tag_7 = _RAND_7[51:0];
  _RAND_8 = {2{`RANDOM}};
  tag_8 = _RAND_8[51:0];
  _RAND_9 = {2{`RANDOM}};
  tag_9 = _RAND_9[51:0];
  _RAND_10 = {2{`RANDOM}};
  tag_10 = _RAND_10[51:0];
  _RAND_11 = {2{`RANDOM}};
  tag_11 = _RAND_11[51:0];
  _RAND_12 = {2{`RANDOM}};
  tag_12 = _RAND_12[51:0];
  _RAND_13 = {2{`RANDOM}};
  tag_13 = _RAND_13[51:0];
  _RAND_14 = {2{`RANDOM}};
  tag_14 = _RAND_14[51:0];
  _RAND_15 = {2{`RANDOM}};
  tag_15 = _RAND_15[51:0];
  _RAND_16 = {1{`RANDOM}};
  paddr_0 = _RAND_16[19:0];
  _RAND_17 = {1{`RANDOM}};
  paddr_1 = _RAND_17[19:0];
  _RAND_18 = {1{`RANDOM}};
  paddr_2 = _RAND_18[19:0];
  _RAND_19 = {1{`RANDOM}};
  paddr_3 = _RAND_19[19:0];
  _RAND_20 = {1{`RANDOM}};
  paddr_4 = _RAND_20[19:0];
  _RAND_21 = {1{`RANDOM}};
  paddr_5 = _RAND_21[19:0];
  _RAND_22 = {1{`RANDOM}};
  paddr_6 = _RAND_22[19:0];
  _RAND_23 = {1{`RANDOM}};
  paddr_7 = _RAND_23[19:0];
  _RAND_24 = {1{`RANDOM}};
  paddr_8 = _RAND_24[19:0];
  _RAND_25 = {1{`RANDOM}};
  paddr_9 = _RAND_25[19:0];
  _RAND_26 = {1{`RANDOM}};
  paddr_10 = _RAND_26[19:0];
  _RAND_27 = {1{`RANDOM}};
  paddr_11 = _RAND_27[19:0];
  _RAND_28 = {1{`RANDOM}};
  paddr_12 = _RAND_28[19:0];
  _RAND_29 = {1{`RANDOM}};
  paddr_13 = _RAND_29[19:0];
  _RAND_30 = {1{`RANDOM}};
  paddr_14 = _RAND_30[19:0];
  _RAND_31 = {1{`RANDOM}};
  paddr_15 = _RAND_31[19:0];
  _RAND_32 = {1{`RANDOM}};
  info_0 = _RAND_32[9:0];
  _RAND_33 = {1{`RANDOM}};
  info_1 = _RAND_33[9:0];
  _RAND_34 = {1{`RANDOM}};
  info_2 = _RAND_34[9:0];
  _RAND_35 = {1{`RANDOM}};
  info_3 = _RAND_35[9:0];
  _RAND_36 = {1{`RANDOM}};
  info_4 = _RAND_36[9:0];
  _RAND_37 = {1{`RANDOM}};
  info_5 = _RAND_37[9:0];
  _RAND_38 = {1{`RANDOM}};
  info_6 = _RAND_38[9:0];
  _RAND_39 = {1{`RANDOM}};
  info_7 = _RAND_39[9:0];
  _RAND_40 = {1{`RANDOM}};
  info_8 = _RAND_40[9:0];
  _RAND_41 = {1{`RANDOM}};
  info_9 = _RAND_41[9:0];
  _RAND_42 = {1{`RANDOM}};
  info_10 = _RAND_42[9:0];
  _RAND_43 = {1{`RANDOM}};
  info_11 = _RAND_43[9:0];
  _RAND_44 = {1{`RANDOM}};
  info_12 = _RAND_44[9:0];
  _RAND_45 = {1{`RANDOM}};
  info_13 = _RAND_45[9:0];
  _RAND_46 = {1{`RANDOM}};
  info_14 = _RAND_46[9:0];
  _RAND_47 = {1{`RANDOM}};
  info_15 = _RAND_47[9:0];
  _RAND_48 = {1{`RANDOM}};
  pte_addr_0 = _RAND_48[31:0];
  _RAND_49 = {1{`RANDOM}};
  pte_addr_1 = _RAND_49[31:0];
  _RAND_50 = {1{`RANDOM}};
  pte_addr_2 = _RAND_50[31:0];
  _RAND_51 = {1{`RANDOM}};
  pte_addr_3 = _RAND_51[31:0];
  _RAND_52 = {1{`RANDOM}};
  pte_addr_4 = _RAND_52[31:0];
  _RAND_53 = {1{`RANDOM}};
  pte_addr_5 = _RAND_53[31:0];
  _RAND_54 = {1{`RANDOM}};
  pte_addr_6 = _RAND_54[31:0];
  _RAND_55 = {1{`RANDOM}};
  pte_addr_7 = _RAND_55[31:0];
  _RAND_56 = {1{`RANDOM}};
  pte_addr_8 = _RAND_56[31:0];
  _RAND_57 = {1{`RANDOM}};
  pte_addr_9 = _RAND_57[31:0];
  _RAND_58 = {1{`RANDOM}};
  pte_addr_10 = _RAND_58[31:0];
  _RAND_59 = {1{`RANDOM}};
  pte_addr_11 = _RAND_59[31:0];
  _RAND_60 = {1{`RANDOM}};
  pte_addr_12 = _RAND_60[31:0];
  _RAND_61 = {1{`RANDOM}};
  pte_addr_13 = _RAND_61[31:0];
  _RAND_62 = {1{`RANDOM}};
  pte_addr_14 = _RAND_62[31:0];
  _RAND_63 = {1{`RANDOM}};
  pte_addr_15 = _RAND_63[31:0];
  _RAND_64 = {1{`RANDOM}};
  pte_level_0 = _RAND_64[1:0];
  _RAND_65 = {1{`RANDOM}};
  pte_level_1 = _RAND_65[1:0];
  _RAND_66 = {1{`RANDOM}};
  pte_level_2 = _RAND_66[1:0];
  _RAND_67 = {1{`RANDOM}};
  pte_level_3 = _RAND_67[1:0];
  _RAND_68 = {1{`RANDOM}};
  pte_level_4 = _RAND_68[1:0];
  _RAND_69 = {1{`RANDOM}};
  pte_level_5 = _RAND_69[1:0];
  _RAND_70 = {1{`RANDOM}};
  pte_level_6 = _RAND_70[1:0];
  _RAND_71 = {1{`RANDOM}};
  pte_level_7 = _RAND_71[1:0];
  _RAND_72 = {1{`RANDOM}};
  pte_level_8 = _RAND_72[1:0];
  _RAND_73 = {1{`RANDOM}};
  pte_level_9 = _RAND_73[1:0];
  _RAND_74 = {1{`RANDOM}};
  pte_level_10 = _RAND_74[1:0];
  _RAND_75 = {1{`RANDOM}};
  pte_level_11 = _RAND_75[1:0];
  _RAND_76 = {1{`RANDOM}};
  pte_level_12 = _RAND_76[1:0];
  _RAND_77 = {1{`RANDOM}};
  pte_level_13 = _RAND_77[1:0];
  _RAND_78 = {1{`RANDOM}};
  pte_level_14 = _RAND_78[1:0];
  _RAND_79 = {1{`RANDOM}};
  pte_level_15 = _RAND_79[1:0];
  _RAND_80 = {1{`RANDOM}};
  valid_0 = _RAND_80[0:0];
  _RAND_81 = {1{`RANDOM}};
  valid_1 = _RAND_81[0:0];
  _RAND_82 = {1{`RANDOM}};
  valid_2 = _RAND_82[0:0];
  _RAND_83 = {1{`RANDOM}};
  valid_3 = _RAND_83[0:0];
  _RAND_84 = {1{`RANDOM}};
  valid_4 = _RAND_84[0:0];
  _RAND_85 = {1{`RANDOM}};
  valid_5 = _RAND_85[0:0];
  _RAND_86 = {1{`RANDOM}};
  valid_6 = _RAND_86[0:0];
  _RAND_87 = {1{`RANDOM}};
  valid_7 = _RAND_87[0:0];
  _RAND_88 = {1{`RANDOM}};
  valid_8 = _RAND_88[0:0];
  _RAND_89 = {1{`RANDOM}};
  valid_9 = _RAND_89[0:0];
  _RAND_90 = {1{`RANDOM}};
  valid_10 = _RAND_90[0:0];
  _RAND_91 = {1{`RANDOM}};
  valid_11 = _RAND_91[0:0];
  _RAND_92 = {1{`RANDOM}};
  valid_12 = _RAND_92[0:0];
  _RAND_93 = {1{`RANDOM}};
  valid_13 = _RAND_93[0:0];
  _RAND_94 = {1{`RANDOM}};
  valid_14 = _RAND_94[0:0];
  _RAND_95 = {1{`RANDOM}};
  valid_15 = _RAND_95[0:0];
  _RAND_96 = {2{`RANDOM}};
  pre_addr = _RAND_96[63:0];
  _RAND_97 = {1{`RANDOM}};
  pte_addr_r = _RAND_97[31:0];
  _RAND_98 = {2{`RANDOM}};
  wpte_data_r = _RAND_98[63:0];
  _RAND_99 = {1{`RANDOM}};
  dc_mode_r = _RAND_99[4:0];
  _RAND_100 = {1{`RANDOM}};
  out_valid_r = _RAND_100[0:0];
  _RAND_101 = {1{`RANDOM}};
  out_paddr_r = _RAND_101[31:0];
  _RAND_102 = {2{`RANDOM}};
  out_excep_r_cause = _RAND_102[63:0];
  _RAND_103 = {2{`RANDOM}};
  out_excep_r_tval = _RAND_103[63:0];
  _RAND_104 = {1{`RANDOM}};
  out_excep_r_en = _RAND_104[0:0];
  _RAND_105 = {1{`RANDOM}};
  state = _RAND_105[1:0];
  _RAND_106 = {1{`RANDOM}};
  flush_r = _RAND_106[0:0];
  _RAND_107 = {1{`RANDOM}};
  m_type_r = _RAND_107[1:0];
  _RAND_108 = {1{`RANDOM}};
  select_r = _RAND_108[3:0];
  _RAND_109 = {1{`RANDOM}};
  offset = _RAND_109[7:0];
  _RAND_110 = {1{`RANDOM}};
  level = _RAND_110[1:0];
  _RAND_111 = {1{`RANDOM}};
  wpte_hs_r = _RAND_111[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module DcacheSelector(
  input         clock,
  input         reset,
  input  [31:0] io_tlb_if2dc_addr, // @[playground/src/noop/dcache.scala 15:16]
  output [63:0] io_tlb_if2dc_rdata, // @[playground/src/noop/dcache.scala 15:16]
  output        io_tlb_if2dc_rvalid, // @[playground/src/noop/dcache.scala 15:16]
  input  [63:0] io_tlb_if2dc_wdata, // @[playground/src/noop/dcache.scala 15:16]
  input  [4:0]  io_tlb_if2dc_dc_mode, // @[playground/src/noop/dcache.scala 15:16]
  output        io_tlb_if2dc_ready, // @[playground/src/noop/dcache.scala 15:16]
  input  [31:0] io_tlb_mem2dc_addr, // @[playground/src/noop/dcache.scala 15:16]
  output [63:0] io_tlb_mem2dc_rdata, // @[playground/src/noop/dcache.scala 15:16]
  output        io_tlb_mem2dc_rvalid, // @[playground/src/noop/dcache.scala 15:16]
  input  [63:0] io_tlb_mem2dc_wdata, // @[playground/src/noop/dcache.scala 15:16]
  input  [4:0]  io_tlb_mem2dc_dc_mode, // @[playground/src/noop/dcache.scala 15:16]
  output        io_tlb_mem2dc_ready, // @[playground/src/noop/dcache.scala 15:16]
  input  [31:0] io_mem2dc_addr, // @[playground/src/noop/dcache.scala 15:16]
  output [63:0] io_mem2dc_rdata, // @[playground/src/noop/dcache.scala 15:16]
  output        io_mem2dc_rvalid, // @[playground/src/noop/dcache.scala 15:16]
  input  [63:0] io_mem2dc_wdata, // @[playground/src/noop/dcache.scala 15:16]
  input  [4:0]  io_mem2dc_dc_mode, // @[playground/src/noop/dcache.scala 15:16]
  input  [4:0]  io_mem2dc_amo, // @[playground/src/noop/dcache.scala 15:16]
  output        io_mem2dc_ready, // @[playground/src/noop/dcache.scala 15:16]
  input  [31:0] io_dma2dc_addr, // @[playground/src/noop/dcache.scala 15:16]
  output [63:0] io_dma2dc_rdata, // @[playground/src/noop/dcache.scala 15:16]
  output        io_dma2dc_rvalid, // @[playground/src/noop/dcache.scala 15:16]
  input  [63:0] io_dma2dc_wdata, // @[playground/src/noop/dcache.scala 15:16]
  input  [4:0]  io_dma2dc_dc_mode, // @[playground/src/noop/dcache.scala 15:16]
  output        io_dma2dc_ready, // @[playground/src/noop/dcache.scala 15:16]
  output [31:0] io_select_addr, // @[playground/src/noop/dcache.scala 15:16]
  input  [63:0] io_select_rdata, // @[playground/src/noop/dcache.scala 15:16]
  input         io_select_rvalid, // @[playground/src/noop/dcache.scala 15:16]
  output [63:0] io_select_wdata, // @[playground/src/noop/dcache.scala 15:16]
  output [4:0]  io_select_dc_mode, // @[playground/src/noop/dcache.scala 15:16]
  output [4:0]  io_select_amo, // @[playground/src/noop/dcache.scala 15:16]
  input         io_select_ready // @[playground/src/noop/dcache.scala 15:16]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg [1:0] pre_idx; // @[playground/src/noop/dcache.scala 30:26]
  reg  busy; // @[playground/src/noop/dcache.scala 31:26]
  wire  _GEN_0 = io_select_rvalid ? 1'h0 : busy; // @[playground/src/noop/dcache.scala 37:27 38:14 31:26]
  wire [1:0] _GEN_1 = io_dma2dc_dc_mode != 5'h0 ? 2'h3 : pre_idx; // @[playground/src/noop/dcache.scala 65:47 66:17 30:26]
  wire  _GEN_2 = io_dma2dc_dc_mode != 5'h0 ? io_select_ready : _GEN_0; // @[playground/src/noop/dcache.scala 65:47 67:17]
  wire [31:0] _GEN_3 = io_dma2dc_dc_mode != 5'h0 ? io_dma2dc_addr : 32'h0; // @[playground/src/noop/dcache.scala 32:25 65:47 68:29]
  wire [63:0] _GEN_4 = io_dma2dc_dc_mode != 5'h0 ? io_dma2dc_wdata : 64'h0; // @[playground/src/noop/dcache.scala 33:25 65:47 69:29]
  wire [4:0] _GEN_5 = io_dma2dc_dc_mode != 5'h0 ? io_dma2dc_dc_mode : 5'h0; // @[playground/src/noop/dcache.scala 34:25 65:47 70:29]
  wire  _GEN_7 = io_dma2dc_dc_mode != 5'h0 & io_select_ready; // @[playground/src/noop/dcache.scala 65:47 72:29 29:69]
  wire [1:0] _GEN_8 = io_tlb_if2dc_dc_mode != 5'h0 ? 2'h2 : _GEN_1; // @[playground/src/noop/dcache.scala 57:50 58:17]
  wire  _GEN_9 = io_tlb_if2dc_dc_mode != 5'h0 ? io_select_ready : _GEN_2; // @[playground/src/noop/dcache.scala 57:50 59:17]
  wire [31:0] _GEN_10 = io_tlb_if2dc_dc_mode != 5'h0 ? io_tlb_if2dc_addr : _GEN_3; // @[playground/src/noop/dcache.scala 57:50 60:29]
  wire [63:0] _GEN_11 = io_tlb_if2dc_dc_mode != 5'h0 ? io_tlb_if2dc_wdata : _GEN_4; // @[playground/src/noop/dcache.scala 57:50 61:29]
  wire [4:0] _GEN_12 = io_tlb_if2dc_dc_mode != 5'h0 ? io_tlb_if2dc_dc_mode : _GEN_5; // @[playground/src/noop/dcache.scala 57:50 62:29]
  wire  _GEN_14 = io_tlb_if2dc_dc_mode != 5'h0 & io_select_ready; // @[playground/src/noop/dcache.scala 57:50 64:29 23:69]
  wire  _GEN_15 = io_tlb_if2dc_dc_mode != 5'h0 ? 1'h0 : _GEN_7; // @[playground/src/noop/dcache.scala 57:50 29:69]
  wire [31:0] _GEN_18 = io_tlb_mem2dc_dc_mode != 5'h0 ? io_tlb_mem2dc_addr : _GEN_10; // @[playground/src/noop/dcache.scala 49:51 52:29]
  wire [63:0] _GEN_19 = io_tlb_mem2dc_dc_mode != 5'h0 ? io_tlb_mem2dc_wdata : _GEN_11; // @[playground/src/noop/dcache.scala 49:51 53:29]
  wire [4:0] _GEN_20 = io_tlb_mem2dc_dc_mode != 5'h0 ? io_tlb_mem2dc_dc_mode : _GEN_12; // @[playground/src/noop/dcache.scala 49:51 54:29]
  wire  _GEN_22 = io_tlb_mem2dc_dc_mode != 5'h0 & io_select_ready; // @[playground/src/noop/dcache.scala 49:51 56:29 25:69]
  wire  _GEN_23 = io_tlb_mem2dc_dc_mode != 5'h0 ? 1'h0 : _GEN_14; // @[playground/src/noop/dcache.scala 49:51 23:69]
  wire  _GEN_24 = io_tlb_mem2dc_dc_mode != 5'h0 ? 1'h0 : _GEN_15; // @[playground/src/noop/dcache.scala 49:51 29:69]
  wire [31:0] _GEN_27 = io_mem2dc_dc_mode != 5'h0 ? io_mem2dc_addr : _GEN_18; // @[playground/src/noop/dcache.scala 41:47 44:29]
  wire [63:0] _GEN_28 = io_mem2dc_dc_mode != 5'h0 ? io_mem2dc_wdata : _GEN_19; // @[playground/src/noop/dcache.scala 41:47 45:29]
  wire [4:0] _GEN_29 = io_mem2dc_dc_mode != 5'h0 ? io_mem2dc_dc_mode : _GEN_20; // @[playground/src/noop/dcache.scala 41:47 46:29]
  wire [4:0] _GEN_30 = io_mem2dc_dc_mode != 5'h0 ? io_mem2dc_amo : 5'h0; // @[playground/src/noop/dcache.scala 41:47 47:29]
  wire  _GEN_31 = io_mem2dc_dc_mode != 5'h0 & io_select_ready; // @[playground/src/noop/dcache.scala 36:25 41:47 48:29]
  wire  _GEN_32 = io_mem2dc_dc_mode != 5'h0 ? 1'h0 : _GEN_22; // @[playground/src/noop/dcache.scala 41:47 25:69]
  wire  _GEN_33 = io_mem2dc_dc_mode != 5'h0 ? 1'h0 : _GEN_23; // @[playground/src/noop/dcache.scala 41:47 23:69]
  wire  _GEN_34 = io_mem2dc_dc_mode != 5'h0 ? 1'h0 : _GEN_24; // @[playground/src/noop/dcache.scala 41:47 29:69]
  assign io_tlb_if2dc_rdata = io_select_rdata; // @[playground/src/noop/dcache.scala 22:29]
  assign io_tlb_if2dc_rvalid = io_select_rvalid & pre_idx == 2'h2; // @[playground/src/noop/dcache.scala 76:49]
  assign io_tlb_if2dc_ready = busy & ~io_select_rvalid ? 1'h0 : _GEN_33; // @[playground/src/noop/dcache.scala 40:36 23:69]
  assign io_tlb_mem2dc_rdata = io_select_rdata; // @[playground/src/noop/dcache.scala 24:29]
  assign io_tlb_mem2dc_rvalid = io_select_rvalid & pre_idx == 2'h1; // @[playground/src/noop/dcache.scala 75:49]
  assign io_tlb_mem2dc_ready = busy & ~io_select_rvalid ? 1'h0 : _GEN_32; // @[playground/src/noop/dcache.scala 40:36 25:69]
  assign io_mem2dc_rdata = io_select_rdata; // @[playground/src/noop/dcache.scala 26:29]
  assign io_mem2dc_rvalid = io_select_rvalid & pre_idx == 2'h0; // @[playground/src/noop/dcache.scala 74:49]
  assign io_mem2dc_ready = busy & ~io_select_rvalid ? 1'h0 : _GEN_31; // @[playground/src/noop/dcache.scala 36:25 40:36]
  assign io_dma2dc_rdata = io_select_rdata; // @[playground/src/noop/dcache.scala 28:29]
  assign io_dma2dc_rvalid = io_select_rvalid & pre_idx == 2'h3; // @[playground/src/noop/dcache.scala 77:49]
  assign io_dma2dc_ready = busy & ~io_select_rvalid ? 1'h0 : _GEN_34; // @[playground/src/noop/dcache.scala 40:36 29:69]
  assign io_select_addr = busy & ~io_select_rvalid ? 32'h0 : _GEN_27; // @[playground/src/noop/dcache.scala 32:25 40:36]
  assign io_select_wdata = busy & ~io_select_rvalid ? 64'h0 : _GEN_28; // @[playground/src/noop/dcache.scala 33:25 40:36]
  assign io_select_dc_mode = busy & ~io_select_rvalid ? 5'h0 : _GEN_29; // @[playground/src/noop/dcache.scala 34:25 40:36]
  assign io_select_amo = busy & ~io_select_rvalid ? 5'h0 : _GEN_30; // @[playground/src/noop/dcache.scala 35:25 40:36]
  always @(posedge clock) begin
    if (reset) begin // @[playground/src/noop/dcache.scala 30:26]
      pre_idx <= 2'h0; // @[playground/src/noop/dcache.scala 30:26]
    end else if (!(busy & ~io_select_rvalid)) begin // @[playground/src/noop/dcache.scala 40:36]
      if (io_mem2dc_dc_mode != 5'h0) begin // @[playground/src/noop/dcache.scala 41:47]
        pre_idx <= 2'h0; // @[playground/src/noop/dcache.scala 42:17]
      end else if (io_tlb_mem2dc_dc_mode != 5'h0) begin // @[playground/src/noop/dcache.scala 49:51]
        pre_idx <= 2'h1; // @[playground/src/noop/dcache.scala 50:17]
      end else begin
        pre_idx <= _GEN_8;
      end
    end
    if (reset) begin // @[playground/src/noop/dcache.scala 31:26]
      busy <= 1'h0; // @[playground/src/noop/dcache.scala 31:26]
    end else if (busy & ~io_select_rvalid) begin // @[playground/src/noop/dcache.scala 40:36]
      if (io_select_rvalid) begin // @[playground/src/noop/dcache.scala 37:27]
        busy <= 1'h0; // @[playground/src/noop/dcache.scala 38:14]
      end
    end else if (io_mem2dc_dc_mode != 5'h0) begin // @[playground/src/noop/dcache.scala 41:47]
      busy <= io_select_ready; // @[playground/src/noop/dcache.scala 43:17]
    end else if (io_tlb_mem2dc_dc_mode != 5'h0) begin // @[playground/src/noop/dcache.scala 49:51]
      busy <= io_select_ready; // @[playground/src/noop/dcache.scala 51:17]
    end else begin
      busy <= _GEN_9;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  pre_idx = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  busy = _RAND_1[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module CLINT(
  input         clock,
  input         reset,
  input  [31:0] io_rw_addr, // @[playground/src/noop/clint.scala 16:16]
  output [63:0] io_rw_rdata, // @[playground/src/noop/clint.scala 16:16]
  input  [63:0] io_rw_wdata, // @[playground/src/noop/clint.scala 16:16]
  input         io_rw_wvalid, // @[playground/src/noop/clint.scala 16:16]
  output        io_intr_raise, // @[playground/src/noop/clint.scala 16:16]
  output        io_intr_clear, // @[playground/src/noop/clint.scala 16:16]
  output        io_intr_msip_raise, // @[playground/src/noop/clint.scala 16:16]
  output        io_intr_msip_clear // @[playground/src/noop/clint.scala 16:16]
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  reg [63:0] mtime; // @[playground/src/noop/clint.scala 21:24]
  reg [63:0] mtimecmp; // @[playground/src/noop/clint.scala 22:27]
  reg [63:0] ipi; // @[playground/src/noop/clint.scala 23:22]
  reg [1:0] count; // @[playground/src/noop/clint.scala 24:24]
  reg  clear_r; // @[playground/src/noop/clint.scala 25:26]
  wire [1:0] _count_T_1 = count + 2'h1; // @[playground/src/noop/clint.scala 27:20]
  wire [63:0] _mtime_T_1 = mtime + 64'h1; // @[playground/src/noop/clint.scala 29:24]
  wire [63:0] _GEN_0 = count == 2'h0 ? _mtime_T_1 : mtime; // @[playground/src/noop/clint.scala 28:24 29:15 21:24]
  wire [63:0] _GEN_2 = io_rw_addr == 32'h200bff8 ? mtime : 64'h0; // @[playground/src/noop/clint.scala 34:17 35:31 36:24]
  wire [63:0] _GEN_6 = io_rw_addr == 32'h2004000 ? mtimecmp : _GEN_2; // @[playground/src/noop/clint.scala 41:34 42:24]
  wire  _GEN_8 = io_rw_addr == 32'h2004000 & io_rw_wvalid; // @[playground/src/noop/clint.scala 26:13 41:34]
  wire  _GEN_10 = io_rw_wvalid & io_rw_wdata[0]; // @[playground/src/noop/clint.scala 33:20 50:27 52:32]
  wire  _GEN_11 = io_rw_wvalid & ~io_rw_wdata[0]; // @[playground/src/noop/clint.scala 33:20 50:27 53:32]
  assign io_rw_rdata = io_rw_addr == 32'h2000000 ? ipi : _GEN_6; // @[playground/src/noop/clint.scala 48:29 49:24]
  assign io_intr_raise = mtime > mtimecmp; // @[playground/src/noop/clint.scala 31:28]
  assign io_intr_clear = clear_r; // @[playground/src/noop/clint.scala 32:19]
  assign io_intr_msip_raise = io_rw_addr == 32'h2000000 & _GEN_10; // @[playground/src/noop/clint.scala 33:20 48:29]
  assign io_intr_msip_clear = io_rw_addr == 32'h2000000 & _GEN_11; // @[playground/src/noop/clint.scala 33:20 48:29]
  always @(posedge clock) begin
    if (reset) begin // @[playground/src/noop/clint.scala 21:24]
      mtime <= 64'h0; // @[playground/src/noop/clint.scala 21:24]
    end else if (io_rw_addr == 32'h200bff8) begin // @[playground/src/noop/clint.scala 35:31]
      if (io_rw_wvalid) begin // @[playground/src/noop/clint.scala 37:27]
        mtime <= io_rw_wdata; // @[playground/src/noop/clint.scala 38:19]
      end else begin
        mtime <= _GEN_0;
      end
    end else begin
      mtime <= _GEN_0;
    end
    if (reset) begin // @[playground/src/noop/clint.scala 22:27]
      mtimecmp <= 64'h0; // @[playground/src/noop/clint.scala 22:27]
    end else if (io_rw_addr == 32'h2004000) begin // @[playground/src/noop/clint.scala 41:34]
      if (io_rw_wvalid) begin // @[playground/src/noop/clint.scala 43:27]
        mtimecmp <= io_rw_wdata; // @[playground/src/noop/clint.scala 44:22]
      end
    end
    if (reset) begin // @[playground/src/noop/clint.scala 23:22]
      ipi <= 64'h0; // @[playground/src/noop/clint.scala 23:22]
    end else if (io_rw_addr == 32'h2000000) begin // @[playground/src/noop/clint.scala 48:29]
      if (io_rw_wvalid) begin // @[playground/src/noop/clint.scala 50:27]
        ipi <= io_rw_wdata; // @[playground/src/noop/clint.scala 51:17]
      end
    end
    if (reset) begin // @[playground/src/noop/clint.scala 24:24]
      count <= 2'h0; // @[playground/src/noop/clint.scala 24:24]
    end else begin
      count <= _count_T_1; // @[playground/src/noop/clint.scala 27:11]
    end
    if (reset) begin // @[playground/src/noop/clint.scala 25:26]
      clear_r <= 1'h0; // @[playground/src/noop/clint.scala 25:26]
    end else begin
      clear_r <= _GEN_8;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  mtime = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  mtimecmp = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  ipi = _RAND_2[63:0];
  _RAND_3 = {1{`RANDOM}};
  count = _RAND_3[1:0];
  _RAND_4 = {1{`RANDOM}};
  clear_r = _RAND_4[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Plic(
  input         clock,
  input         reset,
  input         io_intr_in1, // @[playground/src/noop/plic.scala 28:16]
  output        io_intr_out_m_raise, // @[playground/src/noop/plic.scala 28:16]
  output        io_intr_out_m_clear, // @[playground/src/noop/plic.scala 28:16]
  output        io_intr_out_s_raise, // @[playground/src/noop/plic.scala 28:16]
  output        io_intr_out_s_clear, // @[playground/src/noop/plic.scala 28:16]
  input  [31:0] io_rw_addr, // @[playground/src/noop/plic.scala 28:16]
  output [63:0] io_rw_rdata, // @[playground/src/noop/plic.scala 28:16]
  input  [63:0] io_rw_wdata, // @[playground/src/noop/plic.scala 28:16]
  input         io_rw_wvalid, // @[playground/src/noop/plic.scala 28:16]
  input         io_rw_arvalid // @[playground/src/noop/plic.scala 28:16]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] priority_; // @[playground/src/noop/plic.scala 34:27]
  reg [31:0] pending; // @[playground/src/noop/plic.scala 35:26]
  reg [31:0] intr_enable1; // @[playground/src/noop/plic.scala 36:31]
  reg [31:0] intr_enable2; // @[playground/src/noop/plic.scala 37:31]
  reg [31:0] threshold1; // @[playground/src/noop/plic.scala 38:29]
  reg [31:0] threshold2; // @[playground/src/noop/plic.scala 39:29]
  reg [31:0] claim1; // @[playground/src/noop/plic.scala 40:25]
  reg [31:0] claim2; // @[playground/src/noop/plic.scala 41:25]
  reg  clear_r; // @[playground/src/noop/plic.scala 43:26]
  wire [63:0] _GEN_32 = {{32'd0}, pending}; // @[playground/src/noop/plic.scala 23:18]
  wire [63:0] _pending_T_1 = _GEN_32 & 64'hfffffffffffffffd; // @[playground/src/noop/plic.scala 23:18]
  wire [63:0] _pending_T_4 = _pending_T_1 | 64'h2; // @[playground/src/noop/plic.scala 23:27]
  wire [63:0] _GEN_0 = io_intr_in1 ? _pending_T_4 : {{32'd0}, pending}; // @[playground/src/noop/plic.scala 51:22 52:17 35:26]
  wire [31:0] _GEN_1 = io_intr_out_m_raise ? 32'h1 : claim1; // @[playground/src/noop/plic.scala 54:30 55:16 40:25]
  wire [31:0] _GEN_2 = io_intr_out_s_raise ? 32'h1 : claim2; // @[playground/src/noop/plic.scala 57:30 58:16 41:25]
  wire [63:0] _GEN_3 = io_rw_wvalid ? io_rw_wdata : {{32'd0}, priority_}; // @[playground/src/noop/plic.scala 63:27 64:22 34:27]
  wire [31:0] _GEN_4 = io_rw_addr == 32'hc000004 ? priority_ : 32'h0; // @[playground/src/noop/plic.scala 50:17 61:39 62:21]
  wire [63:0] _GEN_5 = io_rw_addr == 32'hc000004 ? _GEN_3 : {{32'd0}, priority_}; // @[playground/src/noop/plic.scala 34:27 61:39]
  wire [63:0] _GEN_6 = io_rw_wvalid ? io_rw_wdata : {{32'd0}, intr_enable1}; // @[playground/src/noop/plic.scala 69:27 70:26 36:31]
  wire [31:0] _GEN_7 = io_rw_addr == 32'hc002000 ? intr_enable1 : _GEN_4; // @[playground/src/noop/plic.scala 67:38 68:21]
  wire [63:0] _GEN_8 = io_rw_addr == 32'hc002000 ? _GEN_6 : {{32'd0}, intr_enable1}; // @[playground/src/noop/plic.scala 36:31 67:38]
  wire [63:0] _GEN_9 = io_rw_wvalid ? io_rw_wdata : {{32'd0}, intr_enable2}; // @[playground/src/noop/plic.scala 75:27 76:26 37:31]
  wire [31:0] _GEN_10 = io_rw_addr == 32'hc002100 ? intr_enable2 : _GEN_7; // @[playground/src/noop/plic.scala 73:38 74:21]
  wire [63:0] _GEN_11 = io_rw_addr == 32'hc002100 ? _GEN_9 : {{32'd0}, intr_enable2}; // @[playground/src/noop/plic.scala 37:31 73:38]
  wire [5:0] pending_bit_idx = claim1[5:0]; // @[playground/src/noop/plic.scala 21:26]
  wire [63:0] pending_mask_1 = 64'h1 << pending_bit_idx; // @[playground/src/noop/plic.scala 22:24]
  wire [63:0] _pending_T_5 = ~pending_mask_1; // @[playground/src/noop/plic.scala 23:20]
  wire [63:0] _pending_T_6 = _GEN_32 & _pending_T_5; // @[playground/src/noop/plic.scala 23:18]
  wire [63:0] _pending_T_7 = 64'h0 << pending_bit_idx; // @[playground/src/noop/plic.scala 23:37]
  wire [63:0] _pending_T_8 = _pending_T_7 & pending_mask_1; // @[playground/src/noop/plic.scala 23:49]
  wire [63:0] _pending_T_9 = _pending_T_6 | _pending_T_8; // @[playground/src/noop/plic.scala 23:27]
  wire [63:0] _GEN_12 = io_rw_arvalid ? _pending_T_9 : _GEN_0; // @[playground/src/noop/plic.scala 81:28 82:21]
  wire [31:0] _GEN_15 = io_rw_addr == 32'hc200004 ? claim1 : _GEN_10; // @[playground/src/noop/plic.scala 79:37 80:21]
  wire [63:0] _GEN_16 = io_rw_addr == 32'hc200004 ? _GEN_12 : _GEN_0; // @[playground/src/noop/plic.scala 79:37]
  wire  _GEN_17 = io_rw_addr == 32'hc200004 & io_rw_arvalid; // @[playground/src/noop/plic.scala 44:13 79:37]
  wire [5:0] pending_bit_idx_1 = claim2[5:0]; // @[playground/src/noop/plic.scala 21:26]
  wire [63:0] pending_mask_2 = 64'h1 << pending_bit_idx_1; // @[playground/src/noop/plic.scala 22:24]
  wire [63:0] _pending_T_10 = ~pending_mask_2; // @[playground/src/noop/plic.scala 23:20]
  wire [63:0] _pending_T_11 = _GEN_32 & _pending_T_10; // @[playground/src/noop/plic.scala 23:18]
  wire [63:0] _pending_T_12 = 64'h0 << pending_bit_idx_1; // @[playground/src/noop/plic.scala 23:37]
  wire [63:0] _pending_T_13 = _pending_T_12 & pending_mask_2; // @[playground/src/noop/plic.scala 23:49]
  wire [63:0] _pending_T_14 = _pending_T_11 | _pending_T_13; // @[playground/src/noop/plic.scala 23:27]
  wire [63:0] _GEN_19 = io_rw_arvalid ? _pending_T_14 : _GEN_16; // @[playground/src/noop/plic.scala 91:28 92:21]
  wire  _GEN_20 = io_rw_arvalid | _GEN_17; // @[playground/src/noop/plic.scala 91:28 93:21]
  wire [31:0] _GEN_22 = io_rw_addr == 32'hc201004 ? claim2 : _GEN_15; // @[playground/src/noop/plic.scala 89:37 90:21]
  wire [63:0] _GEN_23 = io_rw_addr == 32'hc201004 ? _GEN_19 : _GEN_16; // @[playground/src/noop/plic.scala 89:37]
  wire [63:0] _GEN_26 = io_rw_wvalid ? io_rw_wdata : {{32'd0}, threshold1}; // @[playground/src/noop/plic.scala 101:27 102:24 38:29]
  wire [31:0] _GEN_27 = io_rw_addr == 32'hc200000 ? threshold1 : _GEN_22; // @[playground/src/noop/plic.scala 100:21 99:41]
  wire [63:0] _GEN_28 = io_rw_addr == 32'hc200000 ? _GEN_26 : {{32'd0}, threshold1}; // @[playground/src/noop/plic.scala 38:29 99:41]
  wire [63:0] _GEN_29 = io_rw_wvalid ? io_rw_wdata : {{32'd0}, threshold2}; // @[playground/src/noop/plic.scala 107:27 108:24 39:29]
  wire [31:0] _GEN_30 = io_rw_addr == 32'hc201000 ? threshold2 : _GEN_27; // @[playground/src/noop/plic.scala 105:41 106:21]
  wire [63:0] _GEN_31 = io_rw_addr == 32'hc201000 ? _GEN_29 : {{32'd0}, threshold2}; // @[playground/src/noop/plic.scala 105:41 39:29]
  wire [63:0] _GEN_35 = reset ? 64'h0 : _GEN_5; // @[playground/src/noop/plic.scala 34:{27,27}]
  wire [63:0] _GEN_36 = reset ? 64'h0 : _GEN_23; // @[playground/src/noop/plic.scala 35:{26,26}]
  wire [63:0] _GEN_37 = reset ? 64'h0 : _GEN_8; // @[playground/src/noop/plic.scala 36:{31,31}]
  wire [63:0] _GEN_38 = reset ? 64'h0 : _GEN_11; // @[playground/src/noop/plic.scala 37:{31,31}]
  wire [63:0] _GEN_39 = reset ? 64'h0 : _GEN_28; // @[playground/src/noop/plic.scala 38:{29,29}]
  wire [63:0] _GEN_40 = reset ? 64'h0 : _GEN_31; // @[playground/src/noop/plic.scala 39:{29,29}]
  assign io_intr_out_m_raise = pending[1] & priority_ >= threshold1; // @[playground/src/noop/plic.scala 48:39]
  assign io_intr_out_m_clear = clear_r; // @[playground/src/noop/plic.scala 49:25]
  assign io_intr_out_s_raise = pending[1] & priority_ >= threshold2; // @[playground/src/noop/plic.scala 46:39]
  assign io_intr_out_s_clear = clear_r; // @[playground/src/noop/plic.scala 47:25]
  assign io_rw_rdata = {{32'd0}, _GEN_30};
  always @(posedge clock) begin
    priority_ <= _GEN_35[31:0]; // @[playground/src/noop/plic.scala 34:{27,27}]
    pending <= _GEN_36[31:0]; // @[playground/src/noop/plic.scala 35:{26,26}]
    intr_enable1 <= _GEN_37[31:0]; // @[playground/src/noop/plic.scala 36:{31,31}]
    intr_enable2 <= _GEN_38[31:0]; // @[playground/src/noop/plic.scala 37:{31,31}]
    threshold1 <= _GEN_39[31:0]; // @[playground/src/noop/plic.scala 38:{29,29}]
    threshold2 <= _GEN_40[31:0]; // @[playground/src/noop/plic.scala 39:{29,29}]
    if (reset) begin // @[playground/src/noop/plic.scala 40:25]
      claim1 <= 32'h0; // @[playground/src/noop/plic.scala 40:25]
    end else if (io_rw_addr == 32'hc200004) begin // @[playground/src/noop/plic.scala 79:37]
      if (io_rw_arvalid) begin // @[playground/src/noop/plic.scala 81:28]
        claim1 <= 32'h0; // @[playground/src/noop/plic.scala 84:20]
      end else begin
        claim1 <= _GEN_1;
      end
    end else begin
      claim1 <= _GEN_1;
    end
    if (reset) begin // @[playground/src/noop/plic.scala 41:25]
      claim2 <= 32'h0; // @[playground/src/noop/plic.scala 41:25]
    end else if (io_rw_addr == 32'hc201004) begin // @[playground/src/noop/plic.scala 89:37]
      if (io_rw_arvalid) begin // @[playground/src/noop/plic.scala 91:28]
        claim2 <= 32'h0; // @[playground/src/noop/plic.scala 94:20]
      end else begin
        claim2 <= _GEN_2;
      end
    end else begin
      claim2 <= _GEN_2;
    end
    if (reset) begin // @[playground/src/noop/plic.scala 43:26]
      clear_r <= 1'h0; // @[playground/src/noop/plic.scala 43:26]
    end else if (io_rw_addr == 32'hc201004) begin // @[playground/src/noop/plic.scala 89:37]
      clear_r <= _GEN_20;
    end else begin
      clear_r <= _GEN_17;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  priority_ = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  pending = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  intr_enable1 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  intr_enable2 = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  threshold1 = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  threshold2 = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  claim1 = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  claim2 = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  clear_r = _RAND_8[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module DmaBridge(
  input         clock,
  input         reset,
  output        io_dmaAxi_awready, // @[playground/src/noop/dma.scala 13:16]
  input         io_dmaAxi_awvalid, // @[playground/src/noop/dma.scala 13:16]
  input  [31:0] io_dmaAxi_awaddr, // @[playground/src/noop/dma.scala 13:16]
  input  [3:0]  io_dmaAxi_awid, // @[playground/src/noop/dma.scala 13:16]
  input  [7:0]  io_dmaAxi_awlen, // @[playground/src/noop/dma.scala 13:16]
  input  [2:0]  io_dmaAxi_awsize, // @[playground/src/noop/dma.scala 13:16]
  output        io_dmaAxi_wready, // @[playground/src/noop/dma.scala 13:16]
  input         io_dmaAxi_wvalid, // @[playground/src/noop/dma.scala 13:16]
  input  [63:0] io_dmaAxi_wdata, // @[playground/src/noop/dma.scala 13:16]
  input  [7:0]  io_dmaAxi_wstrb, // @[playground/src/noop/dma.scala 13:16]
  input         io_dmaAxi_bready, // @[playground/src/noop/dma.scala 13:16]
  output        io_dmaAxi_bvalid, // @[playground/src/noop/dma.scala 13:16]
  output [3:0]  io_dmaAxi_bid, // @[playground/src/noop/dma.scala 13:16]
  output        io_dmaAxi_arready, // @[playground/src/noop/dma.scala 13:16]
  input         io_dmaAxi_arvalid, // @[playground/src/noop/dma.scala 13:16]
  input  [31:0] io_dmaAxi_araddr, // @[playground/src/noop/dma.scala 13:16]
  input  [3:0]  io_dmaAxi_arid, // @[playground/src/noop/dma.scala 13:16]
  input  [7:0]  io_dmaAxi_arlen, // @[playground/src/noop/dma.scala 13:16]
  input  [2:0]  io_dmaAxi_arsize, // @[playground/src/noop/dma.scala 13:16]
  input         io_dmaAxi_rready, // @[playground/src/noop/dma.scala 13:16]
  output        io_dmaAxi_rvalid, // @[playground/src/noop/dma.scala 13:16]
  output [63:0] io_dmaAxi_rdata, // @[playground/src/noop/dma.scala 13:16]
  output        io_dmaAxi_rlast, // @[playground/src/noop/dma.scala 13:16]
  output [3:0]  io_dmaAxi_rid, // @[playground/src/noop/dma.scala 13:16]
  output [31:0] io_dcRW_addr, // @[playground/src/noop/dma.scala 13:16]
  input  [63:0] io_dcRW_rdata, // @[playground/src/noop/dma.scala 13:16]
  input         io_dcRW_rvalid, // @[playground/src/noop/dma.scala 13:16]
  output [63:0] io_dcRW_wdata, // @[playground/src/noop/dma.scala 13:16]
  output [4:0]  io_dcRW_dc_mode, // @[playground/src/noop/dma.scala 13:16]
  input         io_dcRW_ready // @[playground/src/noop/dma.scala 13:16]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [63:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
`endif // RANDOMIZE_REG_INIT
  reg [2:0] state; // @[playground/src/noop/dma.scala 18:24]
  reg  awready_r; // @[playground/src/noop/dma.scala 20:30]
  reg  wready_r; // @[playground/src/noop/dma.scala 21:30]
  reg  bvalid_r; // @[playground/src/noop/dma.scala 22:30]
  reg [3:0] bid_r; // @[playground/src/noop/dma.scala 24:30]
  reg  arready_r; // @[playground/src/noop/dma.scala 25:30]
  reg  rvalid_r; // @[playground/src/noop/dma.scala 26:30]
  reg [63:0] rdata_r; // @[playground/src/noop/dma.scala 28:30]
  reg  rlast_r; // @[playground/src/noop/dma.scala 29:30]
  reg [3:0] rid_r; // @[playground/src/noop/dma.scala 30:30]
  reg [31:0] dc_addr_r; // @[playground/src/noop/dma.scala 32:30]
  reg [63:0] dc_wdata_r; // @[playground/src/noop/dma.scala 33:30]
  reg [4:0] dc_mode_r; // @[playground/src/noop/dma.scala 34:30]
  reg [63:0] data_buf_r; // @[playground/src/noop/dma.scala 35:30]
  reg [7:0] data_strb_r; // @[playground/src/noop/dma.scala 36:30]
  reg [31:0] addr_r; // @[playground/src/noop/dma.scala 39:30]
  reg [3:0] id_r; // @[playground/src/noop/dma.scala 40:30]
  reg [7:0] len_r; // @[playground/src/noop/dma.scala 41:30]
  reg [7:0] size_r; // @[playground/src/noop/dma.scala 42:30]
  wire  _GEN_1 = io_dmaAxi_arvalid | arready_r; // @[playground/src/noop/dma.scala 48:36 50:29 25:30]
  wire  _GEN_3 = io_dmaAxi_awvalid | awready_r; // @[playground/src/noop/dma.scala 52:36 54:29 20:30]
  wire [7:0] _size_r_T = 8'h1 << io_dmaAxi_arsize; // @[playground/src/noop/dma.scala 62:32]
  wire [31:0] _dc_addr_r_T_1 = io_dmaAxi_araddr & 32'hfffffff8; // @[playground/src/noop/dma.scala 65:45]
  wire  _T_4 = io_dcRW_ready & dc_mode_r != 5'h0; // @[playground/src/noop/dma.scala 69:32]
  wire [4:0] _GEN_4 = io_dcRW_ready & dc_mode_r != 5'h0 ? 5'h0 : dc_mode_r; // @[playground/src/noop/dma.scala 69:60 70:27 34:30]
  wire [63:0] _GEN_5 = io_dcRW_rvalid ? io_dcRW_rdata : data_buf_r; // @[playground/src/noop/dma.scala 72:33 73:28 35:30]
  wire [2:0] _GEN_6 = io_dcRW_rvalid ? 3'h2 : state; // @[playground/src/noop/dma.scala 72:33 74:23 18:24]
  wire  _rlast_r_T = len_r == 8'h0; // @[playground/src/noop/dma.scala 80:30]
  wire [7:0] _len_r_T_1 = len_r - 8'h1; // @[playground/src/noop/dma.scala 88:36]
  wire [31:0] _GEN_21 = {{24'd0}, size_r}; // @[playground/src/noop/dma.scala 89:42]
  wire [31:0] _dc_addr_r_T_3 = addr_r + _GEN_21; // @[playground/src/noop/dma.scala 89:42]
  wire [31:0] _dc_addr_r_T_5 = _dc_addr_r_T_3 & 32'hfffffff8; // @[playground/src/noop/dma.scala 89:52]
  wire [2:0] _GEN_7 = rlast_r ? 3'h0 : 3'h6; // @[playground/src/noop/dma.scala 85:30 86:27 92:27]
  wire [7:0] _GEN_8 = rlast_r ? len_r : _len_r_T_1; // @[playground/src/noop/dma.scala 41:30 85:30 88:27]
  wire [31:0] _GEN_9 = rlast_r ? dc_addr_r : _dc_addr_r_T_5; // @[playground/src/noop/dma.scala 32:30 85:30 89:31]
  wire [31:0] _GEN_10 = rlast_r ? addr_r : _dc_addr_r_T_3; // @[playground/src/noop/dma.scala 39:30 85:30 90:28]
  wire [4:0] _GEN_11 = rlast_r ? dc_mode_r : 5'h7; // @[playground/src/noop/dma.scala 34:30 85:30 91:31]
  wire  _GEN_12 = io_dmaAxi_rready & rvalid_r ? 1'h0 : 1'h1; // @[playground/src/noop/dma.scala 79:22 83:47 84:26]
  wire [2:0] _GEN_13 = io_dmaAxi_rready & rvalid_r ? _GEN_7 : state; // @[playground/src/noop/dma.scala 18:24 83:47]
  wire [7:0] _GEN_14 = io_dmaAxi_rready & rvalid_r ? _GEN_8 : len_r; // @[playground/src/noop/dma.scala 41:30 83:47]
  wire [31:0] _GEN_15 = io_dmaAxi_rready & rvalid_r ? _GEN_9 : dc_addr_r; // @[playground/src/noop/dma.scala 32:30 83:47]
  wire [31:0] _GEN_16 = io_dmaAxi_rready & rvalid_r ? _GEN_10 : addr_r; // @[playground/src/noop/dma.scala 39:30 83:47]
  wire [4:0] _GEN_17 = io_dmaAxi_rready & rvalid_r ? _GEN_11 : dc_mode_r; // @[playground/src/noop/dma.scala 34:30 83:47]
  wire [31:0] _dc_addr_r_T_7 = io_dmaAxi_awaddr & 32'hfffffff8; // @[playground/src/noop/dma.scala 99:45]
  wire [7:0] _size_r_T_1 = 8'h1 << io_dmaAxi_awsize; // @[playground/src/noop/dma.scala 102:32]
  wire  _GEN_18 = io_dmaAxi_wvalid & wready_r ? 1'h0 : wready_r; // @[playground/src/noop/dma.scala 108:47 109:29 21:30]
  wire [63:0] _GEN_19 = io_dmaAxi_wvalid & wready_r ? io_dmaAxi_wdata : data_buf_r; // @[playground/src/noop/dma.scala 108:47 110:29 35:30]
  wire [7:0] _GEN_20 = io_dmaAxi_wvalid & wready_r ? io_dmaAxi_wstrb : data_strb_r; // @[playground/src/noop/dma.scala 108:47 111:29 36:30]
  wire [2:0] _GEN_22 = io_dmaAxi_wvalid & wready_r ? 3'h7 : state; // @[playground/src/noop/dma.scala 108:47 113:29 18:24]
  wire  _GEN_23 = _rlast_r_T | bvalid_r; // @[playground/src/noop/dma.scala 120:36 121:30 22:30]
  wire [3:0] _GEN_25 = _rlast_r_T ? id_r : bid_r; // @[playground/src/noop/dma.scala 120:36 123:29 24:30]
  wire [2:0] _GEN_26 = _rlast_r_T ? 3'h5 : 3'h4; // @[playground/src/noop/dma.scala 120:36 124:29 126:27]
  wire  _GEN_27 = _rlast_r_T ? wready_r : 1'h1; // @[playground/src/noop/dma.scala 120:36 127:30 21:30]
  wire [7:0] _GEN_28 = _rlast_r_T ? len_r : _len_r_T_1; // @[playground/src/noop/dma.scala 120:36 128:27 41:30]
  wire [7:0] _data_strb_r_T = {{1'd0}, data_strb_r[7:1]}; // @[playground/src/noop/dma.scala 135:48]
  wire [63:0] _data_buf_r_T = {{8'd0}, data_buf_r[63:8]}; // @[playground/src/noop/dma.scala 136:47]
  wire [31:0] _dc_addr_r_T_13 = dc_addr_r + 32'h1; // @[playground/src/noop/dma.scala 137:46]
  wire [4:0] _GEN_29 = data_strb_r[0] ? 5'h8 : dc_mode_r; // @[playground/src/noop/dma.scala 131:37 132:33 34:30]
  wire [63:0] _GEN_30 = data_strb_r[0] ? data_buf_r : dc_wdata_r; // @[playground/src/noop/dma.scala 131:37 133:33 33:30]
  wire [7:0] _GEN_31 = data_strb_r[0] ? data_strb_r : _data_strb_r_T; // @[playground/src/noop/dma.scala 131:37 36:30 135:33]
  wire [63:0] _GEN_32 = data_strb_r[0] ? data_buf_r : _data_buf_r_T; // @[playground/src/noop/dma.scala 131:37 35:30 136:33]
  wire [31:0] _GEN_33 = data_strb_r[0] ? dc_addr_r : _dc_addr_r_T_13; // @[playground/src/noop/dma.scala 131:37 32:30 137:33]
  wire [4:0] _GEN_35 = _T_4 ? 5'h0 : _GEN_29; // @[playground/src/noop/dma.scala 140:62 141:33]
  wire [7:0] _GEN_36 = _T_4 ? _data_strb_r_T : _GEN_31; // @[playground/src/noop/dma.scala 140:62 142:33]
  wire [63:0] _GEN_37 = _T_4 ? _data_buf_r_T : _GEN_32; // @[playground/src/noop/dma.scala 140:62 143:33]
  wire [31:0] _GEN_38 = _T_4 ? _dc_addr_r_T_13 : _GEN_33; // @[playground/src/noop/dma.scala 140:62 144:33]
  wire [31:0] _GEN_40 = data_strb_r == 8'h0 ? _dc_addr_r_T_3 : addr_r; // @[playground/src/noop/dma.scala 117:38 118:24 39:30]
  wire [31:0] _GEN_41 = data_strb_r == 8'h0 ? _dc_addr_r_T_5 : _GEN_38; // @[playground/src/noop/dma.scala 117:38 119:27]
  wire  _GEN_42 = data_strb_r == 8'h0 ? _GEN_23 : bvalid_r; // @[playground/src/noop/dma.scala 117:38 22:30]
  wire [3:0] _GEN_44 = data_strb_r == 8'h0 ? _GEN_25 : bid_r; // @[playground/src/noop/dma.scala 117:38 24:30]
  wire [2:0] _GEN_45 = data_strb_r == 8'h0 ? _GEN_26 : state; // @[playground/src/noop/dma.scala 117:38 18:24]
  wire  _GEN_46 = data_strb_r == 8'h0 ? _GEN_27 : wready_r; // @[playground/src/noop/dma.scala 117:38 21:30]
  wire [7:0] _GEN_47 = data_strb_r == 8'h0 ? _GEN_28 : len_r; // @[playground/src/noop/dma.scala 117:38 41:30]
  wire [4:0] _GEN_48 = data_strb_r == 8'h0 ? dc_mode_r : _GEN_35; // @[playground/src/noop/dma.scala 117:38 34:30]
  wire [63:0] _GEN_49 = data_strb_r == 8'h0 ? dc_wdata_r : _GEN_30; // @[playground/src/noop/dma.scala 117:38 33:30]
  wire [7:0] _GEN_50 = data_strb_r == 8'h0 ? data_strb_r : _GEN_36; // @[playground/src/noop/dma.scala 117:38 36:30]
  wire [63:0] _GEN_51 = data_strb_r == 8'h0 ? data_buf_r : _GEN_37; // @[playground/src/noop/dma.scala 117:38 35:30]
  wire [2:0] _GEN_53 = io_dmaAxi_bready & bvalid_r ? 3'h0 : state; // @[playground/src/noop/dma.scala 150:47 151:23 18:24]
  wire [2:0] _GEN_55 = 3'h5 == state ? _GEN_53 : state; // @[playground/src/noop/dma.scala 46:18 18:24]
  wire [31:0] _GEN_57 = 3'h7 == state ? _GEN_40 : addr_r; // @[playground/src/noop/dma.scala 46:18 39:30]
  wire [31:0] _GEN_58 = 3'h7 == state ? _GEN_41 : dc_addr_r; // @[playground/src/noop/dma.scala 46:18 32:30]
  wire  _GEN_59 = 3'h7 == state ? _GEN_42 : bvalid_r; // @[playground/src/noop/dma.scala 46:18 22:30]
  wire [3:0] _GEN_61 = 3'h7 == state ? _GEN_44 : bid_r; // @[playground/src/noop/dma.scala 46:18 24:30]
  wire [2:0] _GEN_62 = 3'h7 == state ? _GEN_45 : _GEN_55; // @[playground/src/noop/dma.scala 46:18]
  wire  _GEN_63 = 3'h7 == state ? _GEN_46 : wready_r; // @[playground/src/noop/dma.scala 46:18 21:30]
  wire [7:0] _GEN_64 = 3'h7 == state ? _GEN_47 : len_r; // @[playground/src/noop/dma.scala 46:18 41:30]
  wire [4:0] _GEN_65 = 3'h7 == state ? _GEN_48 : dc_mode_r; // @[playground/src/noop/dma.scala 46:18 34:30]
  wire [63:0] _GEN_66 = 3'h7 == state ? _GEN_49 : dc_wdata_r; // @[playground/src/noop/dma.scala 46:18 33:30]
  wire [7:0] _GEN_67 = 3'h7 == state ? _GEN_50 : data_strb_r; // @[playground/src/noop/dma.scala 46:18 36:30]
  wire [63:0] _GEN_68 = 3'h7 == state ? _GEN_51 : data_buf_r; // @[playground/src/noop/dma.scala 46:18 35:30]
  wire  _GEN_70 = 3'h4 == state ? _GEN_18 : _GEN_63; // @[playground/src/noop/dma.scala 46:18]
  wire [63:0] _GEN_71 = 3'h4 == state ? _GEN_19 : _GEN_68; // @[playground/src/noop/dma.scala 46:18]
  wire [7:0] _GEN_72 = 3'h4 == state ? _GEN_20 : _GEN_67; // @[playground/src/noop/dma.scala 46:18]
  wire [2:0] _GEN_74 = 3'h4 == state ? _GEN_22 : _GEN_62; // @[playground/src/noop/dma.scala 46:18]
  wire [31:0] _GEN_75 = 3'h4 == state ? addr_r : _GEN_57; // @[playground/src/noop/dma.scala 46:18 39:30]
  wire [31:0] _GEN_76 = 3'h4 == state ? dc_addr_r : _GEN_58; // @[playground/src/noop/dma.scala 46:18 32:30]
  wire  _GEN_77 = 3'h4 == state ? bvalid_r : _GEN_59; // @[playground/src/noop/dma.scala 46:18 22:30]
  wire [3:0] _GEN_79 = 3'h4 == state ? bid_r : _GEN_61; // @[playground/src/noop/dma.scala 46:18 24:30]
  wire [7:0] _GEN_80 = 3'h4 == state ? len_r : _GEN_64; // @[playground/src/noop/dma.scala 46:18 41:30]
  wire [4:0] _GEN_81 = 3'h4 == state ? dc_mode_r : _GEN_65; // @[playground/src/noop/dma.scala 46:18 34:30]
  wire [63:0] _GEN_82 = 3'h4 == state ? dc_wdata_r : _GEN_66; // @[playground/src/noop/dma.scala 46:18 33:30]
  wire  _GEN_83 = 3'h3 == state ? 1'h0 : awready_r; // @[playground/src/noop/dma.scala 46:18 97:25 20:30]
  wire [31:0] _GEN_84 = 3'h3 == state ? io_dmaAxi_awaddr : _GEN_75; // @[playground/src/noop/dma.scala 46:18 98:25]
  wire [31:0] _GEN_85 = 3'h3 == state ? _dc_addr_r_T_7 : _GEN_76; // @[playground/src/noop/dma.scala 46:18 99:25]
  wire [3:0] _GEN_86 = 3'h3 == state ? io_dmaAxi_awid : id_r; // @[playground/src/noop/dma.scala 46:18 100:25 40:30]
  wire [7:0] _GEN_87 = 3'h3 == state ? io_dmaAxi_awlen : _GEN_80; // @[playground/src/noop/dma.scala 46:18 101:25]
  wire [7:0] _GEN_88 = 3'h3 == state ? _size_r_T_1 : size_r; // @[playground/src/noop/dma.scala 46:18 102:25 42:30]
  wire  _GEN_90 = 3'h3 == state | _GEN_70; // @[playground/src/noop/dma.scala 46:18 104:25]
  wire [2:0] _GEN_91 = 3'h3 == state ? 3'h4 : _GEN_74; // @[playground/src/noop/dma.scala 46:18 105:25]
  wire [63:0] _GEN_92 = 3'h3 == state ? data_buf_r : _GEN_71; // @[playground/src/noop/dma.scala 46:18 35:30]
  wire [7:0] _GEN_93 = 3'h3 == state ? data_strb_r : _GEN_72; // @[playground/src/noop/dma.scala 46:18 36:30]
  wire  _GEN_95 = 3'h3 == state ? bvalid_r : _GEN_77; // @[playground/src/noop/dma.scala 46:18 22:30]
  wire [3:0] _GEN_97 = 3'h3 == state ? bid_r : _GEN_79; // @[playground/src/noop/dma.scala 46:18 24:30]
  wire [4:0] _GEN_98 = 3'h3 == state ? dc_mode_r : _GEN_81; // @[playground/src/noop/dma.scala 46:18 34:30]
  wire [63:0] _GEN_99 = 3'h3 == state ? dc_wdata_r : _GEN_82; // @[playground/src/noop/dma.scala 46:18 33:30]
  wire [63:0] _GEN_100 = 3'h2 == state ? data_buf_r : rdata_r; // @[playground/src/noop/dma.scala 46:18 78:21 28:30]
  wire  _GEN_101 = 3'h2 == state ? _GEN_12 : rvalid_r; // @[playground/src/noop/dma.scala 46:18 26:30]
  wire  _GEN_102 = 3'h2 == state ? len_r == 8'h0 : rlast_r; // @[playground/src/noop/dma.scala 46:18 80:21 29:30]
  wire [3:0] _GEN_103 = 3'h2 == state ? id_r : rid_r; // @[playground/src/noop/dma.scala 46:18 81:21 30:30]
  wire [2:0] _GEN_105 = 3'h2 == state ? _GEN_13 : _GEN_91; // @[playground/src/noop/dma.scala 46:18]
  wire [7:0] _GEN_106 = 3'h2 == state ? _GEN_14 : _GEN_87; // @[playground/src/noop/dma.scala 46:18]
  wire [31:0] _GEN_107 = 3'h2 == state ? _GEN_15 : _GEN_85; // @[playground/src/noop/dma.scala 46:18]
  wire [31:0] _GEN_108 = 3'h2 == state ? _GEN_16 : _GEN_84; // @[playground/src/noop/dma.scala 46:18]
  wire [4:0] _GEN_109 = 3'h2 == state ? _GEN_17 : _GEN_98; // @[playground/src/noop/dma.scala 46:18]
  wire  _GEN_110 = 3'h2 == state ? awready_r : _GEN_83; // @[playground/src/noop/dma.scala 46:18 20:30]
  wire [3:0] _GEN_111 = 3'h2 == state ? id_r : _GEN_86; // @[playground/src/noop/dma.scala 46:18 40:30]
  wire [7:0] _GEN_112 = 3'h2 == state ? size_r : _GEN_88; // @[playground/src/noop/dma.scala 46:18 42:30]
  wire  _GEN_114 = 3'h2 == state ? wready_r : _GEN_90; // @[playground/src/noop/dma.scala 46:18 21:30]
  wire [63:0] _GEN_115 = 3'h2 == state ? data_buf_r : _GEN_92; // @[playground/src/noop/dma.scala 46:18 35:30]
  wire [7:0] _GEN_116 = 3'h2 == state ? data_strb_r : _GEN_93; // @[playground/src/noop/dma.scala 46:18 36:30]
  wire  _GEN_118 = 3'h2 == state ? bvalid_r : _GEN_95; // @[playground/src/noop/dma.scala 46:18 22:30]
  wire [3:0] _GEN_120 = 3'h2 == state ? bid_r : _GEN_97; // @[playground/src/noop/dma.scala 46:18 24:30]
  wire [63:0] _GEN_121 = 3'h2 == state ? dc_wdata_r : _GEN_99; // @[playground/src/noop/dma.scala 46:18 33:30]
  assign io_dmaAxi_awready = awready_r; // @[playground/src/noop/dma.scala 156:25]
  assign io_dmaAxi_wready = wready_r; // @[playground/src/noop/dma.scala 157:25]
  assign io_dmaAxi_bvalid = bvalid_r; // @[playground/src/noop/dma.scala 158:25]
  assign io_dmaAxi_bid = bid_r; // @[playground/src/noop/dma.scala 160:25]
  assign io_dmaAxi_arready = arready_r; // @[playground/src/noop/dma.scala 161:25]
  assign io_dmaAxi_rvalid = rvalid_r; // @[playground/src/noop/dma.scala 162:25]
  assign io_dmaAxi_rdata = rdata_r; // @[playground/src/noop/dma.scala 164:25]
  assign io_dmaAxi_rlast = rlast_r; // @[playground/src/noop/dma.scala 165:25]
  assign io_dmaAxi_rid = rid_r; // @[playground/src/noop/dma.scala 166:25]
  assign io_dcRW_addr = dc_addr_r; // @[playground/src/noop/dma.scala 168:21]
  assign io_dcRW_wdata = dc_wdata_r; // @[playground/src/noop/dma.scala 169:21]
  assign io_dcRW_dc_mode = dc_mode_r; // @[playground/src/noop/dma.scala 170:21]
  always @(posedge clock) begin
    if (reset) begin // @[playground/src/noop/dma.scala 18:24]
      state <= 3'h0; // @[playground/src/noop/dma.scala 18:24]
    end else if (3'h0 == state) begin // @[playground/src/noop/dma.scala 46:18]
      if (io_dmaAxi_awvalid) begin // @[playground/src/noop/dma.scala 52:36]
        state <= 3'h3; // @[playground/src/noop/dma.scala 53:29]
      end else if (io_dmaAxi_arvalid) begin // @[playground/src/noop/dma.scala 48:36]
        state <= 3'h1; // @[playground/src/noop/dma.scala 49:29]
      end
    end else if (3'h1 == state) begin // @[playground/src/noop/dma.scala 46:18]
      state <= 3'h6; // @[playground/src/noop/dma.scala 64:25]
    end else if (3'h6 == state) begin // @[playground/src/noop/dma.scala 46:18]
      state <= _GEN_6;
    end else begin
      state <= _GEN_105;
    end
    if (reset) begin // @[playground/src/noop/dma.scala 20:30]
      awready_r <= 1'h0; // @[playground/src/noop/dma.scala 20:30]
    end else if (3'h0 == state) begin // @[playground/src/noop/dma.scala 46:18]
      awready_r <= _GEN_3;
    end else if (!(3'h1 == state)) begin // @[playground/src/noop/dma.scala 46:18]
      if (!(3'h6 == state)) begin // @[playground/src/noop/dma.scala 46:18]
        awready_r <= _GEN_110;
      end
    end
    if (reset) begin // @[playground/src/noop/dma.scala 21:30]
      wready_r <= 1'h0; // @[playground/src/noop/dma.scala 21:30]
    end else if (!(3'h0 == state)) begin // @[playground/src/noop/dma.scala 46:18]
      if (!(3'h1 == state)) begin // @[playground/src/noop/dma.scala 46:18]
        if (!(3'h6 == state)) begin // @[playground/src/noop/dma.scala 46:18]
          wready_r <= _GEN_114;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/dma.scala 22:30]
      bvalid_r <= 1'h0; // @[playground/src/noop/dma.scala 22:30]
    end else if (!(3'h0 == state)) begin // @[playground/src/noop/dma.scala 46:18]
      if (!(3'h1 == state)) begin // @[playground/src/noop/dma.scala 46:18]
        if (!(3'h6 == state)) begin // @[playground/src/noop/dma.scala 46:18]
          bvalid_r <= _GEN_118;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/dma.scala 24:30]
      bid_r <= 4'h0; // @[playground/src/noop/dma.scala 24:30]
    end else if (!(3'h0 == state)) begin // @[playground/src/noop/dma.scala 46:18]
      if (!(3'h1 == state)) begin // @[playground/src/noop/dma.scala 46:18]
        if (!(3'h6 == state)) begin // @[playground/src/noop/dma.scala 46:18]
          bid_r <= _GEN_120;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/dma.scala 25:30]
      arready_r <= 1'h0; // @[playground/src/noop/dma.scala 25:30]
    end else if (3'h0 == state) begin // @[playground/src/noop/dma.scala 46:18]
      arready_r <= _GEN_1;
    end else if (3'h1 == state) begin // @[playground/src/noop/dma.scala 46:18]
      arready_r <= 1'h0; // @[playground/src/noop/dma.scala 58:25]
    end
    if (reset) begin // @[playground/src/noop/dma.scala 26:30]
      rvalid_r <= 1'h0; // @[playground/src/noop/dma.scala 26:30]
    end else if (!(3'h0 == state)) begin // @[playground/src/noop/dma.scala 46:18]
      if (!(3'h1 == state)) begin // @[playground/src/noop/dma.scala 46:18]
        if (!(3'h6 == state)) begin // @[playground/src/noop/dma.scala 46:18]
          rvalid_r <= _GEN_101;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/dma.scala 28:30]
      rdata_r <= 64'h0; // @[playground/src/noop/dma.scala 28:30]
    end else if (!(3'h0 == state)) begin // @[playground/src/noop/dma.scala 46:18]
      if (!(3'h1 == state)) begin // @[playground/src/noop/dma.scala 46:18]
        if (!(3'h6 == state)) begin // @[playground/src/noop/dma.scala 46:18]
          rdata_r <= _GEN_100;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/dma.scala 29:30]
      rlast_r <= 1'h0; // @[playground/src/noop/dma.scala 29:30]
    end else if (!(3'h0 == state)) begin // @[playground/src/noop/dma.scala 46:18]
      if (!(3'h1 == state)) begin // @[playground/src/noop/dma.scala 46:18]
        if (!(3'h6 == state)) begin // @[playground/src/noop/dma.scala 46:18]
          rlast_r <= _GEN_102;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/dma.scala 30:30]
      rid_r <= 4'h0; // @[playground/src/noop/dma.scala 30:30]
    end else if (!(3'h0 == state)) begin // @[playground/src/noop/dma.scala 46:18]
      if (!(3'h1 == state)) begin // @[playground/src/noop/dma.scala 46:18]
        if (!(3'h6 == state)) begin // @[playground/src/noop/dma.scala 46:18]
          rid_r <= _GEN_103;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/dma.scala 32:30]
      dc_addr_r <= 32'h0; // @[playground/src/noop/dma.scala 32:30]
    end else if (!(3'h0 == state)) begin // @[playground/src/noop/dma.scala 46:18]
      if (3'h1 == state) begin // @[playground/src/noop/dma.scala 46:18]
        dc_addr_r <= _dc_addr_r_T_1; // @[playground/src/noop/dma.scala 65:25]
      end else if (!(3'h6 == state)) begin // @[playground/src/noop/dma.scala 46:18]
        dc_addr_r <= _GEN_107;
      end
    end
    if (reset) begin // @[playground/src/noop/dma.scala 33:30]
      dc_wdata_r <= 64'h0; // @[playground/src/noop/dma.scala 33:30]
    end else if (!(3'h0 == state)) begin // @[playground/src/noop/dma.scala 46:18]
      if (!(3'h1 == state)) begin // @[playground/src/noop/dma.scala 46:18]
        if (!(3'h6 == state)) begin // @[playground/src/noop/dma.scala 46:18]
          dc_wdata_r <= _GEN_121;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/dma.scala 34:30]
      dc_mode_r <= 5'h0; // @[playground/src/noop/dma.scala 34:30]
    end else if (!(3'h0 == state)) begin // @[playground/src/noop/dma.scala 46:18]
      if (3'h1 == state) begin // @[playground/src/noop/dma.scala 46:18]
        dc_mode_r <= 5'h7; // @[playground/src/noop/dma.scala 66:25]
      end else if (3'h6 == state) begin // @[playground/src/noop/dma.scala 46:18]
        dc_mode_r <= _GEN_4;
      end else begin
        dc_mode_r <= _GEN_109;
      end
    end
    if (reset) begin // @[playground/src/noop/dma.scala 35:30]
      data_buf_r <= 64'h0; // @[playground/src/noop/dma.scala 35:30]
    end else if (!(3'h0 == state)) begin // @[playground/src/noop/dma.scala 46:18]
      if (!(3'h1 == state)) begin // @[playground/src/noop/dma.scala 46:18]
        if (3'h6 == state) begin // @[playground/src/noop/dma.scala 46:18]
          data_buf_r <= _GEN_5;
        end else begin
          data_buf_r <= _GEN_115;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/dma.scala 36:30]
      data_strb_r <= 8'h0; // @[playground/src/noop/dma.scala 36:30]
    end else if (!(3'h0 == state)) begin // @[playground/src/noop/dma.scala 46:18]
      if (!(3'h1 == state)) begin // @[playground/src/noop/dma.scala 46:18]
        if (!(3'h6 == state)) begin // @[playground/src/noop/dma.scala 46:18]
          data_strb_r <= _GEN_116;
        end
      end
    end
    if (reset) begin // @[playground/src/noop/dma.scala 39:30]
      addr_r <= 32'h0; // @[playground/src/noop/dma.scala 39:30]
    end else if (!(3'h0 == state)) begin // @[playground/src/noop/dma.scala 46:18]
      if (3'h1 == state) begin // @[playground/src/noop/dma.scala 46:18]
        addr_r <= io_dmaAxi_araddr; // @[playground/src/noop/dma.scala 59:25]
      end else if (!(3'h6 == state)) begin // @[playground/src/noop/dma.scala 46:18]
        addr_r <= _GEN_108;
      end
    end
    if (reset) begin // @[playground/src/noop/dma.scala 40:30]
      id_r <= 4'h0; // @[playground/src/noop/dma.scala 40:30]
    end else if (!(3'h0 == state)) begin // @[playground/src/noop/dma.scala 46:18]
      if (3'h1 == state) begin // @[playground/src/noop/dma.scala 46:18]
        id_r <= io_dmaAxi_arid; // @[playground/src/noop/dma.scala 60:25]
      end else if (!(3'h6 == state)) begin // @[playground/src/noop/dma.scala 46:18]
        id_r <= _GEN_111;
      end
    end
    if (reset) begin // @[playground/src/noop/dma.scala 41:30]
      len_r <= 8'h0; // @[playground/src/noop/dma.scala 41:30]
    end else if (!(3'h0 == state)) begin // @[playground/src/noop/dma.scala 46:18]
      if (3'h1 == state) begin // @[playground/src/noop/dma.scala 46:18]
        len_r <= io_dmaAxi_arlen; // @[playground/src/noop/dma.scala 61:25]
      end else if (!(3'h6 == state)) begin // @[playground/src/noop/dma.scala 46:18]
        len_r <= _GEN_106;
      end
    end
    if (reset) begin // @[playground/src/noop/dma.scala 42:30]
      size_r <= 8'h0; // @[playground/src/noop/dma.scala 42:30]
    end else if (!(3'h0 == state)) begin // @[playground/src/noop/dma.scala 46:18]
      if (3'h1 == state) begin // @[playground/src/noop/dma.scala 46:18]
        size_r <= _size_r_T; // @[playground/src/noop/dma.scala 62:25]
      end else if (!(3'h6 == state)) begin // @[playground/src/noop/dma.scala 46:18]
        size_r <= _GEN_112;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  awready_r = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  wready_r = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  bvalid_r = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  bid_r = _RAND_4[3:0];
  _RAND_5 = {1{`RANDOM}};
  arready_r = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  rvalid_r = _RAND_6[0:0];
  _RAND_7 = {2{`RANDOM}};
  rdata_r = _RAND_7[63:0];
  _RAND_8 = {1{`RANDOM}};
  rlast_r = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  rid_r = _RAND_9[3:0];
  _RAND_10 = {1{`RANDOM}};
  dc_addr_r = _RAND_10[31:0];
  _RAND_11 = {2{`RANDOM}};
  dc_wdata_r = _RAND_11[63:0];
  _RAND_12 = {1{`RANDOM}};
  dc_mode_r = _RAND_12[4:0];
  _RAND_13 = {2{`RANDOM}};
  data_buf_r = _RAND_13[63:0];
  _RAND_14 = {1{`RANDOM}};
  data_strb_r = _RAND_14[7:0];
  _RAND_15 = {1{`RANDOM}};
  addr_r = _RAND_15[31:0];
  _RAND_16 = {1{`RANDOM}};
  id_r = _RAND_16[3:0];
  _RAND_17 = {1{`RANDOM}};
  len_r = _RAND_17[7:0];
  _RAND_18 = {1{`RANDOM}};
  size_r = _RAND_18[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module CPU(
  input         clock,
  input         reset,
  input         io_master_awready, // @[playground/src/noop/cpu.scala 94:16]
  output        io_master_awvalid, // @[playground/src/noop/cpu.scala 94:16]
  output [31:0] io_master_awaddr, // @[playground/src/noop/cpu.scala 94:16]
  output [3:0]  io_master_awid, // @[playground/src/noop/cpu.scala 94:16]
  output [7:0]  io_master_awlen, // @[playground/src/noop/cpu.scala 94:16]
  output [2:0]  io_master_awsize, // @[playground/src/noop/cpu.scala 94:16]
  output [1:0]  io_master_awburst, // @[playground/src/noop/cpu.scala 94:16]
  input         io_master_wready, // @[playground/src/noop/cpu.scala 94:16]
  output        io_master_wvalid, // @[playground/src/noop/cpu.scala 94:16]
  output [63:0] io_master_wdata, // @[playground/src/noop/cpu.scala 94:16]
  output [7:0]  io_master_wstrb, // @[playground/src/noop/cpu.scala 94:16]
  output        io_master_wlast, // @[playground/src/noop/cpu.scala 94:16]
  output        io_master_bready, // @[playground/src/noop/cpu.scala 94:16]
  input         io_master_bvalid, // @[playground/src/noop/cpu.scala 94:16]
  input  [1:0]  io_master_bresp, // @[playground/src/noop/cpu.scala 94:16]
  input  [3:0]  io_master_bid, // @[playground/src/noop/cpu.scala 94:16]
  input         io_master_arready, // @[playground/src/noop/cpu.scala 94:16]
  output        io_master_arvalid, // @[playground/src/noop/cpu.scala 94:16]
  output [31:0] io_master_araddr, // @[playground/src/noop/cpu.scala 94:16]
  output [3:0]  io_master_arid, // @[playground/src/noop/cpu.scala 94:16]
  output [7:0]  io_master_arlen, // @[playground/src/noop/cpu.scala 94:16]
  output [2:0]  io_master_arsize, // @[playground/src/noop/cpu.scala 94:16]
  output [1:0]  io_master_arburst, // @[playground/src/noop/cpu.scala 94:16]
  output        io_master_rready, // @[playground/src/noop/cpu.scala 94:16]
  input         io_master_rvalid, // @[playground/src/noop/cpu.scala 94:16]
  input  [1:0]  io_master_rresp, // @[playground/src/noop/cpu.scala 94:16]
  input  [63:0] io_master_rdata, // @[playground/src/noop/cpu.scala 94:16]
  input         io_master_rlast, // @[playground/src/noop/cpu.scala 94:16]
  input  [3:0]  io_master_rid, // @[playground/src/noop/cpu.scala 94:16]
  output        io_slave_awready, // @[playground/src/noop/cpu.scala 94:16]
  input         io_slave_awvalid, // @[playground/src/noop/cpu.scala 94:16]
  input  [31:0] io_slave_awaddr, // @[playground/src/noop/cpu.scala 94:16]
  input  [3:0]  io_slave_awid, // @[playground/src/noop/cpu.scala 94:16]
  input  [7:0]  io_slave_awlen, // @[playground/src/noop/cpu.scala 94:16]
  input  [2:0]  io_slave_awsize, // @[playground/src/noop/cpu.scala 94:16]
  input  [1:0]  io_slave_awburst, // @[playground/src/noop/cpu.scala 94:16]
  output        io_slave_wready, // @[playground/src/noop/cpu.scala 94:16]
  input         io_slave_wvalid, // @[playground/src/noop/cpu.scala 94:16]
  input  [63:0] io_slave_wdata, // @[playground/src/noop/cpu.scala 94:16]
  input  [7:0]  io_slave_wstrb, // @[playground/src/noop/cpu.scala 94:16]
  input         io_slave_wlast, // @[playground/src/noop/cpu.scala 94:16]
  input         io_slave_bready, // @[playground/src/noop/cpu.scala 94:16]
  output        io_slave_bvalid, // @[playground/src/noop/cpu.scala 94:16]
  output [1:0]  io_slave_bresp, // @[playground/src/noop/cpu.scala 94:16]
  output [3:0]  io_slave_bid, // @[playground/src/noop/cpu.scala 94:16]
  output        io_slave_arready, // @[playground/src/noop/cpu.scala 94:16]
  input         io_slave_arvalid, // @[playground/src/noop/cpu.scala 94:16]
  input  [31:0] io_slave_araddr, // @[playground/src/noop/cpu.scala 94:16]
  input  [3:0]  io_slave_arid, // @[playground/src/noop/cpu.scala 94:16]
  input  [7:0]  io_slave_arlen, // @[playground/src/noop/cpu.scala 94:16]
  input  [2:0]  io_slave_arsize, // @[playground/src/noop/cpu.scala 94:16]
  input  [1:0]  io_slave_arburst, // @[playground/src/noop/cpu.scala 94:16]
  input         io_slave_rready, // @[playground/src/noop/cpu.scala 94:16]
  output        io_slave_rvalid, // @[playground/src/noop/cpu.scala 94:16]
  output [1:0]  io_slave_rresp, // @[playground/src/noop/cpu.scala 94:16]
  output [63:0] io_slave_rdata, // @[playground/src/noop/cpu.scala 94:16]
  output        io_slave_rlast, // @[playground/src/noop/cpu.scala 94:16]
  output [3:0]  io_slave_rid, // @[playground/src/noop/cpu.scala 94:16]
  input         io_interrupt // @[playground/src/noop/cpu.scala 94:16]
);
  wire  fetch_clock; // @[playground/src/noop/cpu.scala 96:29]
  wire  fetch_reset; // @[playground/src/noop/cpu.scala 96:29]
  wire [31:0] fetch_io_instRead_addr; // @[playground/src/noop/cpu.scala 96:29]
  wire [63:0] fetch_io_instRead_inst; // @[playground/src/noop/cpu.scala 96:29]
  wire  fetch_io_instRead_arvalid; // @[playground/src/noop/cpu.scala 96:29]
  wire  fetch_io_instRead_rvalid; // @[playground/src/noop/cpu.scala 96:29]
  wire [63:0] fetch_io_va2pa_vaddr; // @[playground/src/noop/cpu.scala 96:29]
  wire  fetch_io_va2pa_vvalid; // @[playground/src/noop/cpu.scala 96:29]
  wire [31:0] fetch_io_va2pa_paddr; // @[playground/src/noop/cpu.scala 96:29]
  wire  fetch_io_va2pa_pvalid; // @[playground/src/noop/cpu.scala 96:29]
  wire [63:0] fetch_io_va2pa_tlb_excep_cause; // @[playground/src/noop/cpu.scala 96:29]
  wire [63:0] fetch_io_va2pa_tlb_excep_tval; // @[playground/src/noop/cpu.scala 96:29]
  wire  fetch_io_va2pa_tlb_excep_en; // @[playground/src/noop/cpu.scala 96:29]
  wire [63:0] fetch_io_reg2if_seq_pc; // @[playground/src/noop/cpu.scala 96:29]
  wire  fetch_io_reg2if_valid; // @[playground/src/noop/cpu.scala 96:29]
  wire [63:0] fetch_io_wb2if_seq_pc; // @[playground/src/noop/cpu.scala 96:29]
  wire  fetch_io_wb2if_valid; // @[playground/src/noop/cpu.scala 96:29]
  wire  fetch_io_recov; // @[playground/src/noop/cpu.scala 96:29]
  wire  fetch_io_intr_in_en; // @[playground/src/noop/cpu.scala 96:29]
  wire [63:0] fetch_io_intr_in_cause; // @[playground/src/noop/cpu.scala 96:29]
  wire [63:0] fetch_io_branchFail_seq_pc; // @[playground/src/noop/cpu.scala 96:29]
  wire  fetch_io_branchFail_valid; // @[playground/src/noop/cpu.scala 96:29]
  wire [31:0] fetch_io_if2id_inst; // @[playground/src/noop/cpu.scala 96:29]
  wire [63:0] fetch_io_if2id_pc; // @[playground/src/noop/cpu.scala 96:29]
  wire [63:0] fetch_io_if2id_excep_cause; // @[playground/src/noop/cpu.scala 96:29]
  wire [63:0] fetch_io_if2id_excep_tval; // @[playground/src/noop/cpu.scala 96:29]
  wire  fetch_io_if2id_excep_en; // @[playground/src/noop/cpu.scala 96:29]
  wire [63:0] fetch_io_if2id_excep_pc; // @[playground/src/noop/cpu.scala 96:29]
  wire  fetch_io_if2id_drop; // @[playground/src/noop/cpu.scala 96:29]
  wire  fetch_io_if2id_stall; // @[playground/src/noop/cpu.scala 96:29]
  wire  fetch_io_if2id_recov; // @[playground/src/noop/cpu.scala 96:29]
  wire  fetch_io_if2id_valid; // @[playground/src/noop/cpu.scala 96:29]
  wire  fetch_io_if2id_ready; // @[playground/src/noop/cpu.scala 96:29]
  wire  decode_clock; // @[playground/src/noop/cpu.scala 97:29]
  wire  decode_reset; // @[playground/src/noop/cpu.scala 97:29]
  wire [31:0] decode_io_if2id_inst; // @[playground/src/noop/cpu.scala 97:29]
  wire [63:0] decode_io_if2id_pc; // @[playground/src/noop/cpu.scala 97:29]
  wire [63:0] decode_io_if2id_excep_cause; // @[playground/src/noop/cpu.scala 97:29]
  wire [63:0] decode_io_if2id_excep_tval; // @[playground/src/noop/cpu.scala 97:29]
  wire  decode_io_if2id_excep_en; // @[playground/src/noop/cpu.scala 97:29]
  wire [63:0] decode_io_if2id_excep_pc; // @[playground/src/noop/cpu.scala 97:29]
  wire  decode_io_if2id_drop; // @[playground/src/noop/cpu.scala 97:29]
  wire  decode_io_if2id_stall; // @[playground/src/noop/cpu.scala 97:29]
  wire  decode_io_if2id_recov; // @[playground/src/noop/cpu.scala 97:29]
  wire  decode_io_if2id_valid; // @[playground/src/noop/cpu.scala 97:29]
  wire  decode_io_if2id_ready; // @[playground/src/noop/cpu.scala 97:29]
  wire [31:0] decode_io_id2df_inst; // @[playground/src/noop/cpu.scala 97:29]
  wire [63:0] decode_io_id2df_pc; // @[playground/src/noop/cpu.scala 97:29]
  wire [63:0] decode_io_id2df_excep_cause; // @[playground/src/noop/cpu.scala 97:29]
  wire [63:0] decode_io_id2df_excep_tval; // @[playground/src/noop/cpu.scala 97:29]
  wire  decode_io_id2df_excep_en; // @[playground/src/noop/cpu.scala 97:29]
  wire [63:0] decode_io_id2df_excep_pc; // @[playground/src/noop/cpu.scala 97:29]
  wire [1:0] decode_io_id2df_excep_etype; // @[playground/src/noop/cpu.scala 97:29]
  wire [4:0] decode_io_id2df_ctrl_aluOp; // @[playground/src/noop/cpu.scala 97:29]
  wire  decode_io_id2df_ctrl_aluWidth; // @[playground/src/noop/cpu.scala 97:29]
  wire [4:0] decode_io_id2df_ctrl_dcMode; // @[playground/src/noop/cpu.scala 97:29]
  wire  decode_io_id2df_ctrl_writeRegEn; // @[playground/src/noop/cpu.scala 97:29]
  wire  decode_io_id2df_ctrl_writeCSREn; // @[playground/src/noop/cpu.scala 97:29]
  wire [2:0] decode_io_id2df_ctrl_brType; // @[playground/src/noop/cpu.scala 97:29]
  wire [4:0] decode_io_id2df_rs1; // @[playground/src/noop/cpu.scala 97:29]
  wire  decode_io_id2df_rrs1; // @[playground/src/noop/cpu.scala 97:29]
  wire [63:0] decode_io_id2df_rs1_d; // @[playground/src/noop/cpu.scala 97:29]
  wire [11:0] decode_io_id2df_rs2; // @[playground/src/noop/cpu.scala 97:29]
  wire  decode_io_id2df_rrs2; // @[playground/src/noop/cpu.scala 97:29]
  wire [63:0] decode_io_id2df_rs2_d; // @[playground/src/noop/cpu.scala 97:29]
  wire [4:0] decode_io_id2df_dst; // @[playground/src/noop/cpu.scala 97:29]
  wire [63:0] decode_io_id2df_dst_d; // @[playground/src/noop/cpu.scala 97:29]
  wire [1:0] decode_io_id2df_jmp_type; // @[playground/src/noop/cpu.scala 97:29]
  wire [1:0] decode_io_id2df_special; // @[playground/src/noop/cpu.scala 97:29]
  wire [5:0] decode_io_id2df_swap; // @[playground/src/noop/cpu.scala 97:29]
  wire [1:0] decode_io_id2df_indi; // @[playground/src/noop/cpu.scala 97:29]
  wire  decode_io_id2df_drop; // @[playground/src/noop/cpu.scala 97:29]
  wire  decode_io_id2df_stall; // @[playground/src/noop/cpu.scala 97:29]
  wire  decode_io_id2df_recov; // @[playground/src/noop/cpu.scala 97:29]
  wire  decode_io_id2df_valid; // @[playground/src/noop/cpu.scala 97:29]
  wire  decode_io_id2df_ready; // @[playground/src/noop/cpu.scala 97:29]
  wire [1:0] decode_io_idState_priv; // @[playground/src/noop/cpu.scala 97:29]
  wire  forwading_clock; // @[playground/src/noop/cpu.scala 98:29]
  wire  forwading_reset; // @[playground/src/noop/cpu.scala 98:29]
  wire [31:0] forwading_io_id2df_inst; // @[playground/src/noop/cpu.scala 98:29]
  wire [63:0] forwading_io_id2df_pc; // @[playground/src/noop/cpu.scala 98:29]
  wire [63:0] forwading_io_id2df_excep_cause; // @[playground/src/noop/cpu.scala 98:29]
  wire [63:0] forwading_io_id2df_excep_tval; // @[playground/src/noop/cpu.scala 98:29]
  wire  forwading_io_id2df_excep_en; // @[playground/src/noop/cpu.scala 98:29]
  wire [63:0] forwading_io_id2df_excep_pc; // @[playground/src/noop/cpu.scala 98:29]
  wire [1:0] forwading_io_id2df_excep_etype; // @[playground/src/noop/cpu.scala 98:29]
  wire [4:0] forwading_io_id2df_ctrl_aluOp; // @[playground/src/noop/cpu.scala 98:29]
  wire  forwading_io_id2df_ctrl_aluWidth; // @[playground/src/noop/cpu.scala 98:29]
  wire [4:0] forwading_io_id2df_ctrl_dcMode; // @[playground/src/noop/cpu.scala 98:29]
  wire  forwading_io_id2df_ctrl_writeRegEn; // @[playground/src/noop/cpu.scala 98:29]
  wire  forwading_io_id2df_ctrl_writeCSREn; // @[playground/src/noop/cpu.scala 98:29]
  wire [2:0] forwading_io_id2df_ctrl_brType; // @[playground/src/noop/cpu.scala 98:29]
  wire [4:0] forwading_io_id2df_rs1; // @[playground/src/noop/cpu.scala 98:29]
  wire  forwading_io_id2df_rrs1; // @[playground/src/noop/cpu.scala 98:29]
  wire [63:0] forwading_io_id2df_rs1_d; // @[playground/src/noop/cpu.scala 98:29]
  wire [11:0] forwading_io_id2df_rs2; // @[playground/src/noop/cpu.scala 98:29]
  wire  forwading_io_id2df_rrs2; // @[playground/src/noop/cpu.scala 98:29]
  wire [63:0] forwading_io_id2df_rs2_d; // @[playground/src/noop/cpu.scala 98:29]
  wire [4:0] forwading_io_id2df_dst; // @[playground/src/noop/cpu.scala 98:29]
  wire [63:0] forwading_io_id2df_dst_d; // @[playground/src/noop/cpu.scala 98:29]
  wire [1:0] forwading_io_id2df_jmp_type; // @[playground/src/noop/cpu.scala 98:29]
  wire [1:0] forwading_io_id2df_special; // @[playground/src/noop/cpu.scala 98:29]
  wire [5:0] forwading_io_id2df_swap; // @[playground/src/noop/cpu.scala 98:29]
  wire [1:0] forwading_io_id2df_indi; // @[playground/src/noop/cpu.scala 98:29]
  wire  forwading_io_id2df_drop; // @[playground/src/noop/cpu.scala 98:29]
  wire  forwading_io_id2df_stall; // @[playground/src/noop/cpu.scala 98:29]
  wire  forwading_io_id2df_recov; // @[playground/src/noop/cpu.scala 98:29]
  wire  forwading_io_id2df_valid; // @[playground/src/noop/cpu.scala 98:29]
  wire  forwading_io_id2df_ready; // @[playground/src/noop/cpu.scala 98:29]
  wire [31:0] forwading_io_df2rr_inst; // @[playground/src/noop/cpu.scala 98:29]
  wire [63:0] forwading_io_df2rr_pc; // @[playground/src/noop/cpu.scala 98:29]
  wire [63:0] forwading_io_df2rr_excep_cause; // @[playground/src/noop/cpu.scala 98:29]
  wire [63:0] forwading_io_df2rr_excep_tval; // @[playground/src/noop/cpu.scala 98:29]
  wire  forwading_io_df2rr_excep_en; // @[playground/src/noop/cpu.scala 98:29]
  wire [63:0] forwading_io_df2rr_excep_pc; // @[playground/src/noop/cpu.scala 98:29]
  wire [1:0] forwading_io_df2rr_excep_etype; // @[playground/src/noop/cpu.scala 98:29]
  wire [4:0] forwading_io_df2rr_ctrl_aluOp; // @[playground/src/noop/cpu.scala 98:29]
  wire  forwading_io_df2rr_ctrl_aluWidth; // @[playground/src/noop/cpu.scala 98:29]
  wire [4:0] forwading_io_df2rr_ctrl_dcMode; // @[playground/src/noop/cpu.scala 98:29]
  wire  forwading_io_df2rr_ctrl_writeRegEn; // @[playground/src/noop/cpu.scala 98:29]
  wire  forwading_io_df2rr_ctrl_writeCSREn; // @[playground/src/noop/cpu.scala 98:29]
  wire [2:0] forwading_io_df2rr_ctrl_brType; // @[playground/src/noop/cpu.scala 98:29]
  wire [4:0] forwading_io_df2rr_rs1; // @[playground/src/noop/cpu.scala 98:29]
  wire  forwading_io_df2rr_rrs1; // @[playground/src/noop/cpu.scala 98:29]
  wire [63:0] forwading_io_df2rr_rs1_d; // @[playground/src/noop/cpu.scala 98:29]
  wire [11:0] forwading_io_df2rr_rs2; // @[playground/src/noop/cpu.scala 98:29]
  wire  forwading_io_df2rr_rrs2; // @[playground/src/noop/cpu.scala 98:29]
  wire [63:0] forwading_io_df2rr_rs2_d; // @[playground/src/noop/cpu.scala 98:29]
  wire [4:0] forwading_io_df2rr_dst; // @[playground/src/noop/cpu.scala 98:29]
  wire [63:0] forwading_io_df2rr_dst_d; // @[playground/src/noop/cpu.scala 98:29]
  wire [1:0] forwading_io_df2rr_jmp_type; // @[playground/src/noop/cpu.scala 98:29]
  wire [1:0] forwading_io_df2rr_special; // @[playground/src/noop/cpu.scala 98:29]
  wire [5:0] forwading_io_df2rr_swap; // @[playground/src/noop/cpu.scala 98:29]
  wire [1:0] forwading_io_df2rr_indi; // @[playground/src/noop/cpu.scala 98:29]
  wire  forwading_io_df2rr_drop; // @[playground/src/noop/cpu.scala 98:29]
  wire  forwading_io_df2rr_stall; // @[playground/src/noop/cpu.scala 98:29]
  wire  forwading_io_df2rr_recov; // @[playground/src/noop/cpu.scala 98:29]
  wire  forwading_io_df2rr_valid; // @[playground/src/noop/cpu.scala 98:29]
  wire  forwading_io_df2rr_ready; // @[playground/src/noop/cpu.scala 98:29]
  wire [4:0] forwading_io_d_rr_id; // @[playground/src/noop/cpu.scala 98:29]
  wire [63:0] forwading_io_d_rr_data; // @[playground/src/noop/cpu.scala 98:29]
  wire [1:0] forwading_io_d_rr_state; // @[playground/src/noop/cpu.scala 98:29]
  wire [4:0] forwading_io_d_ex_id; // @[playground/src/noop/cpu.scala 98:29]
  wire [63:0] forwading_io_d_ex_data; // @[playground/src/noop/cpu.scala 98:29]
  wire [1:0] forwading_io_d_ex_state; // @[playground/src/noop/cpu.scala 98:29]
  wire [4:0] forwading_io_d_mem1_id; // @[playground/src/noop/cpu.scala 98:29]
  wire [63:0] forwading_io_d_mem1_data; // @[playground/src/noop/cpu.scala 98:29]
  wire [1:0] forwading_io_d_mem1_state; // @[playground/src/noop/cpu.scala 98:29]
  wire [4:0] forwading_io_d_mem2_id; // @[playground/src/noop/cpu.scala 98:29]
  wire [63:0] forwading_io_d_mem2_data; // @[playground/src/noop/cpu.scala 98:29]
  wire [1:0] forwading_io_d_mem2_state; // @[playground/src/noop/cpu.scala 98:29]
  wire [4:0] forwading_io_d_mem3_id; // @[playground/src/noop/cpu.scala 98:29]
  wire [63:0] forwading_io_d_mem3_data; // @[playground/src/noop/cpu.scala 98:29]
  wire [1:0] forwading_io_d_mem3_state; // @[playground/src/noop/cpu.scala 98:29]
  wire  readregs_clock; // @[playground/src/noop/cpu.scala 99:29]
  wire  readregs_reset; // @[playground/src/noop/cpu.scala 99:29]
  wire [31:0] readregs_io_df2rr_inst; // @[playground/src/noop/cpu.scala 99:29]
  wire [63:0] readregs_io_df2rr_pc; // @[playground/src/noop/cpu.scala 99:29]
  wire [63:0] readregs_io_df2rr_excep_cause; // @[playground/src/noop/cpu.scala 99:29]
  wire [63:0] readregs_io_df2rr_excep_tval; // @[playground/src/noop/cpu.scala 99:29]
  wire  readregs_io_df2rr_excep_en; // @[playground/src/noop/cpu.scala 99:29]
  wire [63:0] readregs_io_df2rr_excep_pc; // @[playground/src/noop/cpu.scala 99:29]
  wire [1:0] readregs_io_df2rr_excep_etype; // @[playground/src/noop/cpu.scala 99:29]
  wire [4:0] readregs_io_df2rr_ctrl_aluOp; // @[playground/src/noop/cpu.scala 99:29]
  wire  readregs_io_df2rr_ctrl_aluWidth; // @[playground/src/noop/cpu.scala 99:29]
  wire [4:0] readregs_io_df2rr_ctrl_dcMode; // @[playground/src/noop/cpu.scala 99:29]
  wire  readregs_io_df2rr_ctrl_writeRegEn; // @[playground/src/noop/cpu.scala 99:29]
  wire  readregs_io_df2rr_ctrl_writeCSREn; // @[playground/src/noop/cpu.scala 99:29]
  wire [2:0] readregs_io_df2rr_ctrl_brType; // @[playground/src/noop/cpu.scala 99:29]
  wire [4:0] readregs_io_df2rr_rs1; // @[playground/src/noop/cpu.scala 99:29]
  wire  readregs_io_df2rr_rrs1; // @[playground/src/noop/cpu.scala 99:29]
  wire [63:0] readregs_io_df2rr_rs1_d; // @[playground/src/noop/cpu.scala 99:29]
  wire [11:0] readregs_io_df2rr_rs2; // @[playground/src/noop/cpu.scala 99:29]
  wire  readregs_io_df2rr_rrs2; // @[playground/src/noop/cpu.scala 99:29]
  wire [63:0] readregs_io_df2rr_rs2_d; // @[playground/src/noop/cpu.scala 99:29]
  wire [4:0] readregs_io_df2rr_dst; // @[playground/src/noop/cpu.scala 99:29]
  wire [63:0] readregs_io_df2rr_dst_d; // @[playground/src/noop/cpu.scala 99:29]
  wire [1:0] readregs_io_df2rr_jmp_type; // @[playground/src/noop/cpu.scala 99:29]
  wire [1:0] readregs_io_df2rr_special; // @[playground/src/noop/cpu.scala 99:29]
  wire [5:0] readregs_io_df2rr_swap; // @[playground/src/noop/cpu.scala 99:29]
  wire [1:0] readregs_io_df2rr_indi; // @[playground/src/noop/cpu.scala 99:29]
  wire  readregs_io_df2rr_drop; // @[playground/src/noop/cpu.scala 99:29]
  wire  readregs_io_df2rr_stall; // @[playground/src/noop/cpu.scala 99:29]
  wire  readregs_io_df2rr_recov; // @[playground/src/noop/cpu.scala 99:29]
  wire  readregs_io_df2rr_valid; // @[playground/src/noop/cpu.scala 99:29]
  wire  readregs_io_df2rr_ready; // @[playground/src/noop/cpu.scala 99:29]
  wire [31:0] readregs_io_rr2ex_inst; // @[playground/src/noop/cpu.scala 99:29]
  wire [63:0] readregs_io_rr2ex_pc; // @[playground/src/noop/cpu.scala 99:29]
  wire [63:0] readregs_io_rr2ex_excep_cause; // @[playground/src/noop/cpu.scala 99:29]
  wire [63:0] readregs_io_rr2ex_excep_tval; // @[playground/src/noop/cpu.scala 99:29]
  wire  readregs_io_rr2ex_excep_en; // @[playground/src/noop/cpu.scala 99:29]
  wire [63:0] readregs_io_rr2ex_excep_pc; // @[playground/src/noop/cpu.scala 99:29]
  wire [1:0] readregs_io_rr2ex_excep_etype; // @[playground/src/noop/cpu.scala 99:29]
  wire [4:0] readregs_io_rr2ex_ctrl_aluOp; // @[playground/src/noop/cpu.scala 99:29]
  wire  readregs_io_rr2ex_ctrl_aluWidth; // @[playground/src/noop/cpu.scala 99:29]
  wire [4:0] readregs_io_rr2ex_ctrl_dcMode; // @[playground/src/noop/cpu.scala 99:29]
  wire  readregs_io_rr2ex_ctrl_writeRegEn; // @[playground/src/noop/cpu.scala 99:29]
  wire  readregs_io_rr2ex_ctrl_writeCSREn; // @[playground/src/noop/cpu.scala 99:29]
  wire [2:0] readregs_io_rr2ex_ctrl_brType; // @[playground/src/noop/cpu.scala 99:29]
  wire [63:0] readregs_io_rr2ex_rs1_d; // @[playground/src/noop/cpu.scala 99:29]
  wire [11:0] readregs_io_rr2ex_rs2; // @[playground/src/noop/cpu.scala 99:29]
  wire [63:0] readregs_io_rr2ex_rs2_d; // @[playground/src/noop/cpu.scala 99:29]
  wire [4:0] readregs_io_rr2ex_dst; // @[playground/src/noop/cpu.scala 99:29]
  wire [63:0] readregs_io_rr2ex_dst_d; // @[playground/src/noop/cpu.scala 99:29]
  wire [11:0] readregs_io_rr2ex_rcsr_id; // @[playground/src/noop/cpu.scala 99:29]
  wire [1:0] readregs_io_rr2ex_jmp_type; // @[playground/src/noop/cpu.scala 99:29]
  wire [1:0] readregs_io_rr2ex_special; // @[playground/src/noop/cpu.scala 99:29]
  wire [1:0] readregs_io_rr2ex_indi; // @[playground/src/noop/cpu.scala 99:29]
  wire  readregs_io_rr2ex_drop; // @[playground/src/noop/cpu.scala 99:29]
  wire  readregs_io_rr2ex_stall; // @[playground/src/noop/cpu.scala 99:29]
  wire  readregs_io_rr2ex_recov; // @[playground/src/noop/cpu.scala 99:29]
  wire  readregs_io_rr2ex_valid; // @[playground/src/noop/cpu.scala 99:29]
  wire  readregs_io_rr2ex_ready; // @[playground/src/noop/cpu.scala 99:29]
  wire [4:0] readregs_io_rs1Read_id; // @[playground/src/noop/cpu.scala 99:29]
  wire [63:0] readregs_io_rs1Read_data; // @[playground/src/noop/cpu.scala 99:29]
  wire [4:0] readregs_io_rs2Read_id; // @[playground/src/noop/cpu.scala 99:29]
  wire [63:0] readregs_io_rs2Read_data; // @[playground/src/noop/cpu.scala 99:29]
  wire [11:0] readregs_io_csrRead_id; // @[playground/src/noop/cpu.scala 99:29]
  wire [63:0] readregs_io_csrRead_data; // @[playground/src/noop/cpu.scala 99:29]
  wire  readregs_io_csrRead_is_err; // @[playground/src/noop/cpu.scala 99:29]
  wire [4:0] readregs_io_d_rr_id; // @[playground/src/noop/cpu.scala 99:29]
  wire [63:0] readregs_io_d_rr_data; // @[playground/src/noop/cpu.scala 99:29]
  wire [1:0] readregs_io_d_rr_state; // @[playground/src/noop/cpu.scala 99:29]
  wire  execute_clock; // @[playground/src/noop/cpu.scala 100:29]
  wire  execute_reset; // @[playground/src/noop/cpu.scala 100:29]
  wire [31:0] execute_io_rr2ex_inst; // @[playground/src/noop/cpu.scala 100:29]
  wire [63:0] execute_io_rr2ex_pc; // @[playground/src/noop/cpu.scala 100:29]
  wire [63:0] execute_io_rr2ex_excep_cause; // @[playground/src/noop/cpu.scala 100:29]
  wire [63:0] execute_io_rr2ex_excep_tval; // @[playground/src/noop/cpu.scala 100:29]
  wire  execute_io_rr2ex_excep_en; // @[playground/src/noop/cpu.scala 100:29]
  wire [63:0] execute_io_rr2ex_excep_pc; // @[playground/src/noop/cpu.scala 100:29]
  wire [1:0] execute_io_rr2ex_excep_etype; // @[playground/src/noop/cpu.scala 100:29]
  wire [4:0] execute_io_rr2ex_ctrl_aluOp; // @[playground/src/noop/cpu.scala 100:29]
  wire  execute_io_rr2ex_ctrl_aluWidth; // @[playground/src/noop/cpu.scala 100:29]
  wire [4:0] execute_io_rr2ex_ctrl_dcMode; // @[playground/src/noop/cpu.scala 100:29]
  wire  execute_io_rr2ex_ctrl_writeRegEn; // @[playground/src/noop/cpu.scala 100:29]
  wire  execute_io_rr2ex_ctrl_writeCSREn; // @[playground/src/noop/cpu.scala 100:29]
  wire [2:0] execute_io_rr2ex_ctrl_brType; // @[playground/src/noop/cpu.scala 100:29]
  wire [63:0] execute_io_rr2ex_rs1_d; // @[playground/src/noop/cpu.scala 100:29]
  wire [11:0] execute_io_rr2ex_rs2; // @[playground/src/noop/cpu.scala 100:29]
  wire [63:0] execute_io_rr2ex_rs2_d; // @[playground/src/noop/cpu.scala 100:29]
  wire [4:0] execute_io_rr2ex_dst; // @[playground/src/noop/cpu.scala 100:29]
  wire [63:0] execute_io_rr2ex_dst_d; // @[playground/src/noop/cpu.scala 100:29]
  wire [11:0] execute_io_rr2ex_rcsr_id; // @[playground/src/noop/cpu.scala 100:29]
  wire [1:0] execute_io_rr2ex_jmp_type; // @[playground/src/noop/cpu.scala 100:29]
  wire [1:0] execute_io_rr2ex_special; // @[playground/src/noop/cpu.scala 100:29]
  wire [1:0] execute_io_rr2ex_indi; // @[playground/src/noop/cpu.scala 100:29]
  wire  execute_io_rr2ex_drop; // @[playground/src/noop/cpu.scala 100:29]
  wire  execute_io_rr2ex_stall; // @[playground/src/noop/cpu.scala 100:29]
  wire  execute_io_rr2ex_recov; // @[playground/src/noop/cpu.scala 100:29]
  wire  execute_io_rr2ex_valid; // @[playground/src/noop/cpu.scala 100:29]
  wire  execute_io_rr2ex_ready; // @[playground/src/noop/cpu.scala 100:29]
  wire [31:0] execute_io_ex2mem_inst; // @[playground/src/noop/cpu.scala 100:29]
  wire [63:0] execute_io_ex2mem_pc; // @[playground/src/noop/cpu.scala 100:29]
  wire [63:0] execute_io_ex2mem_excep_cause; // @[playground/src/noop/cpu.scala 100:29]
  wire [63:0] execute_io_ex2mem_excep_tval; // @[playground/src/noop/cpu.scala 100:29]
  wire  execute_io_ex2mem_excep_en; // @[playground/src/noop/cpu.scala 100:29]
  wire [63:0] execute_io_ex2mem_excep_pc; // @[playground/src/noop/cpu.scala 100:29]
  wire [1:0] execute_io_ex2mem_excep_etype; // @[playground/src/noop/cpu.scala 100:29]
  wire [4:0] execute_io_ex2mem_ctrl_dcMode; // @[playground/src/noop/cpu.scala 100:29]
  wire  execute_io_ex2mem_ctrl_writeRegEn; // @[playground/src/noop/cpu.scala 100:29]
  wire  execute_io_ex2mem_ctrl_writeCSREn; // @[playground/src/noop/cpu.scala 100:29]
  wire [63:0] execute_io_ex2mem_mem_addr; // @[playground/src/noop/cpu.scala 100:29]
  wire [63:0] execute_io_ex2mem_mem_data; // @[playground/src/noop/cpu.scala 100:29]
  wire [11:0] execute_io_ex2mem_csr_id; // @[playground/src/noop/cpu.scala 100:29]
  wire [63:0] execute_io_ex2mem_csr_d; // @[playground/src/noop/cpu.scala 100:29]
  wire [4:0] execute_io_ex2mem_dst; // @[playground/src/noop/cpu.scala 100:29]
  wire [63:0] execute_io_ex2mem_dst_d; // @[playground/src/noop/cpu.scala 100:29]
  wire [11:0] execute_io_ex2mem_rcsr_id; // @[playground/src/noop/cpu.scala 100:29]
  wire [1:0] execute_io_ex2mem_special; // @[playground/src/noop/cpu.scala 100:29]
  wire [1:0] execute_io_ex2mem_indi; // @[playground/src/noop/cpu.scala 100:29]
  wire  execute_io_ex2mem_drop; // @[playground/src/noop/cpu.scala 100:29]
  wire  execute_io_ex2mem_stall; // @[playground/src/noop/cpu.scala 100:29]
  wire  execute_io_ex2mem_recov; // @[playground/src/noop/cpu.scala 100:29]
  wire  execute_io_ex2mem_valid; // @[playground/src/noop/cpu.scala 100:29]
  wire  execute_io_ex2mem_ready; // @[playground/src/noop/cpu.scala 100:29]
  wire [4:0] execute_io_d_ex_id; // @[playground/src/noop/cpu.scala 100:29]
  wire [63:0] execute_io_d_ex_data; // @[playground/src/noop/cpu.scala 100:29]
  wire [1:0] execute_io_d_ex_state; // @[playground/src/noop/cpu.scala 100:29]
  wire [63:0] execute_io_ex2if_seq_pc; // @[playground/src/noop/cpu.scala 100:29]
  wire  execute_io_ex2if_valid; // @[playground/src/noop/cpu.scala 100:29]
  wire [63:0] execute_io_updateNextPc_seq_pc; // @[playground/src/noop/cpu.scala 100:29]
  wire  execute_io_updateNextPc_valid; // @[playground/src/noop/cpu.scala 100:29]
  wire  memory_clock; // @[playground/src/noop/cpu.scala 101:29]
  wire  memory_reset; // @[playground/src/noop/cpu.scala 101:29]
  wire [31:0] memory_io_ex2mem_inst; // @[playground/src/noop/cpu.scala 101:29]
  wire [63:0] memory_io_ex2mem_pc; // @[playground/src/noop/cpu.scala 101:29]
  wire [63:0] memory_io_ex2mem_excep_cause; // @[playground/src/noop/cpu.scala 101:29]
  wire [63:0] memory_io_ex2mem_excep_tval; // @[playground/src/noop/cpu.scala 101:29]
  wire  memory_io_ex2mem_excep_en; // @[playground/src/noop/cpu.scala 101:29]
  wire [63:0] memory_io_ex2mem_excep_pc; // @[playground/src/noop/cpu.scala 101:29]
  wire [1:0] memory_io_ex2mem_excep_etype; // @[playground/src/noop/cpu.scala 101:29]
  wire [4:0] memory_io_ex2mem_ctrl_dcMode; // @[playground/src/noop/cpu.scala 101:29]
  wire  memory_io_ex2mem_ctrl_writeRegEn; // @[playground/src/noop/cpu.scala 101:29]
  wire  memory_io_ex2mem_ctrl_writeCSREn; // @[playground/src/noop/cpu.scala 101:29]
  wire [63:0] memory_io_ex2mem_mem_addr; // @[playground/src/noop/cpu.scala 101:29]
  wire [63:0] memory_io_ex2mem_mem_data; // @[playground/src/noop/cpu.scala 101:29]
  wire [11:0] memory_io_ex2mem_csr_id; // @[playground/src/noop/cpu.scala 101:29]
  wire [63:0] memory_io_ex2mem_csr_d; // @[playground/src/noop/cpu.scala 101:29]
  wire [4:0] memory_io_ex2mem_dst; // @[playground/src/noop/cpu.scala 101:29]
  wire [63:0] memory_io_ex2mem_dst_d; // @[playground/src/noop/cpu.scala 101:29]
  wire [11:0] memory_io_ex2mem_rcsr_id; // @[playground/src/noop/cpu.scala 101:29]
  wire [1:0] memory_io_ex2mem_special; // @[playground/src/noop/cpu.scala 101:29]
  wire [1:0] memory_io_ex2mem_indi; // @[playground/src/noop/cpu.scala 101:29]
  wire  memory_io_ex2mem_drop; // @[playground/src/noop/cpu.scala 101:29]
  wire  memory_io_ex2mem_stall; // @[playground/src/noop/cpu.scala 101:29]
  wire  memory_io_ex2mem_recov; // @[playground/src/noop/cpu.scala 101:29]
  wire  memory_io_ex2mem_valid; // @[playground/src/noop/cpu.scala 101:29]
  wire  memory_io_ex2mem_ready; // @[playground/src/noop/cpu.scala 101:29]
  wire [31:0] memory_io_mem2rb_inst; // @[playground/src/noop/cpu.scala 101:29]
  wire [63:0] memory_io_mem2rb_pc; // @[playground/src/noop/cpu.scala 101:29]
  wire [63:0] memory_io_mem2rb_excep_cause; // @[playground/src/noop/cpu.scala 101:29]
  wire [63:0] memory_io_mem2rb_excep_tval; // @[playground/src/noop/cpu.scala 101:29]
  wire  memory_io_mem2rb_excep_en; // @[playground/src/noop/cpu.scala 101:29]
  wire [63:0] memory_io_mem2rb_excep_pc; // @[playground/src/noop/cpu.scala 101:29]
  wire [1:0] memory_io_mem2rb_excep_etype; // @[playground/src/noop/cpu.scala 101:29]
  wire [11:0] memory_io_mem2rb_csr_id; // @[playground/src/noop/cpu.scala 101:29]
  wire [63:0] memory_io_mem2rb_csr_d; // @[playground/src/noop/cpu.scala 101:29]
  wire  memory_io_mem2rb_csr_en; // @[playground/src/noop/cpu.scala 101:29]
  wire [4:0] memory_io_mem2rb_dst; // @[playground/src/noop/cpu.scala 101:29]
  wire [63:0] memory_io_mem2rb_dst_d; // @[playground/src/noop/cpu.scala 101:29]
  wire  memory_io_mem2rb_dst_en; // @[playground/src/noop/cpu.scala 101:29]
  wire [11:0] memory_io_mem2rb_rcsr_id; // @[playground/src/noop/cpu.scala 101:29]
  wire [1:0] memory_io_mem2rb_special; // @[playground/src/noop/cpu.scala 101:29]
  wire  memory_io_mem2rb_is_mmio; // @[playground/src/noop/cpu.scala 101:29]
  wire  memory_io_mem2rb_drop; // @[playground/src/noop/cpu.scala 101:29]
  wire  memory_io_mem2rb_stall; // @[playground/src/noop/cpu.scala 101:29]
  wire  memory_io_mem2rb_recov; // @[playground/src/noop/cpu.scala 101:29]
  wire  memory_io_mem2rb_valid; // @[playground/src/noop/cpu.scala 101:29]
  wire  memory_io_mem2rb_ready; // @[playground/src/noop/cpu.scala 101:29]
  wire [31:0] memory_io_dataRW_addr; // @[playground/src/noop/cpu.scala 101:29]
  wire [63:0] memory_io_dataRW_rdata; // @[playground/src/noop/cpu.scala 101:29]
  wire  memory_io_dataRW_rvalid; // @[playground/src/noop/cpu.scala 101:29]
  wire [63:0] memory_io_dataRW_wdata; // @[playground/src/noop/cpu.scala 101:29]
  wire [4:0] memory_io_dataRW_dc_mode; // @[playground/src/noop/cpu.scala 101:29]
  wire [4:0] memory_io_dataRW_amo; // @[playground/src/noop/cpu.scala 101:29]
  wire  memory_io_dataRW_ready; // @[playground/src/noop/cpu.scala 101:29]
  wire [63:0] memory_io_va2pa_vaddr; // @[playground/src/noop/cpu.scala 101:29]
  wire  memory_io_va2pa_vvalid; // @[playground/src/noop/cpu.scala 101:29]
  wire [1:0] memory_io_va2pa_m_type; // @[playground/src/noop/cpu.scala 101:29]
  wire [31:0] memory_io_va2pa_paddr; // @[playground/src/noop/cpu.scala 101:29]
  wire  memory_io_va2pa_pvalid; // @[playground/src/noop/cpu.scala 101:29]
  wire [63:0] memory_io_va2pa_tlb_excep_cause; // @[playground/src/noop/cpu.scala 101:29]
  wire [63:0] memory_io_va2pa_tlb_excep_tval; // @[playground/src/noop/cpu.scala 101:29]
  wire  memory_io_va2pa_tlb_excep_en; // @[playground/src/noop/cpu.scala 101:29]
  wire [4:0] memory_io_d_mem1_id; // @[playground/src/noop/cpu.scala 101:29]
  wire [63:0] memory_io_d_mem1_data; // @[playground/src/noop/cpu.scala 101:29]
  wire [1:0] memory_io_d_mem1_state; // @[playground/src/noop/cpu.scala 101:29]
  wire [4:0] memory_io_d_mem2_id; // @[playground/src/noop/cpu.scala 101:29]
  wire [63:0] memory_io_d_mem2_data; // @[playground/src/noop/cpu.scala 101:29]
  wire [1:0] memory_io_d_mem2_state; // @[playground/src/noop/cpu.scala 101:29]
  wire [4:0] memory_io_d_mem3_id; // @[playground/src/noop/cpu.scala 101:29]
  wire [63:0] memory_io_d_mem3_data; // @[playground/src/noop/cpu.scala 101:29]
  wire [1:0] memory_io_d_mem3_state; // @[playground/src/noop/cpu.scala 101:29]
  wire  writeback_clock; // @[playground/src/noop/cpu.scala 102:29]
  wire  writeback_reset; // @[playground/src/noop/cpu.scala 102:29]
  wire [31:0] writeback_io_mem2rb_inst; // @[playground/src/noop/cpu.scala 102:29]
  wire [63:0] writeback_io_mem2rb_pc; // @[playground/src/noop/cpu.scala 102:29]
  wire [63:0] writeback_io_mem2rb_excep_cause; // @[playground/src/noop/cpu.scala 102:29]
  wire [63:0] writeback_io_mem2rb_excep_tval; // @[playground/src/noop/cpu.scala 102:29]
  wire  writeback_io_mem2rb_excep_en; // @[playground/src/noop/cpu.scala 102:29]
  wire [63:0] writeback_io_mem2rb_excep_pc; // @[playground/src/noop/cpu.scala 102:29]
  wire [1:0] writeback_io_mem2rb_excep_etype; // @[playground/src/noop/cpu.scala 102:29]
  wire [11:0] writeback_io_mem2rb_csr_id; // @[playground/src/noop/cpu.scala 102:29]
  wire [63:0] writeback_io_mem2rb_csr_d; // @[playground/src/noop/cpu.scala 102:29]
  wire  writeback_io_mem2rb_csr_en; // @[playground/src/noop/cpu.scala 102:29]
  wire [4:0] writeback_io_mem2rb_dst; // @[playground/src/noop/cpu.scala 102:29]
  wire [63:0] writeback_io_mem2rb_dst_d; // @[playground/src/noop/cpu.scala 102:29]
  wire  writeback_io_mem2rb_dst_en; // @[playground/src/noop/cpu.scala 102:29]
  wire [11:0] writeback_io_mem2rb_rcsr_id; // @[playground/src/noop/cpu.scala 102:29]
  wire [1:0] writeback_io_mem2rb_special; // @[playground/src/noop/cpu.scala 102:29]
  wire  writeback_io_mem2rb_is_mmio; // @[playground/src/noop/cpu.scala 102:29]
  wire  writeback_io_mem2rb_drop; // @[playground/src/noop/cpu.scala 102:29]
  wire  writeback_io_mem2rb_stall; // @[playground/src/noop/cpu.scala 102:29]
  wire  writeback_io_mem2rb_recov; // @[playground/src/noop/cpu.scala 102:29]
  wire  writeback_io_mem2rb_valid; // @[playground/src/noop/cpu.scala 102:29]
  wire  writeback_io_mem2rb_ready; // @[playground/src/noop/cpu.scala 102:29]
  wire [4:0] writeback_io_wReg_id; // @[playground/src/noop/cpu.scala 102:29]
  wire [63:0] writeback_io_wReg_data; // @[playground/src/noop/cpu.scala 102:29]
  wire  writeback_io_wReg_en; // @[playground/src/noop/cpu.scala 102:29]
  wire [11:0] writeback_io_wCsr_id; // @[playground/src/noop/cpu.scala 102:29]
  wire [63:0] writeback_io_wCsr_data; // @[playground/src/noop/cpu.scala 102:29]
  wire  writeback_io_wCsr_en; // @[playground/src/noop/cpu.scala 102:29]
  wire [63:0] writeback_io_excep_cause; // @[playground/src/noop/cpu.scala 102:29]
  wire [63:0] writeback_io_excep_tval; // @[playground/src/noop/cpu.scala 102:29]
  wire  writeback_io_excep_en; // @[playground/src/noop/cpu.scala 102:29]
  wire [63:0] writeback_io_excep_pc; // @[playground/src/noop/cpu.scala 102:29]
  wire [1:0] writeback_io_excep_etype; // @[playground/src/noop/cpu.scala 102:29]
  wire [63:0] writeback_io_wb2if_seq_pc; // @[playground/src/noop/cpu.scala 102:29]
  wire  writeback_io_wb2if_valid; // @[playground/src/noop/cpu.scala 102:29]
  wire  writeback_io_recov; // @[playground/src/noop/cpu.scala 102:29]
  wire  writeback_io_flush_tlb; // @[playground/src/noop/cpu.scala 102:29]
  wire  writeback_io_flush_cache; // @[playground/src/noop/cpu.scala 102:29]
  wire  regs_clock; // @[playground/src/noop/cpu.scala 104:29]
  wire  regs_reset; // @[playground/src/noop/cpu.scala 104:29]
  wire [4:0] regs_io_rs1_id; // @[playground/src/noop/cpu.scala 104:29]
  wire [63:0] regs_io_rs1_data; // @[playground/src/noop/cpu.scala 104:29]
  wire [4:0] regs_io_rs2_id; // @[playground/src/noop/cpu.scala 104:29]
  wire [63:0] regs_io_rs2_data; // @[playground/src/noop/cpu.scala 104:29]
  wire [4:0] regs_io_dst_id; // @[playground/src/noop/cpu.scala 104:29]
  wire [63:0] regs_io_dst_data; // @[playground/src/noop/cpu.scala 104:29]
  wire  regs_io_dst_en; // @[playground/src/noop/cpu.scala 104:29]
  wire  csrs_clock; // @[playground/src/noop/cpu.scala 105:29]
  wire  csrs_reset; // @[playground/src/noop/cpu.scala 105:29]
  wire [11:0] csrs_io_rs_id; // @[playground/src/noop/cpu.scala 105:29]
  wire [63:0] csrs_io_rs_data; // @[playground/src/noop/cpu.scala 105:29]
  wire  csrs_io_rs_is_err; // @[playground/src/noop/cpu.scala 105:29]
  wire [11:0] csrs_io_rd_id; // @[playground/src/noop/cpu.scala 105:29]
  wire [63:0] csrs_io_rd_data; // @[playground/src/noop/cpu.scala 105:29]
  wire  csrs_io_rd_en; // @[playground/src/noop/cpu.scala 105:29]
  wire [63:0] csrs_io_excep_cause; // @[playground/src/noop/cpu.scala 105:29]
  wire [63:0] csrs_io_excep_tval; // @[playground/src/noop/cpu.scala 105:29]
  wire  csrs_io_excep_en; // @[playground/src/noop/cpu.scala 105:29]
  wire [63:0] csrs_io_excep_pc; // @[playground/src/noop/cpu.scala 105:29]
  wire [1:0] csrs_io_excep_etype; // @[playground/src/noop/cpu.scala 105:29]
  wire [1:0] csrs_io_mmuState_priv; // @[playground/src/noop/cpu.scala 105:29]
  wire [63:0] csrs_io_mmuState_mstatus; // @[playground/src/noop/cpu.scala 105:29]
  wire [63:0] csrs_io_mmuState_satp; // @[playground/src/noop/cpu.scala 105:29]
  wire [1:0] csrs_io_idState_priv; // @[playground/src/noop/cpu.scala 105:29]
  wire [63:0] csrs_io_reg2if_seq_pc; // @[playground/src/noop/cpu.scala 105:29]
  wire  csrs_io_reg2if_valid; // @[playground/src/noop/cpu.scala 105:29]
  wire  csrs_io_intr_out_en; // @[playground/src/noop/cpu.scala 105:29]
  wire [63:0] csrs_io_intr_out_cause; // @[playground/src/noop/cpu.scala 105:29]
  wire  csrs_io_clint_raise; // @[playground/src/noop/cpu.scala 105:29]
  wire  csrs_io_clint_clear; // @[playground/src/noop/cpu.scala 105:29]
  wire  csrs_io_plic_m_raise; // @[playground/src/noop/cpu.scala 105:29]
  wire  csrs_io_plic_m_clear; // @[playground/src/noop/cpu.scala 105:29]
  wire  csrs_io_plic_s_raise; // @[playground/src/noop/cpu.scala 105:29]
  wire  csrs_io_plic_s_clear; // @[playground/src/noop/cpu.scala 105:29]
  wire [63:0] csrs_io_updateNextPc_seq_pc; // @[playground/src/noop/cpu.scala 105:29]
  wire  csrs_io_updateNextPc_valid; // @[playground/src/noop/cpu.scala 105:29]
  wire  csrs_io_intr_msip_raise; // @[playground/src/noop/cpu.scala 105:29]
  wire  csrs_io_intr_msip_clear; // @[playground/src/noop/cpu.scala 105:29]
  wire  icache_clock; // @[playground/src/noop/cpu.scala 106:29]
  wire  icache_reset; // @[playground/src/noop/cpu.scala 106:29]
  wire  icache_io_instAxi_ra_ready; // @[playground/src/noop/cpu.scala 106:29]
  wire  icache_io_instAxi_ra_valid; // @[playground/src/noop/cpu.scala 106:29]
  wire [31:0] icache_io_instAxi_ra_bits_addr; // @[playground/src/noop/cpu.scala 106:29]
  wire  icache_io_instAxi_rd_valid; // @[playground/src/noop/cpu.scala 106:29]
  wire [63:0] icache_io_instAxi_rd_bits_data; // @[playground/src/noop/cpu.scala 106:29]
  wire  icache_io_instAxi_rd_bits_last; // @[playground/src/noop/cpu.scala 106:29]
  wire [31:0] icache_io_icRead_addr; // @[playground/src/noop/cpu.scala 106:29]
  wire [63:0] icache_io_icRead_inst; // @[playground/src/noop/cpu.scala 106:29]
  wire  icache_io_icRead_arvalid; // @[playground/src/noop/cpu.scala 106:29]
  wire  icache_io_icRead_ready; // @[playground/src/noop/cpu.scala 106:29]
  wire  icache_io_icRead_rvalid; // @[playground/src/noop/cpu.scala 106:29]
  wire  icache_io_flush; // @[playground/src/noop/cpu.scala 106:29]
  wire  dcache_clock; // @[playground/src/noop/cpu.scala 107:29]
  wire  dcache_reset; // @[playground/src/noop/cpu.scala 107:29]
  wire  dcache_io_dataAxi_wa_ready; // @[playground/src/noop/cpu.scala 107:29]
  wire  dcache_io_dataAxi_wa_valid; // @[playground/src/noop/cpu.scala 107:29]
  wire [31:0] dcache_io_dataAxi_wa_bits_addr; // @[playground/src/noop/cpu.scala 107:29]
  wire  dcache_io_dataAxi_wd_ready; // @[playground/src/noop/cpu.scala 107:29]
  wire  dcache_io_dataAxi_wd_valid; // @[playground/src/noop/cpu.scala 107:29]
  wire [63:0] dcache_io_dataAxi_wd_bits_data; // @[playground/src/noop/cpu.scala 107:29]
  wire  dcache_io_dataAxi_wd_bits_last; // @[playground/src/noop/cpu.scala 107:29]
  wire  dcache_io_dataAxi_ra_ready; // @[playground/src/noop/cpu.scala 107:29]
  wire  dcache_io_dataAxi_ra_valid; // @[playground/src/noop/cpu.scala 107:29]
  wire [31:0] dcache_io_dataAxi_ra_bits_addr; // @[playground/src/noop/cpu.scala 107:29]
  wire  dcache_io_dataAxi_rd_valid; // @[playground/src/noop/cpu.scala 107:29]
  wire [63:0] dcache_io_dataAxi_rd_bits_data; // @[playground/src/noop/cpu.scala 107:29]
  wire  dcache_io_dataAxi_rd_bits_last; // @[playground/src/noop/cpu.scala 107:29]
  wire [31:0] dcache_io_dcRW_addr; // @[playground/src/noop/cpu.scala 107:29]
  wire [63:0] dcache_io_dcRW_rdata; // @[playground/src/noop/cpu.scala 107:29]
  wire  dcache_io_dcRW_rvalid; // @[playground/src/noop/cpu.scala 107:29]
  wire [63:0] dcache_io_dcRW_wdata; // @[playground/src/noop/cpu.scala 107:29]
  wire [4:0] dcache_io_dcRW_dc_mode; // @[playground/src/noop/cpu.scala 107:29]
  wire [4:0] dcache_io_dcRW_amo; // @[playground/src/noop/cpu.scala 107:29]
  wire  dcache_io_dcRW_ready; // @[playground/src/noop/cpu.scala 107:29]
  wire  dcache_io_flush; // @[playground/src/noop/cpu.scala 107:29]
  wire  dcache_io_flush_out; // @[playground/src/noop/cpu.scala 107:29]
  wire  mem2Axi_clock; // @[playground/src/noop/cpu.scala 109:29]
  wire  mem2Axi_reset; // @[playground/src/noop/cpu.scala 109:29]
  wire [31:0] mem2Axi_io_dataIO_addr; // @[playground/src/noop/cpu.scala 109:29]
  wire [63:0] mem2Axi_io_dataIO_rdata; // @[playground/src/noop/cpu.scala 109:29]
  wire  mem2Axi_io_dataIO_rvalid; // @[playground/src/noop/cpu.scala 109:29]
  wire [63:0] mem2Axi_io_dataIO_wdata; // @[playground/src/noop/cpu.scala 109:29]
  wire [4:0] mem2Axi_io_dataIO_dc_mode; // @[playground/src/noop/cpu.scala 109:29]
  wire  mem2Axi_io_dataIO_ready; // @[playground/src/noop/cpu.scala 109:29]
  wire  mem2Axi_io_outAxi_wa_ready; // @[playground/src/noop/cpu.scala 109:29]
  wire  mem2Axi_io_outAxi_wa_valid; // @[playground/src/noop/cpu.scala 109:29]
  wire [3:0] mem2Axi_io_outAxi_wa_bits_id; // @[playground/src/noop/cpu.scala 109:29]
  wire [31:0] mem2Axi_io_outAxi_wa_bits_addr; // @[playground/src/noop/cpu.scala 109:29]
  wire [7:0] mem2Axi_io_outAxi_wa_bits_len; // @[playground/src/noop/cpu.scala 109:29]
  wire [2:0] mem2Axi_io_outAxi_wa_bits_size; // @[playground/src/noop/cpu.scala 109:29]
  wire [1:0] mem2Axi_io_outAxi_wa_bits_burst; // @[playground/src/noop/cpu.scala 109:29]
  wire  mem2Axi_io_outAxi_wd_ready; // @[playground/src/noop/cpu.scala 109:29]
  wire  mem2Axi_io_outAxi_wd_valid; // @[playground/src/noop/cpu.scala 109:29]
  wire [63:0] mem2Axi_io_outAxi_wd_bits_data; // @[playground/src/noop/cpu.scala 109:29]
  wire [7:0] mem2Axi_io_outAxi_wd_bits_strb; // @[playground/src/noop/cpu.scala 109:29]
  wire  mem2Axi_io_outAxi_wd_bits_last; // @[playground/src/noop/cpu.scala 109:29]
  wire  mem2Axi_io_outAxi_wr_ready; // @[playground/src/noop/cpu.scala 109:29]
  wire  mem2Axi_io_outAxi_wr_valid; // @[playground/src/noop/cpu.scala 109:29]
  wire [3:0] mem2Axi_io_outAxi_wr_bits_id; // @[playground/src/noop/cpu.scala 109:29]
  wire [1:0] mem2Axi_io_outAxi_wr_bits_resp; // @[playground/src/noop/cpu.scala 109:29]
  wire  mem2Axi_io_outAxi_ra_ready; // @[playground/src/noop/cpu.scala 109:29]
  wire  mem2Axi_io_outAxi_ra_valid; // @[playground/src/noop/cpu.scala 109:29]
  wire [3:0] mem2Axi_io_outAxi_ra_bits_id; // @[playground/src/noop/cpu.scala 109:29]
  wire [31:0] mem2Axi_io_outAxi_ra_bits_addr; // @[playground/src/noop/cpu.scala 109:29]
  wire [7:0] mem2Axi_io_outAxi_ra_bits_len; // @[playground/src/noop/cpu.scala 109:29]
  wire [2:0] mem2Axi_io_outAxi_ra_bits_size; // @[playground/src/noop/cpu.scala 109:29]
  wire [1:0] mem2Axi_io_outAxi_ra_bits_burst; // @[playground/src/noop/cpu.scala 109:29]
  wire  mem2Axi_io_outAxi_rd_ready; // @[playground/src/noop/cpu.scala 109:29]
  wire  mem2Axi_io_outAxi_rd_valid; // @[playground/src/noop/cpu.scala 109:29]
  wire [3:0] mem2Axi_io_outAxi_rd_bits_id; // @[playground/src/noop/cpu.scala 109:29]
  wire [63:0] mem2Axi_io_outAxi_rd_bits_data; // @[playground/src/noop/cpu.scala 109:29]
  wire [1:0] mem2Axi_io_outAxi_rd_bits_resp; // @[playground/src/noop/cpu.scala 109:29]
  wire  mem2Axi_io_outAxi_rd_bits_last; // @[playground/src/noop/cpu.scala 109:29]
  wire  flash2Axi_clock; // @[playground/src/noop/cpu.scala 110:29]
  wire  flash2Axi_reset; // @[playground/src/noop/cpu.scala 110:29]
  wire [31:0] flash2Axi_io_dataIO_addr; // @[playground/src/noop/cpu.scala 110:29]
  wire [63:0] flash2Axi_io_dataIO_rdata; // @[playground/src/noop/cpu.scala 110:29]
  wire  flash2Axi_io_dataIO_rvalid; // @[playground/src/noop/cpu.scala 110:29]
  wire [63:0] flash2Axi_io_dataIO_wdata; // @[playground/src/noop/cpu.scala 110:29]
  wire [4:0] flash2Axi_io_dataIO_dc_mode; // @[playground/src/noop/cpu.scala 110:29]
  wire  flash2Axi_io_dataIO_ready; // @[playground/src/noop/cpu.scala 110:29]
  wire  flash2Axi_io_outAxi_wa_ready; // @[playground/src/noop/cpu.scala 110:29]
  wire  flash2Axi_io_outAxi_wa_valid; // @[playground/src/noop/cpu.scala 110:29]
  wire [3:0] flash2Axi_io_outAxi_wa_bits_id; // @[playground/src/noop/cpu.scala 110:29]
  wire [31:0] flash2Axi_io_outAxi_wa_bits_addr; // @[playground/src/noop/cpu.scala 110:29]
  wire [7:0] flash2Axi_io_outAxi_wa_bits_len; // @[playground/src/noop/cpu.scala 110:29]
  wire [2:0] flash2Axi_io_outAxi_wa_bits_size; // @[playground/src/noop/cpu.scala 110:29]
  wire [1:0] flash2Axi_io_outAxi_wa_bits_burst; // @[playground/src/noop/cpu.scala 110:29]
  wire  flash2Axi_io_outAxi_wd_ready; // @[playground/src/noop/cpu.scala 110:29]
  wire  flash2Axi_io_outAxi_wd_valid; // @[playground/src/noop/cpu.scala 110:29]
  wire [63:0] flash2Axi_io_outAxi_wd_bits_data; // @[playground/src/noop/cpu.scala 110:29]
  wire [7:0] flash2Axi_io_outAxi_wd_bits_strb; // @[playground/src/noop/cpu.scala 110:29]
  wire  flash2Axi_io_outAxi_wd_bits_last; // @[playground/src/noop/cpu.scala 110:29]
  wire  flash2Axi_io_outAxi_wr_ready; // @[playground/src/noop/cpu.scala 110:29]
  wire  flash2Axi_io_outAxi_wr_valid; // @[playground/src/noop/cpu.scala 110:29]
  wire [3:0] flash2Axi_io_outAxi_wr_bits_id; // @[playground/src/noop/cpu.scala 110:29]
  wire [1:0] flash2Axi_io_outAxi_wr_bits_resp; // @[playground/src/noop/cpu.scala 110:29]
  wire  flash2Axi_io_outAxi_ra_ready; // @[playground/src/noop/cpu.scala 110:29]
  wire  flash2Axi_io_outAxi_ra_valid; // @[playground/src/noop/cpu.scala 110:29]
  wire [3:0] flash2Axi_io_outAxi_ra_bits_id; // @[playground/src/noop/cpu.scala 110:29]
  wire [31:0] flash2Axi_io_outAxi_ra_bits_addr; // @[playground/src/noop/cpu.scala 110:29]
  wire [7:0] flash2Axi_io_outAxi_ra_bits_len; // @[playground/src/noop/cpu.scala 110:29]
  wire [2:0] flash2Axi_io_outAxi_ra_bits_size; // @[playground/src/noop/cpu.scala 110:29]
  wire [1:0] flash2Axi_io_outAxi_ra_bits_burst; // @[playground/src/noop/cpu.scala 110:29]
  wire  flash2Axi_io_outAxi_rd_ready; // @[playground/src/noop/cpu.scala 110:29]
  wire  flash2Axi_io_outAxi_rd_valid; // @[playground/src/noop/cpu.scala 110:29]
  wire [3:0] flash2Axi_io_outAxi_rd_bits_id; // @[playground/src/noop/cpu.scala 110:29]
  wire [63:0] flash2Axi_io_outAxi_rd_bits_data; // @[playground/src/noop/cpu.scala 110:29]
  wire [1:0] flash2Axi_io_outAxi_rd_bits_resp; // @[playground/src/noop/cpu.scala 110:29]
  wire  flash2Axi_io_outAxi_rd_bits_last; // @[playground/src/noop/cpu.scala 110:29]
  wire  crossBar_clock; // @[playground/src/noop/cpu.scala 112:29]
  wire  crossBar_reset; // @[playground/src/noop/cpu.scala 112:29]
  wire  crossBar_io_icAxi_ra_ready; // @[playground/src/noop/cpu.scala 112:29]
  wire  crossBar_io_icAxi_ra_valid; // @[playground/src/noop/cpu.scala 112:29]
  wire [31:0] crossBar_io_icAxi_ra_bits_addr; // @[playground/src/noop/cpu.scala 112:29]
  wire  crossBar_io_icAxi_rd_valid; // @[playground/src/noop/cpu.scala 112:29]
  wire [63:0] crossBar_io_icAxi_rd_bits_data; // @[playground/src/noop/cpu.scala 112:29]
  wire  crossBar_io_icAxi_rd_bits_last; // @[playground/src/noop/cpu.scala 112:29]
  wire  crossBar_io_flashAxi_wa_ready; // @[playground/src/noop/cpu.scala 112:29]
  wire  crossBar_io_flashAxi_wa_valid; // @[playground/src/noop/cpu.scala 112:29]
  wire [3:0] crossBar_io_flashAxi_wa_bits_id; // @[playground/src/noop/cpu.scala 112:29]
  wire [31:0] crossBar_io_flashAxi_wa_bits_addr; // @[playground/src/noop/cpu.scala 112:29]
  wire [7:0] crossBar_io_flashAxi_wa_bits_len; // @[playground/src/noop/cpu.scala 112:29]
  wire [2:0] crossBar_io_flashAxi_wa_bits_size; // @[playground/src/noop/cpu.scala 112:29]
  wire [1:0] crossBar_io_flashAxi_wa_bits_burst; // @[playground/src/noop/cpu.scala 112:29]
  wire  crossBar_io_flashAxi_wd_ready; // @[playground/src/noop/cpu.scala 112:29]
  wire  crossBar_io_flashAxi_wd_valid; // @[playground/src/noop/cpu.scala 112:29]
  wire [63:0] crossBar_io_flashAxi_wd_bits_data; // @[playground/src/noop/cpu.scala 112:29]
  wire [7:0] crossBar_io_flashAxi_wd_bits_strb; // @[playground/src/noop/cpu.scala 112:29]
  wire  crossBar_io_flashAxi_wd_bits_last; // @[playground/src/noop/cpu.scala 112:29]
  wire  crossBar_io_flashAxi_wr_ready; // @[playground/src/noop/cpu.scala 112:29]
  wire  crossBar_io_flashAxi_wr_valid; // @[playground/src/noop/cpu.scala 112:29]
  wire [3:0] crossBar_io_flashAxi_wr_bits_id; // @[playground/src/noop/cpu.scala 112:29]
  wire [1:0] crossBar_io_flashAxi_wr_bits_resp; // @[playground/src/noop/cpu.scala 112:29]
  wire  crossBar_io_flashAxi_ra_ready; // @[playground/src/noop/cpu.scala 112:29]
  wire  crossBar_io_flashAxi_ra_valid; // @[playground/src/noop/cpu.scala 112:29]
  wire [3:0] crossBar_io_flashAxi_ra_bits_id; // @[playground/src/noop/cpu.scala 112:29]
  wire [31:0] crossBar_io_flashAxi_ra_bits_addr; // @[playground/src/noop/cpu.scala 112:29]
  wire [7:0] crossBar_io_flashAxi_ra_bits_len; // @[playground/src/noop/cpu.scala 112:29]
  wire [2:0] crossBar_io_flashAxi_ra_bits_size; // @[playground/src/noop/cpu.scala 112:29]
  wire [1:0] crossBar_io_flashAxi_ra_bits_burst; // @[playground/src/noop/cpu.scala 112:29]
  wire  crossBar_io_flashAxi_rd_ready; // @[playground/src/noop/cpu.scala 112:29]
  wire  crossBar_io_flashAxi_rd_valid; // @[playground/src/noop/cpu.scala 112:29]
  wire [3:0] crossBar_io_flashAxi_rd_bits_id; // @[playground/src/noop/cpu.scala 112:29]
  wire [63:0] crossBar_io_flashAxi_rd_bits_data; // @[playground/src/noop/cpu.scala 112:29]
  wire [1:0] crossBar_io_flashAxi_rd_bits_resp; // @[playground/src/noop/cpu.scala 112:29]
  wire  crossBar_io_flashAxi_rd_bits_last; // @[playground/src/noop/cpu.scala 112:29]
  wire  crossBar_io_memAxi_wa_ready; // @[playground/src/noop/cpu.scala 112:29]
  wire  crossBar_io_memAxi_wa_valid; // @[playground/src/noop/cpu.scala 112:29]
  wire [31:0] crossBar_io_memAxi_wa_bits_addr; // @[playground/src/noop/cpu.scala 112:29]
  wire  crossBar_io_memAxi_wd_ready; // @[playground/src/noop/cpu.scala 112:29]
  wire  crossBar_io_memAxi_wd_valid; // @[playground/src/noop/cpu.scala 112:29]
  wire [63:0] crossBar_io_memAxi_wd_bits_data; // @[playground/src/noop/cpu.scala 112:29]
  wire  crossBar_io_memAxi_wd_bits_last; // @[playground/src/noop/cpu.scala 112:29]
  wire  crossBar_io_memAxi_ra_ready; // @[playground/src/noop/cpu.scala 112:29]
  wire  crossBar_io_memAxi_ra_valid; // @[playground/src/noop/cpu.scala 112:29]
  wire [31:0] crossBar_io_memAxi_ra_bits_addr; // @[playground/src/noop/cpu.scala 112:29]
  wire  crossBar_io_memAxi_rd_valid; // @[playground/src/noop/cpu.scala 112:29]
  wire [63:0] crossBar_io_memAxi_rd_bits_data; // @[playground/src/noop/cpu.scala 112:29]
  wire  crossBar_io_memAxi_rd_bits_last; // @[playground/src/noop/cpu.scala 112:29]
  wire  crossBar_io_mmioAxi_wa_ready; // @[playground/src/noop/cpu.scala 112:29]
  wire  crossBar_io_mmioAxi_wa_valid; // @[playground/src/noop/cpu.scala 112:29]
  wire [3:0] crossBar_io_mmioAxi_wa_bits_id; // @[playground/src/noop/cpu.scala 112:29]
  wire [31:0] crossBar_io_mmioAxi_wa_bits_addr; // @[playground/src/noop/cpu.scala 112:29]
  wire [7:0] crossBar_io_mmioAxi_wa_bits_len; // @[playground/src/noop/cpu.scala 112:29]
  wire [2:0] crossBar_io_mmioAxi_wa_bits_size; // @[playground/src/noop/cpu.scala 112:29]
  wire [1:0] crossBar_io_mmioAxi_wa_bits_burst; // @[playground/src/noop/cpu.scala 112:29]
  wire  crossBar_io_mmioAxi_wd_ready; // @[playground/src/noop/cpu.scala 112:29]
  wire  crossBar_io_mmioAxi_wd_valid; // @[playground/src/noop/cpu.scala 112:29]
  wire [63:0] crossBar_io_mmioAxi_wd_bits_data; // @[playground/src/noop/cpu.scala 112:29]
  wire [7:0] crossBar_io_mmioAxi_wd_bits_strb; // @[playground/src/noop/cpu.scala 112:29]
  wire  crossBar_io_mmioAxi_wd_bits_last; // @[playground/src/noop/cpu.scala 112:29]
  wire  crossBar_io_mmioAxi_wr_ready; // @[playground/src/noop/cpu.scala 112:29]
  wire  crossBar_io_mmioAxi_wr_valid; // @[playground/src/noop/cpu.scala 112:29]
  wire [3:0] crossBar_io_mmioAxi_wr_bits_id; // @[playground/src/noop/cpu.scala 112:29]
  wire [1:0] crossBar_io_mmioAxi_wr_bits_resp; // @[playground/src/noop/cpu.scala 112:29]
  wire  crossBar_io_mmioAxi_ra_ready; // @[playground/src/noop/cpu.scala 112:29]
  wire  crossBar_io_mmioAxi_ra_valid; // @[playground/src/noop/cpu.scala 112:29]
  wire [3:0] crossBar_io_mmioAxi_ra_bits_id; // @[playground/src/noop/cpu.scala 112:29]
  wire [31:0] crossBar_io_mmioAxi_ra_bits_addr; // @[playground/src/noop/cpu.scala 112:29]
  wire [7:0] crossBar_io_mmioAxi_ra_bits_len; // @[playground/src/noop/cpu.scala 112:29]
  wire [2:0] crossBar_io_mmioAxi_ra_bits_size; // @[playground/src/noop/cpu.scala 112:29]
  wire [1:0] crossBar_io_mmioAxi_ra_bits_burst; // @[playground/src/noop/cpu.scala 112:29]
  wire  crossBar_io_mmioAxi_rd_ready; // @[playground/src/noop/cpu.scala 112:29]
  wire  crossBar_io_mmioAxi_rd_valid; // @[playground/src/noop/cpu.scala 112:29]
  wire [3:0] crossBar_io_mmioAxi_rd_bits_id; // @[playground/src/noop/cpu.scala 112:29]
  wire [63:0] crossBar_io_mmioAxi_rd_bits_data; // @[playground/src/noop/cpu.scala 112:29]
  wire [1:0] crossBar_io_mmioAxi_rd_bits_resp; // @[playground/src/noop/cpu.scala 112:29]
  wire  crossBar_io_mmioAxi_rd_bits_last; // @[playground/src/noop/cpu.scala 112:29]
  wire  crossBar_io_outAxi_wa_ready; // @[playground/src/noop/cpu.scala 112:29]
  wire  crossBar_io_outAxi_wa_valid; // @[playground/src/noop/cpu.scala 112:29]
  wire [3:0] crossBar_io_outAxi_wa_bits_id; // @[playground/src/noop/cpu.scala 112:29]
  wire [31:0] crossBar_io_outAxi_wa_bits_addr; // @[playground/src/noop/cpu.scala 112:29]
  wire [7:0] crossBar_io_outAxi_wa_bits_len; // @[playground/src/noop/cpu.scala 112:29]
  wire [2:0] crossBar_io_outAxi_wa_bits_size; // @[playground/src/noop/cpu.scala 112:29]
  wire [1:0] crossBar_io_outAxi_wa_bits_burst; // @[playground/src/noop/cpu.scala 112:29]
  wire  crossBar_io_outAxi_wd_ready; // @[playground/src/noop/cpu.scala 112:29]
  wire  crossBar_io_outAxi_wd_valid; // @[playground/src/noop/cpu.scala 112:29]
  wire [63:0] crossBar_io_outAxi_wd_bits_data; // @[playground/src/noop/cpu.scala 112:29]
  wire [7:0] crossBar_io_outAxi_wd_bits_strb; // @[playground/src/noop/cpu.scala 112:29]
  wire  crossBar_io_outAxi_wd_bits_last; // @[playground/src/noop/cpu.scala 112:29]
  wire  crossBar_io_outAxi_wr_ready; // @[playground/src/noop/cpu.scala 112:29]
  wire  crossBar_io_outAxi_wr_valid; // @[playground/src/noop/cpu.scala 112:29]
  wire [3:0] crossBar_io_outAxi_wr_bits_id; // @[playground/src/noop/cpu.scala 112:29]
  wire [1:0] crossBar_io_outAxi_wr_bits_resp; // @[playground/src/noop/cpu.scala 112:29]
  wire  crossBar_io_outAxi_ra_ready; // @[playground/src/noop/cpu.scala 112:29]
  wire  crossBar_io_outAxi_ra_valid; // @[playground/src/noop/cpu.scala 112:29]
  wire [3:0] crossBar_io_outAxi_ra_bits_id; // @[playground/src/noop/cpu.scala 112:29]
  wire [31:0] crossBar_io_outAxi_ra_bits_addr; // @[playground/src/noop/cpu.scala 112:29]
  wire [7:0] crossBar_io_outAxi_ra_bits_len; // @[playground/src/noop/cpu.scala 112:29]
  wire [2:0] crossBar_io_outAxi_ra_bits_size; // @[playground/src/noop/cpu.scala 112:29]
  wire [1:0] crossBar_io_outAxi_ra_bits_burst; // @[playground/src/noop/cpu.scala 112:29]
  wire  crossBar_io_outAxi_rd_ready; // @[playground/src/noop/cpu.scala 112:29]
  wire  crossBar_io_outAxi_rd_valid; // @[playground/src/noop/cpu.scala 112:29]
  wire [3:0] crossBar_io_outAxi_rd_bits_id; // @[playground/src/noop/cpu.scala 112:29]
  wire [63:0] crossBar_io_outAxi_rd_bits_data; // @[playground/src/noop/cpu.scala 112:29]
  wire [1:0] crossBar_io_outAxi_rd_bits_resp; // @[playground/src/noop/cpu.scala 112:29]
  wire  crossBar_io_outAxi_rd_bits_last; // @[playground/src/noop/cpu.scala 112:29]
  wire  crossBar_io_selectMem; // @[playground/src/noop/cpu.scala 112:29]
  wire  fetchCrossbar_clock; // @[playground/src/noop/cpu.scala 113:31]
  wire  fetchCrossbar_reset; // @[playground/src/noop/cpu.scala 113:31]
  wire [31:0] fetchCrossbar_io_instIO_addr; // @[playground/src/noop/cpu.scala 113:31]
  wire [63:0] fetchCrossbar_io_instIO_inst; // @[playground/src/noop/cpu.scala 113:31]
  wire  fetchCrossbar_io_instIO_arvalid; // @[playground/src/noop/cpu.scala 113:31]
  wire  fetchCrossbar_io_instIO_rvalid; // @[playground/src/noop/cpu.scala 113:31]
  wire [31:0] fetchCrossbar_io_icRead_addr; // @[playground/src/noop/cpu.scala 113:31]
  wire [63:0] fetchCrossbar_io_icRead_inst; // @[playground/src/noop/cpu.scala 113:31]
  wire  fetchCrossbar_io_icRead_arvalid; // @[playground/src/noop/cpu.scala 113:31]
  wire  fetchCrossbar_io_icRead_rvalid; // @[playground/src/noop/cpu.scala 113:31]
  wire [31:0] fetchCrossbar_io_flashRead_addr; // @[playground/src/noop/cpu.scala 113:31]
  wire [63:0] fetchCrossbar_io_flashRead_rdata; // @[playground/src/noop/cpu.scala 113:31]
  wire  fetchCrossbar_io_flashRead_rvalid; // @[playground/src/noop/cpu.scala 113:31]
  wire [4:0] fetchCrossbar_io_flashRead_dc_mode; // @[playground/src/noop/cpu.scala 113:31]
  wire  split64to32_clock; // @[playground/src/noop/cpu.scala 114:29]
  wire  split64to32_reset; // @[playground/src/noop/cpu.scala 114:29]
  wire [31:0] split64to32_io_data_in_addr; // @[playground/src/noop/cpu.scala 114:29]
  wire [63:0] split64to32_io_data_in_rdata; // @[playground/src/noop/cpu.scala 114:29]
  wire  split64to32_io_data_in_rvalid; // @[playground/src/noop/cpu.scala 114:29]
  wire [4:0] split64to32_io_data_in_dc_mode; // @[playground/src/noop/cpu.scala 114:29]
  wire [31:0] split64to32_io_data_out_addr; // @[playground/src/noop/cpu.scala 114:29]
  wire [63:0] split64to32_io_data_out_rdata; // @[playground/src/noop/cpu.scala 114:29]
  wire  split64to32_io_data_out_rvalid; // @[playground/src/noop/cpu.scala 114:29]
  wire [4:0] split64to32_io_data_out_dc_mode; // @[playground/src/noop/cpu.scala 114:29]
  wire  split64to32_io_data_out_ready; // @[playground/src/noop/cpu.scala 114:29]
  wire  memCrossbar_clock; // @[playground/src/noop/cpu.scala 115:29]
  wire  memCrossbar_reset; // @[playground/src/noop/cpu.scala 115:29]
  wire [31:0] memCrossbar_io_dataRW_addr; // @[playground/src/noop/cpu.scala 115:29]
  wire [63:0] memCrossbar_io_dataRW_rdata; // @[playground/src/noop/cpu.scala 115:29]
  wire  memCrossbar_io_dataRW_rvalid; // @[playground/src/noop/cpu.scala 115:29]
  wire [63:0] memCrossbar_io_dataRW_wdata; // @[playground/src/noop/cpu.scala 115:29]
  wire [4:0] memCrossbar_io_dataRW_dc_mode; // @[playground/src/noop/cpu.scala 115:29]
  wire [4:0] memCrossbar_io_dataRW_amo; // @[playground/src/noop/cpu.scala 115:29]
  wire  memCrossbar_io_dataRW_ready; // @[playground/src/noop/cpu.scala 115:29]
  wire [31:0] memCrossbar_io_mmio_addr; // @[playground/src/noop/cpu.scala 115:29]
  wire [63:0] memCrossbar_io_mmio_rdata; // @[playground/src/noop/cpu.scala 115:29]
  wire  memCrossbar_io_mmio_rvalid; // @[playground/src/noop/cpu.scala 115:29]
  wire [63:0] memCrossbar_io_mmio_wdata; // @[playground/src/noop/cpu.scala 115:29]
  wire [4:0] memCrossbar_io_mmio_dc_mode; // @[playground/src/noop/cpu.scala 115:29]
  wire  memCrossbar_io_mmio_ready; // @[playground/src/noop/cpu.scala 115:29]
  wire [31:0] memCrossbar_io_dcRW_addr; // @[playground/src/noop/cpu.scala 115:29]
  wire [63:0] memCrossbar_io_dcRW_rdata; // @[playground/src/noop/cpu.scala 115:29]
  wire  memCrossbar_io_dcRW_rvalid; // @[playground/src/noop/cpu.scala 115:29]
  wire [63:0] memCrossbar_io_dcRW_wdata; // @[playground/src/noop/cpu.scala 115:29]
  wire [4:0] memCrossbar_io_dcRW_dc_mode; // @[playground/src/noop/cpu.scala 115:29]
  wire [4:0] memCrossbar_io_dcRW_amo; // @[playground/src/noop/cpu.scala 115:29]
  wire  memCrossbar_io_dcRW_ready; // @[playground/src/noop/cpu.scala 115:29]
  wire [31:0] memCrossbar_io_clintIO_addr; // @[playground/src/noop/cpu.scala 115:29]
  wire [63:0] memCrossbar_io_clintIO_rdata; // @[playground/src/noop/cpu.scala 115:29]
  wire [63:0] memCrossbar_io_clintIO_wdata; // @[playground/src/noop/cpu.scala 115:29]
  wire  memCrossbar_io_clintIO_wvalid; // @[playground/src/noop/cpu.scala 115:29]
  wire [31:0] memCrossbar_io_plicIO_addr; // @[playground/src/noop/cpu.scala 115:29]
  wire [63:0] memCrossbar_io_plicIO_rdata; // @[playground/src/noop/cpu.scala 115:29]
  wire [63:0] memCrossbar_io_plicIO_wdata; // @[playground/src/noop/cpu.scala 115:29]
  wire  memCrossbar_io_plicIO_wvalid; // @[playground/src/noop/cpu.scala 115:29]
  wire  memCrossbar_io_plicIO_arvalid; // @[playground/src/noop/cpu.scala 115:29]
  wire  tlb_if_clock; // @[playground/src/noop/cpu.scala 116:30]
  wire  tlb_if_reset; // @[playground/src/noop/cpu.scala 116:30]
  wire [63:0] tlb_if_io_va2pa_vaddr; // @[playground/src/noop/cpu.scala 116:30]
  wire  tlb_if_io_va2pa_vvalid; // @[playground/src/noop/cpu.scala 116:30]
  wire  tlb_if_io_va2pa_ready; // @[playground/src/noop/cpu.scala 116:30]
  wire [31:0] tlb_if_io_va2pa_paddr; // @[playground/src/noop/cpu.scala 116:30]
  wire  tlb_if_io_va2pa_pvalid; // @[playground/src/noop/cpu.scala 116:30]
  wire [63:0] tlb_if_io_va2pa_tlb_excep_cause; // @[playground/src/noop/cpu.scala 116:30]
  wire [63:0] tlb_if_io_va2pa_tlb_excep_tval; // @[playground/src/noop/cpu.scala 116:30]
  wire  tlb_if_io_va2pa_tlb_excep_en; // @[playground/src/noop/cpu.scala 116:30]
  wire [1:0] tlb_if_io_mmuState_priv; // @[playground/src/noop/cpu.scala 116:30]
  wire [63:0] tlb_if_io_mmuState_mstatus; // @[playground/src/noop/cpu.scala 116:30]
  wire [63:0] tlb_if_io_mmuState_satp; // @[playground/src/noop/cpu.scala 116:30]
  wire  tlb_if_io_flush; // @[playground/src/noop/cpu.scala 116:30]
  wire [31:0] tlb_if_io_dcacheRW_addr; // @[playground/src/noop/cpu.scala 116:30]
  wire [63:0] tlb_if_io_dcacheRW_rdata; // @[playground/src/noop/cpu.scala 116:30]
  wire  tlb_if_io_dcacheRW_rvalid; // @[playground/src/noop/cpu.scala 116:30]
  wire [63:0] tlb_if_io_dcacheRW_wdata; // @[playground/src/noop/cpu.scala 116:30]
  wire [4:0] tlb_if_io_dcacheRW_dc_mode; // @[playground/src/noop/cpu.scala 116:30]
  wire  tlb_if_io_dcacheRW_ready; // @[playground/src/noop/cpu.scala 116:30]
  wire  tlb_mem_clock; // @[playground/src/noop/cpu.scala 117:30]
  wire  tlb_mem_reset; // @[playground/src/noop/cpu.scala 117:30]
  wire [63:0] tlb_mem_io_va2pa_vaddr; // @[playground/src/noop/cpu.scala 117:30]
  wire  tlb_mem_io_va2pa_vvalid; // @[playground/src/noop/cpu.scala 117:30]
  wire [1:0] tlb_mem_io_va2pa_m_type; // @[playground/src/noop/cpu.scala 117:30]
  wire  tlb_mem_io_va2pa_ready; // @[playground/src/noop/cpu.scala 117:30]
  wire [31:0] tlb_mem_io_va2pa_paddr; // @[playground/src/noop/cpu.scala 117:30]
  wire  tlb_mem_io_va2pa_pvalid; // @[playground/src/noop/cpu.scala 117:30]
  wire [63:0] tlb_mem_io_va2pa_tlb_excep_cause; // @[playground/src/noop/cpu.scala 117:30]
  wire [63:0] tlb_mem_io_va2pa_tlb_excep_tval; // @[playground/src/noop/cpu.scala 117:30]
  wire  tlb_mem_io_va2pa_tlb_excep_en; // @[playground/src/noop/cpu.scala 117:30]
  wire [1:0] tlb_mem_io_mmuState_priv; // @[playground/src/noop/cpu.scala 117:30]
  wire [63:0] tlb_mem_io_mmuState_mstatus; // @[playground/src/noop/cpu.scala 117:30]
  wire [63:0] tlb_mem_io_mmuState_satp; // @[playground/src/noop/cpu.scala 117:30]
  wire  tlb_mem_io_flush; // @[playground/src/noop/cpu.scala 117:30]
  wire [31:0] tlb_mem_io_dcacheRW_addr; // @[playground/src/noop/cpu.scala 117:30]
  wire [63:0] tlb_mem_io_dcacheRW_rdata; // @[playground/src/noop/cpu.scala 117:30]
  wire  tlb_mem_io_dcacheRW_rvalid; // @[playground/src/noop/cpu.scala 117:30]
  wire [63:0] tlb_mem_io_dcacheRW_wdata; // @[playground/src/noop/cpu.scala 117:30]
  wire [4:0] tlb_mem_io_dcacheRW_dc_mode; // @[playground/src/noop/cpu.scala 117:30]
  wire  tlb_mem_io_dcacheRW_ready; // @[playground/src/noop/cpu.scala 117:30]
  wire  dcSelector_clock; // @[playground/src/noop/cpu.scala 118:29]
  wire  dcSelector_reset; // @[playground/src/noop/cpu.scala 118:29]
  wire [31:0] dcSelector_io_tlb_if2dc_addr; // @[playground/src/noop/cpu.scala 118:29]
  wire [63:0] dcSelector_io_tlb_if2dc_rdata; // @[playground/src/noop/cpu.scala 118:29]
  wire  dcSelector_io_tlb_if2dc_rvalid; // @[playground/src/noop/cpu.scala 118:29]
  wire [63:0] dcSelector_io_tlb_if2dc_wdata; // @[playground/src/noop/cpu.scala 118:29]
  wire [4:0] dcSelector_io_tlb_if2dc_dc_mode; // @[playground/src/noop/cpu.scala 118:29]
  wire  dcSelector_io_tlb_if2dc_ready; // @[playground/src/noop/cpu.scala 118:29]
  wire [31:0] dcSelector_io_tlb_mem2dc_addr; // @[playground/src/noop/cpu.scala 118:29]
  wire [63:0] dcSelector_io_tlb_mem2dc_rdata; // @[playground/src/noop/cpu.scala 118:29]
  wire  dcSelector_io_tlb_mem2dc_rvalid; // @[playground/src/noop/cpu.scala 118:29]
  wire [63:0] dcSelector_io_tlb_mem2dc_wdata; // @[playground/src/noop/cpu.scala 118:29]
  wire [4:0] dcSelector_io_tlb_mem2dc_dc_mode; // @[playground/src/noop/cpu.scala 118:29]
  wire  dcSelector_io_tlb_mem2dc_ready; // @[playground/src/noop/cpu.scala 118:29]
  wire [31:0] dcSelector_io_mem2dc_addr; // @[playground/src/noop/cpu.scala 118:29]
  wire [63:0] dcSelector_io_mem2dc_rdata; // @[playground/src/noop/cpu.scala 118:29]
  wire  dcSelector_io_mem2dc_rvalid; // @[playground/src/noop/cpu.scala 118:29]
  wire [63:0] dcSelector_io_mem2dc_wdata; // @[playground/src/noop/cpu.scala 118:29]
  wire [4:0] dcSelector_io_mem2dc_dc_mode; // @[playground/src/noop/cpu.scala 118:29]
  wire [4:0] dcSelector_io_mem2dc_amo; // @[playground/src/noop/cpu.scala 118:29]
  wire  dcSelector_io_mem2dc_ready; // @[playground/src/noop/cpu.scala 118:29]
  wire [31:0] dcSelector_io_dma2dc_addr; // @[playground/src/noop/cpu.scala 118:29]
  wire [63:0] dcSelector_io_dma2dc_rdata; // @[playground/src/noop/cpu.scala 118:29]
  wire  dcSelector_io_dma2dc_rvalid; // @[playground/src/noop/cpu.scala 118:29]
  wire [63:0] dcSelector_io_dma2dc_wdata; // @[playground/src/noop/cpu.scala 118:29]
  wire [4:0] dcSelector_io_dma2dc_dc_mode; // @[playground/src/noop/cpu.scala 118:29]
  wire  dcSelector_io_dma2dc_ready; // @[playground/src/noop/cpu.scala 118:29]
  wire [31:0] dcSelector_io_select_addr; // @[playground/src/noop/cpu.scala 118:29]
  wire [63:0] dcSelector_io_select_rdata; // @[playground/src/noop/cpu.scala 118:29]
  wire  dcSelector_io_select_rvalid; // @[playground/src/noop/cpu.scala 118:29]
  wire [63:0] dcSelector_io_select_wdata; // @[playground/src/noop/cpu.scala 118:29]
  wire [4:0] dcSelector_io_select_dc_mode; // @[playground/src/noop/cpu.scala 118:29]
  wire [4:0] dcSelector_io_select_amo; // @[playground/src/noop/cpu.scala 118:29]
  wire  dcSelector_io_select_ready; // @[playground/src/noop/cpu.scala 118:29]
  wire  clint_clock; // @[playground/src/noop/cpu.scala 119:29]
  wire  clint_reset; // @[playground/src/noop/cpu.scala 119:29]
  wire [31:0] clint_io_rw_addr; // @[playground/src/noop/cpu.scala 119:29]
  wire [63:0] clint_io_rw_rdata; // @[playground/src/noop/cpu.scala 119:29]
  wire [63:0] clint_io_rw_wdata; // @[playground/src/noop/cpu.scala 119:29]
  wire  clint_io_rw_wvalid; // @[playground/src/noop/cpu.scala 119:29]
  wire  clint_io_intr_raise; // @[playground/src/noop/cpu.scala 119:29]
  wire  clint_io_intr_clear; // @[playground/src/noop/cpu.scala 119:29]
  wire  clint_io_intr_msip_raise; // @[playground/src/noop/cpu.scala 119:29]
  wire  clint_io_intr_msip_clear; // @[playground/src/noop/cpu.scala 119:29]
  wire  plic_clock; // @[playground/src/noop/cpu.scala 120:29]
  wire  plic_reset; // @[playground/src/noop/cpu.scala 120:29]
  wire  plic_io_intr_in1; // @[playground/src/noop/cpu.scala 120:29]
  wire  plic_io_intr_out_m_raise; // @[playground/src/noop/cpu.scala 120:29]
  wire  plic_io_intr_out_m_clear; // @[playground/src/noop/cpu.scala 120:29]
  wire  plic_io_intr_out_s_raise; // @[playground/src/noop/cpu.scala 120:29]
  wire  plic_io_intr_out_s_clear; // @[playground/src/noop/cpu.scala 120:29]
  wire [31:0] plic_io_rw_addr; // @[playground/src/noop/cpu.scala 120:29]
  wire [63:0] plic_io_rw_rdata; // @[playground/src/noop/cpu.scala 120:29]
  wire [63:0] plic_io_rw_wdata; // @[playground/src/noop/cpu.scala 120:29]
  wire  plic_io_rw_wvalid; // @[playground/src/noop/cpu.scala 120:29]
  wire  plic_io_rw_arvalid; // @[playground/src/noop/cpu.scala 120:29]
  wire  dmaBridge_clock; // @[playground/src/noop/cpu.scala 121:29]
  wire  dmaBridge_reset; // @[playground/src/noop/cpu.scala 121:29]
  wire  dmaBridge_io_dmaAxi_awready; // @[playground/src/noop/cpu.scala 121:29]
  wire  dmaBridge_io_dmaAxi_awvalid; // @[playground/src/noop/cpu.scala 121:29]
  wire [31:0] dmaBridge_io_dmaAxi_awaddr; // @[playground/src/noop/cpu.scala 121:29]
  wire [3:0] dmaBridge_io_dmaAxi_awid; // @[playground/src/noop/cpu.scala 121:29]
  wire [7:0] dmaBridge_io_dmaAxi_awlen; // @[playground/src/noop/cpu.scala 121:29]
  wire [2:0] dmaBridge_io_dmaAxi_awsize; // @[playground/src/noop/cpu.scala 121:29]
  wire  dmaBridge_io_dmaAxi_wready; // @[playground/src/noop/cpu.scala 121:29]
  wire  dmaBridge_io_dmaAxi_wvalid; // @[playground/src/noop/cpu.scala 121:29]
  wire [63:0] dmaBridge_io_dmaAxi_wdata; // @[playground/src/noop/cpu.scala 121:29]
  wire [7:0] dmaBridge_io_dmaAxi_wstrb; // @[playground/src/noop/cpu.scala 121:29]
  wire  dmaBridge_io_dmaAxi_bready; // @[playground/src/noop/cpu.scala 121:29]
  wire  dmaBridge_io_dmaAxi_bvalid; // @[playground/src/noop/cpu.scala 121:29]
  wire [3:0] dmaBridge_io_dmaAxi_bid; // @[playground/src/noop/cpu.scala 121:29]
  wire  dmaBridge_io_dmaAxi_arready; // @[playground/src/noop/cpu.scala 121:29]
  wire  dmaBridge_io_dmaAxi_arvalid; // @[playground/src/noop/cpu.scala 121:29]
  wire [31:0] dmaBridge_io_dmaAxi_araddr; // @[playground/src/noop/cpu.scala 121:29]
  wire [3:0] dmaBridge_io_dmaAxi_arid; // @[playground/src/noop/cpu.scala 121:29]
  wire [7:0] dmaBridge_io_dmaAxi_arlen; // @[playground/src/noop/cpu.scala 121:29]
  wire [2:0] dmaBridge_io_dmaAxi_arsize; // @[playground/src/noop/cpu.scala 121:29]
  wire  dmaBridge_io_dmaAxi_rready; // @[playground/src/noop/cpu.scala 121:29]
  wire  dmaBridge_io_dmaAxi_rvalid; // @[playground/src/noop/cpu.scala 121:29]
  wire [63:0] dmaBridge_io_dmaAxi_rdata; // @[playground/src/noop/cpu.scala 121:29]
  wire  dmaBridge_io_dmaAxi_rlast; // @[playground/src/noop/cpu.scala 121:29]
  wire [3:0] dmaBridge_io_dmaAxi_rid; // @[playground/src/noop/cpu.scala 121:29]
  wire [31:0] dmaBridge_io_dcRW_addr; // @[playground/src/noop/cpu.scala 121:29]
  wire [63:0] dmaBridge_io_dcRW_rdata; // @[playground/src/noop/cpu.scala 121:29]
  wire  dmaBridge_io_dcRW_rvalid; // @[playground/src/noop/cpu.scala 121:29]
  wire [63:0] dmaBridge_io_dcRW_wdata; // @[playground/src/noop/cpu.scala 121:29]
  wire [4:0] dmaBridge_io_dcRW_dc_mode; // @[playground/src/noop/cpu.scala 121:29]
  wire  dmaBridge_io_dcRW_ready; // @[playground/src/noop/cpu.scala 121:29]
  Fetch fetch ( // @[playground/src/noop/cpu.scala 96:29]
    .clock(fetch_clock),
    .reset(fetch_reset),
    .io_instRead_addr(fetch_io_instRead_addr),
    .io_instRead_inst(fetch_io_instRead_inst),
    .io_instRead_arvalid(fetch_io_instRead_arvalid),
    .io_instRead_rvalid(fetch_io_instRead_rvalid),
    .io_va2pa_vaddr(fetch_io_va2pa_vaddr),
    .io_va2pa_vvalid(fetch_io_va2pa_vvalid),
    .io_va2pa_paddr(fetch_io_va2pa_paddr),
    .io_va2pa_pvalid(fetch_io_va2pa_pvalid),
    .io_va2pa_tlb_excep_cause(fetch_io_va2pa_tlb_excep_cause),
    .io_va2pa_tlb_excep_tval(fetch_io_va2pa_tlb_excep_tval),
    .io_va2pa_tlb_excep_en(fetch_io_va2pa_tlb_excep_en),
    .io_reg2if_seq_pc(fetch_io_reg2if_seq_pc),
    .io_reg2if_valid(fetch_io_reg2if_valid),
    .io_wb2if_seq_pc(fetch_io_wb2if_seq_pc),
    .io_wb2if_valid(fetch_io_wb2if_valid),
    .io_recov(fetch_io_recov),
    .io_intr_in_en(fetch_io_intr_in_en),
    .io_intr_in_cause(fetch_io_intr_in_cause),
    .io_branchFail_seq_pc(fetch_io_branchFail_seq_pc),
    .io_branchFail_valid(fetch_io_branchFail_valid),
    .io_if2id_inst(fetch_io_if2id_inst),
    .io_if2id_pc(fetch_io_if2id_pc),
    .io_if2id_excep_cause(fetch_io_if2id_excep_cause),
    .io_if2id_excep_tval(fetch_io_if2id_excep_tval),
    .io_if2id_excep_en(fetch_io_if2id_excep_en),
    .io_if2id_excep_pc(fetch_io_if2id_excep_pc),
    .io_if2id_drop(fetch_io_if2id_drop),
    .io_if2id_stall(fetch_io_if2id_stall),
    .io_if2id_recov(fetch_io_if2id_recov),
    .io_if2id_valid(fetch_io_if2id_valid),
    .io_if2id_ready(fetch_io_if2id_ready)
  );
  Decode decode ( // @[playground/src/noop/cpu.scala 97:29]
    .clock(decode_clock),
    .reset(decode_reset),
    .io_if2id_inst(decode_io_if2id_inst),
    .io_if2id_pc(decode_io_if2id_pc),
    .io_if2id_excep_cause(decode_io_if2id_excep_cause),
    .io_if2id_excep_tval(decode_io_if2id_excep_tval),
    .io_if2id_excep_en(decode_io_if2id_excep_en),
    .io_if2id_excep_pc(decode_io_if2id_excep_pc),
    .io_if2id_drop(decode_io_if2id_drop),
    .io_if2id_stall(decode_io_if2id_stall),
    .io_if2id_recov(decode_io_if2id_recov),
    .io_if2id_valid(decode_io_if2id_valid),
    .io_if2id_ready(decode_io_if2id_ready),
    .io_id2df_inst(decode_io_id2df_inst),
    .io_id2df_pc(decode_io_id2df_pc),
    .io_id2df_excep_cause(decode_io_id2df_excep_cause),
    .io_id2df_excep_tval(decode_io_id2df_excep_tval),
    .io_id2df_excep_en(decode_io_id2df_excep_en),
    .io_id2df_excep_pc(decode_io_id2df_excep_pc),
    .io_id2df_excep_etype(decode_io_id2df_excep_etype),
    .io_id2df_ctrl_aluOp(decode_io_id2df_ctrl_aluOp),
    .io_id2df_ctrl_aluWidth(decode_io_id2df_ctrl_aluWidth),
    .io_id2df_ctrl_dcMode(decode_io_id2df_ctrl_dcMode),
    .io_id2df_ctrl_writeRegEn(decode_io_id2df_ctrl_writeRegEn),
    .io_id2df_ctrl_writeCSREn(decode_io_id2df_ctrl_writeCSREn),
    .io_id2df_ctrl_brType(decode_io_id2df_ctrl_brType),
    .io_id2df_rs1(decode_io_id2df_rs1),
    .io_id2df_rrs1(decode_io_id2df_rrs1),
    .io_id2df_rs1_d(decode_io_id2df_rs1_d),
    .io_id2df_rs2(decode_io_id2df_rs2),
    .io_id2df_rrs2(decode_io_id2df_rrs2),
    .io_id2df_rs2_d(decode_io_id2df_rs2_d),
    .io_id2df_dst(decode_io_id2df_dst),
    .io_id2df_dst_d(decode_io_id2df_dst_d),
    .io_id2df_jmp_type(decode_io_id2df_jmp_type),
    .io_id2df_special(decode_io_id2df_special),
    .io_id2df_swap(decode_io_id2df_swap),
    .io_id2df_indi(decode_io_id2df_indi),
    .io_id2df_drop(decode_io_id2df_drop),
    .io_id2df_stall(decode_io_id2df_stall),
    .io_id2df_recov(decode_io_id2df_recov),
    .io_id2df_valid(decode_io_id2df_valid),
    .io_id2df_ready(decode_io_id2df_ready),
    .io_idState_priv(decode_io_idState_priv)
  );
  Forwarding forwading ( // @[playground/src/noop/cpu.scala 98:29]
    .clock(forwading_clock),
    .reset(forwading_reset),
    .io_id2df_inst(forwading_io_id2df_inst),
    .io_id2df_pc(forwading_io_id2df_pc),
    .io_id2df_excep_cause(forwading_io_id2df_excep_cause),
    .io_id2df_excep_tval(forwading_io_id2df_excep_tval),
    .io_id2df_excep_en(forwading_io_id2df_excep_en),
    .io_id2df_excep_pc(forwading_io_id2df_excep_pc),
    .io_id2df_excep_etype(forwading_io_id2df_excep_etype),
    .io_id2df_ctrl_aluOp(forwading_io_id2df_ctrl_aluOp),
    .io_id2df_ctrl_aluWidth(forwading_io_id2df_ctrl_aluWidth),
    .io_id2df_ctrl_dcMode(forwading_io_id2df_ctrl_dcMode),
    .io_id2df_ctrl_writeRegEn(forwading_io_id2df_ctrl_writeRegEn),
    .io_id2df_ctrl_writeCSREn(forwading_io_id2df_ctrl_writeCSREn),
    .io_id2df_ctrl_brType(forwading_io_id2df_ctrl_brType),
    .io_id2df_rs1(forwading_io_id2df_rs1),
    .io_id2df_rrs1(forwading_io_id2df_rrs1),
    .io_id2df_rs1_d(forwading_io_id2df_rs1_d),
    .io_id2df_rs2(forwading_io_id2df_rs2),
    .io_id2df_rrs2(forwading_io_id2df_rrs2),
    .io_id2df_rs2_d(forwading_io_id2df_rs2_d),
    .io_id2df_dst(forwading_io_id2df_dst),
    .io_id2df_dst_d(forwading_io_id2df_dst_d),
    .io_id2df_jmp_type(forwading_io_id2df_jmp_type),
    .io_id2df_special(forwading_io_id2df_special),
    .io_id2df_swap(forwading_io_id2df_swap),
    .io_id2df_indi(forwading_io_id2df_indi),
    .io_id2df_drop(forwading_io_id2df_drop),
    .io_id2df_stall(forwading_io_id2df_stall),
    .io_id2df_recov(forwading_io_id2df_recov),
    .io_id2df_valid(forwading_io_id2df_valid),
    .io_id2df_ready(forwading_io_id2df_ready),
    .io_df2rr_inst(forwading_io_df2rr_inst),
    .io_df2rr_pc(forwading_io_df2rr_pc),
    .io_df2rr_excep_cause(forwading_io_df2rr_excep_cause),
    .io_df2rr_excep_tval(forwading_io_df2rr_excep_tval),
    .io_df2rr_excep_en(forwading_io_df2rr_excep_en),
    .io_df2rr_excep_pc(forwading_io_df2rr_excep_pc),
    .io_df2rr_excep_etype(forwading_io_df2rr_excep_etype),
    .io_df2rr_ctrl_aluOp(forwading_io_df2rr_ctrl_aluOp),
    .io_df2rr_ctrl_aluWidth(forwading_io_df2rr_ctrl_aluWidth),
    .io_df2rr_ctrl_dcMode(forwading_io_df2rr_ctrl_dcMode),
    .io_df2rr_ctrl_writeRegEn(forwading_io_df2rr_ctrl_writeRegEn),
    .io_df2rr_ctrl_writeCSREn(forwading_io_df2rr_ctrl_writeCSREn),
    .io_df2rr_ctrl_brType(forwading_io_df2rr_ctrl_brType),
    .io_df2rr_rs1(forwading_io_df2rr_rs1),
    .io_df2rr_rrs1(forwading_io_df2rr_rrs1),
    .io_df2rr_rs1_d(forwading_io_df2rr_rs1_d),
    .io_df2rr_rs2(forwading_io_df2rr_rs2),
    .io_df2rr_rrs2(forwading_io_df2rr_rrs2),
    .io_df2rr_rs2_d(forwading_io_df2rr_rs2_d),
    .io_df2rr_dst(forwading_io_df2rr_dst),
    .io_df2rr_dst_d(forwading_io_df2rr_dst_d),
    .io_df2rr_jmp_type(forwading_io_df2rr_jmp_type),
    .io_df2rr_special(forwading_io_df2rr_special),
    .io_df2rr_swap(forwading_io_df2rr_swap),
    .io_df2rr_indi(forwading_io_df2rr_indi),
    .io_df2rr_drop(forwading_io_df2rr_drop),
    .io_df2rr_stall(forwading_io_df2rr_stall),
    .io_df2rr_recov(forwading_io_df2rr_recov),
    .io_df2rr_valid(forwading_io_df2rr_valid),
    .io_df2rr_ready(forwading_io_df2rr_ready),
    .io_d_rr_id(forwading_io_d_rr_id),
    .io_d_rr_data(forwading_io_d_rr_data),
    .io_d_rr_state(forwading_io_d_rr_state),
    .io_d_ex_id(forwading_io_d_ex_id),
    .io_d_ex_data(forwading_io_d_ex_data),
    .io_d_ex_state(forwading_io_d_ex_state),
    .io_d_mem1_id(forwading_io_d_mem1_id),
    .io_d_mem1_data(forwading_io_d_mem1_data),
    .io_d_mem1_state(forwading_io_d_mem1_state),
    .io_d_mem2_id(forwading_io_d_mem2_id),
    .io_d_mem2_data(forwading_io_d_mem2_data),
    .io_d_mem2_state(forwading_io_d_mem2_state),
    .io_d_mem3_id(forwading_io_d_mem3_id),
    .io_d_mem3_data(forwading_io_d_mem3_data),
    .io_d_mem3_state(forwading_io_d_mem3_state)
  );
  ReadRegs readregs ( // @[playground/src/noop/cpu.scala 99:29]
    .clock(readregs_clock),
    .reset(readregs_reset),
    .io_df2rr_inst(readregs_io_df2rr_inst),
    .io_df2rr_pc(readregs_io_df2rr_pc),
    .io_df2rr_excep_cause(readregs_io_df2rr_excep_cause),
    .io_df2rr_excep_tval(readregs_io_df2rr_excep_tval),
    .io_df2rr_excep_en(readregs_io_df2rr_excep_en),
    .io_df2rr_excep_pc(readregs_io_df2rr_excep_pc),
    .io_df2rr_excep_etype(readregs_io_df2rr_excep_etype),
    .io_df2rr_ctrl_aluOp(readregs_io_df2rr_ctrl_aluOp),
    .io_df2rr_ctrl_aluWidth(readregs_io_df2rr_ctrl_aluWidth),
    .io_df2rr_ctrl_dcMode(readregs_io_df2rr_ctrl_dcMode),
    .io_df2rr_ctrl_writeRegEn(readregs_io_df2rr_ctrl_writeRegEn),
    .io_df2rr_ctrl_writeCSREn(readregs_io_df2rr_ctrl_writeCSREn),
    .io_df2rr_ctrl_brType(readregs_io_df2rr_ctrl_brType),
    .io_df2rr_rs1(readregs_io_df2rr_rs1),
    .io_df2rr_rrs1(readregs_io_df2rr_rrs1),
    .io_df2rr_rs1_d(readregs_io_df2rr_rs1_d),
    .io_df2rr_rs2(readregs_io_df2rr_rs2),
    .io_df2rr_rrs2(readregs_io_df2rr_rrs2),
    .io_df2rr_rs2_d(readregs_io_df2rr_rs2_d),
    .io_df2rr_dst(readregs_io_df2rr_dst),
    .io_df2rr_dst_d(readregs_io_df2rr_dst_d),
    .io_df2rr_jmp_type(readregs_io_df2rr_jmp_type),
    .io_df2rr_special(readregs_io_df2rr_special),
    .io_df2rr_swap(readregs_io_df2rr_swap),
    .io_df2rr_indi(readregs_io_df2rr_indi),
    .io_df2rr_drop(readregs_io_df2rr_drop),
    .io_df2rr_stall(readregs_io_df2rr_stall),
    .io_df2rr_recov(readregs_io_df2rr_recov),
    .io_df2rr_valid(readregs_io_df2rr_valid),
    .io_df2rr_ready(readregs_io_df2rr_ready),
    .io_rr2ex_inst(readregs_io_rr2ex_inst),
    .io_rr2ex_pc(readregs_io_rr2ex_pc),
    .io_rr2ex_excep_cause(readregs_io_rr2ex_excep_cause),
    .io_rr2ex_excep_tval(readregs_io_rr2ex_excep_tval),
    .io_rr2ex_excep_en(readregs_io_rr2ex_excep_en),
    .io_rr2ex_excep_pc(readregs_io_rr2ex_excep_pc),
    .io_rr2ex_excep_etype(readregs_io_rr2ex_excep_etype),
    .io_rr2ex_ctrl_aluOp(readregs_io_rr2ex_ctrl_aluOp),
    .io_rr2ex_ctrl_aluWidth(readregs_io_rr2ex_ctrl_aluWidth),
    .io_rr2ex_ctrl_dcMode(readregs_io_rr2ex_ctrl_dcMode),
    .io_rr2ex_ctrl_writeRegEn(readregs_io_rr2ex_ctrl_writeRegEn),
    .io_rr2ex_ctrl_writeCSREn(readregs_io_rr2ex_ctrl_writeCSREn),
    .io_rr2ex_ctrl_brType(readregs_io_rr2ex_ctrl_brType),
    .io_rr2ex_rs1_d(readregs_io_rr2ex_rs1_d),
    .io_rr2ex_rs2(readregs_io_rr2ex_rs2),
    .io_rr2ex_rs2_d(readregs_io_rr2ex_rs2_d),
    .io_rr2ex_dst(readregs_io_rr2ex_dst),
    .io_rr2ex_dst_d(readregs_io_rr2ex_dst_d),
    .io_rr2ex_rcsr_id(readregs_io_rr2ex_rcsr_id),
    .io_rr2ex_jmp_type(readregs_io_rr2ex_jmp_type),
    .io_rr2ex_special(readregs_io_rr2ex_special),
    .io_rr2ex_indi(readregs_io_rr2ex_indi),
    .io_rr2ex_drop(readregs_io_rr2ex_drop),
    .io_rr2ex_stall(readregs_io_rr2ex_stall),
    .io_rr2ex_recov(readregs_io_rr2ex_recov),
    .io_rr2ex_valid(readregs_io_rr2ex_valid),
    .io_rr2ex_ready(readregs_io_rr2ex_ready),
    .io_rs1Read_id(readregs_io_rs1Read_id),
    .io_rs1Read_data(readregs_io_rs1Read_data),
    .io_rs2Read_id(readregs_io_rs2Read_id),
    .io_rs2Read_data(readregs_io_rs2Read_data),
    .io_csrRead_id(readregs_io_csrRead_id),
    .io_csrRead_data(readregs_io_csrRead_data),
    .io_csrRead_is_err(readregs_io_csrRead_is_err),
    .io_d_rr_id(readregs_io_d_rr_id),
    .io_d_rr_data(readregs_io_d_rr_data),
    .io_d_rr_state(readregs_io_d_rr_state)
  );
  Execute execute ( // @[playground/src/noop/cpu.scala 100:29]
    .clock(execute_clock),
    .reset(execute_reset),
    .io_rr2ex_inst(execute_io_rr2ex_inst),
    .io_rr2ex_pc(execute_io_rr2ex_pc),
    .io_rr2ex_excep_cause(execute_io_rr2ex_excep_cause),
    .io_rr2ex_excep_tval(execute_io_rr2ex_excep_tval),
    .io_rr2ex_excep_en(execute_io_rr2ex_excep_en),
    .io_rr2ex_excep_pc(execute_io_rr2ex_excep_pc),
    .io_rr2ex_excep_etype(execute_io_rr2ex_excep_etype),
    .io_rr2ex_ctrl_aluOp(execute_io_rr2ex_ctrl_aluOp),
    .io_rr2ex_ctrl_aluWidth(execute_io_rr2ex_ctrl_aluWidth),
    .io_rr2ex_ctrl_dcMode(execute_io_rr2ex_ctrl_dcMode),
    .io_rr2ex_ctrl_writeRegEn(execute_io_rr2ex_ctrl_writeRegEn),
    .io_rr2ex_ctrl_writeCSREn(execute_io_rr2ex_ctrl_writeCSREn),
    .io_rr2ex_ctrl_brType(execute_io_rr2ex_ctrl_brType),
    .io_rr2ex_rs1_d(execute_io_rr2ex_rs1_d),
    .io_rr2ex_rs2(execute_io_rr2ex_rs2),
    .io_rr2ex_rs2_d(execute_io_rr2ex_rs2_d),
    .io_rr2ex_dst(execute_io_rr2ex_dst),
    .io_rr2ex_dst_d(execute_io_rr2ex_dst_d),
    .io_rr2ex_rcsr_id(execute_io_rr2ex_rcsr_id),
    .io_rr2ex_jmp_type(execute_io_rr2ex_jmp_type),
    .io_rr2ex_special(execute_io_rr2ex_special),
    .io_rr2ex_indi(execute_io_rr2ex_indi),
    .io_rr2ex_drop(execute_io_rr2ex_drop),
    .io_rr2ex_stall(execute_io_rr2ex_stall),
    .io_rr2ex_recov(execute_io_rr2ex_recov),
    .io_rr2ex_valid(execute_io_rr2ex_valid),
    .io_rr2ex_ready(execute_io_rr2ex_ready),
    .io_ex2mem_inst(execute_io_ex2mem_inst),
    .io_ex2mem_pc(execute_io_ex2mem_pc),
    .io_ex2mem_excep_cause(execute_io_ex2mem_excep_cause),
    .io_ex2mem_excep_tval(execute_io_ex2mem_excep_tval),
    .io_ex2mem_excep_en(execute_io_ex2mem_excep_en),
    .io_ex2mem_excep_pc(execute_io_ex2mem_excep_pc),
    .io_ex2mem_excep_etype(execute_io_ex2mem_excep_etype),
    .io_ex2mem_ctrl_dcMode(execute_io_ex2mem_ctrl_dcMode),
    .io_ex2mem_ctrl_writeRegEn(execute_io_ex2mem_ctrl_writeRegEn),
    .io_ex2mem_ctrl_writeCSREn(execute_io_ex2mem_ctrl_writeCSREn),
    .io_ex2mem_mem_addr(execute_io_ex2mem_mem_addr),
    .io_ex2mem_mem_data(execute_io_ex2mem_mem_data),
    .io_ex2mem_csr_id(execute_io_ex2mem_csr_id),
    .io_ex2mem_csr_d(execute_io_ex2mem_csr_d),
    .io_ex2mem_dst(execute_io_ex2mem_dst),
    .io_ex2mem_dst_d(execute_io_ex2mem_dst_d),
    .io_ex2mem_rcsr_id(execute_io_ex2mem_rcsr_id),
    .io_ex2mem_special(execute_io_ex2mem_special),
    .io_ex2mem_indi(execute_io_ex2mem_indi),
    .io_ex2mem_drop(execute_io_ex2mem_drop),
    .io_ex2mem_stall(execute_io_ex2mem_stall),
    .io_ex2mem_recov(execute_io_ex2mem_recov),
    .io_ex2mem_valid(execute_io_ex2mem_valid),
    .io_ex2mem_ready(execute_io_ex2mem_ready),
    .io_d_ex_id(execute_io_d_ex_id),
    .io_d_ex_data(execute_io_d_ex_data),
    .io_d_ex_state(execute_io_d_ex_state),
    .io_ex2if_seq_pc(execute_io_ex2if_seq_pc),
    .io_ex2if_valid(execute_io_ex2if_valid),
    .io_updateNextPc_seq_pc(execute_io_updateNextPc_seq_pc),
    .io_updateNextPc_valid(execute_io_updateNextPc_valid)
  );
  Memory memory ( // @[playground/src/noop/cpu.scala 101:29]
    .clock(memory_clock),
    .reset(memory_reset),
    .io_ex2mem_inst(memory_io_ex2mem_inst),
    .io_ex2mem_pc(memory_io_ex2mem_pc),
    .io_ex2mem_excep_cause(memory_io_ex2mem_excep_cause),
    .io_ex2mem_excep_tval(memory_io_ex2mem_excep_tval),
    .io_ex2mem_excep_en(memory_io_ex2mem_excep_en),
    .io_ex2mem_excep_pc(memory_io_ex2mem_excep_pc),
    .io_ex2mem_excep_etype(memory_io_ex2mem_excep_etype),
    .io_ex2mem_ctrl_dcMode(memory_io_ex2mem_ctrl_dcMode),
    .io_ex2mem_ctrl_writeRegEn(memory_io_ex2mem_ctrl_writeRegEn),
    .io_ex2mem_ctrl_writeCSREn(memory_io_ex2mem_ctrl_writeCSREn),
    .io_ex2mem_mem_addr(memory_io_ex2mem_mem_addr),
    .io_ex2mem_mem_data(memory_io_ex2mem_mem_data),
    .io_ex2mem_csr_id(memory_io_ex2mem_csr_id),
    .io_ex2mem_csr_d(memory_io_ex2mem_csr_d),
    .io_ex2mem_dst(memory_io_ex2mem_dst),
    .io_ex2mem_dst_d(memory_io_ex2mem_dst_d),
    .io_ex2mem_rcsr_id(memory_io_ex2mem_rcsr_id),
    .io_ex2mem_special(memory_io_ex2mem_special),
    .io_ex2mem_indi(memory_io_ex2mem_indi),
    .io_ex2mem_drop(memory_io_ex2mem_drop),
    .io_ex2mem_stall(memory_io_ex2mem_stall),
    .io_ex2mem_recov(memory_io_ex2mem_recov),
    .io_ex2mem_valid(memory_io_ex2mem_valid),
    .io_ex2mem_ready(memory_io_ex2mem_ready),
    .io_mem2rb_inst(memory_io_mem2rb_inst),
    .io_mem2rb_pc(memory_io_mem2rb_pc),
    .io_mem2rb_excep_cause(memory_io_mem2rb_excep_cause),
    .io_mem2rb_excep_tval(memory_io_mem2rb_excep_tval),
    .io_mem2rb_excep_en(memory_io_mem2rb_excep_en),
    .io_mem2rb_excep_pc(memory_io_mem2rb_excep_pc),
    .io_mem2rb_excep_etype(memory_io_mem2rb_excep_etype),
    .io_mem2rb_csr_id(memory_io_mem2rb_csr_id),
    .io_mem2rb_csr_d(memory_io_mem2rb_csr_d),
    .io_mem2rb_csr_en(memory_io_mem2rb_csr_en),
    .io_mem2rb_dst(memory_io_mem2rb_dst),
    .io_mem2rb_dst_d(memory_io_mem2rb_dst_d),
    .io_mem2rb_dst_en(memory_io_mem2rb_dst_en),
    .io_mem2rb_rcsr_id(memory_io_mem2rb_rcsr_id),
    .io_mem2rb_special(memory_io_mem2rb_special),
    .io_mem2rb_is_mmio(memory_io_mem2rb_is_mmio),
    .io_mem2rb_drop(memory_io_mem2rb_drop),
    .io_mem2rb_stall(memory_io_mem2rb_stall),
    .io_mem2rb_recov(memory_io_mem2rb_recov),
    .io_mem2rb_valid(memory_io_mem2rb_valid),
    .io_mem2rb_ready(memory_io_mem2rb_ready),
    .io_dataRW_addr(memory_io_dataRW_addr),
    .io_dataRW_rdata(memory_io_dataRW_rdata),
    .io_dataRW_rvalid(memory_io_dataRW_rvalid),
    .io_dataRW_wdata(memory_io_dataRW_wdata),
    .io_dataRW_dc_mode(memory_io_dataRW_dc_mode),
    .io_dataRW_amo(memory_io_dataRW_amo),
    .io_dataRW_ready(memory_io_dataRW_ready),
    .io_va2pa_vaddr(memory_io_va2pa_vaddr),
    .io_va2pa_vvalid(memory_io_va2pa_vvalid),
    .io_va2pa_m_type(memory_io_va2pa_m_type),
    .io_va2pa_paddr(memory_io_va2pa_paddr),
    .io_va2pa_pvalid(memory_io_va2pa_pvalid),
    .io_va2pa_tlb_excep_cause(memory_io_va2pa_tlb_excep_cause),
    .io_va2pa_tlb_excep_tval(memory_io_va2pa_tlb_excep_tval),
    .io_va2pa_tlb_excep_en(memory_io_va2pa_tlb_excep_en),
    .io_d_mem1_id(memory_io_d_mem1_id),
    .io_d_mem1_data(memory_io_d_mem1_data),
    .io_d_mem1_state(memory_io_d_mem1_state),
    .io_d_mem2_id(memory_io_d_mem2_id),
    .io_d_mem2_data(memory_io_d_mem2_data),
    .io_d_mem2_state(memory_io_d_mem2_state),
    .io_d_mem3_id(memory_io_d_mem3_id),
    .io_d_mem3_data(memory_io_d_mem3_data),
    .io_d_mem3_state(memory_io_d_mem3_state)
  );
  Writeback writeback ( // @[playground/src/noop/cpu.scala 102:29]
    .clock(writeback_clock),
    .reset(writeback_reset),
    .io_mem2rb_inst(writeback_io_mem2rb_inst),
    .io_mem2rb_pc(writeback_io_mem2rb_pc),
    .io_mem2rb_excep_cause(writeback_io_mem2rb_excep_cause),
    .io_mem2rb_excep_tval(writeback_io_mem2rb_excep_tval),
    .io_mem2rb_excep_en(writeback_io_mem2rb_excep_en),
    .io_mem2rb_excep_pc(writeback_io_mem2rb_excep_pc),
    .io_mem2rb_excep_etype(writeback_io_mem2rb_excep_etype),
    .io_mem2rb_csr_id(writeback_io_mem2rb_csr_id),
    .io_mem2rb_csr_d(writeback_io_mem2rb_csr_d),
    .io_mem2rb_csr_en(writeback_io_mem2rb_csr_en),
    .io_mem2rb_dst(writeback_io_mem2rb_dst),
    .io_mem2rb_dst_d(writeback_io_mem2rb_dst_d),
    .io_mem2rb_dst_en(writeback_io_mem2rb_dst_en),
    .io_mem2rb_rcsr_id(writeback_io_mem2rb_rcsr_id),
    .io_mem2rb_special(writeback_io_mem2rb_special),
    .io_mem2rb_is_mmio(writeback_io_mem2rb_is_mmio),
    .io_mem2rb_drop(writeback_io_mem2rb_drop),
    .io_mem2rb_stall(writeback_io_mem2rb_stall),
    .io_mem2rb_recov(writeback_io_mem2rb_recov),
    .io_mem2rb_valid(writeback_io_mem2rb_valid),
    .io_mem2rb_ready(writeback_io_mem2rb_ready),
    .io_wReg_id(writeback_io_wReg_id),
    .io_wReg_data(writeback_io_wReg_data),
    .io_wReg_en(writeback_io_wReg_en),
    .io_wCsr_id(writeback_io_wCsr_id),
    .io_wCsr_data(writeback_io_wCsr_data),
    .io_wCsr_en(writeback_io_wCsr_en),
    .io_excep_cause(writeback_io_excep_cause),
    .io_excep_tval(writeback_io_excep_tval),
    .io_excep_en(writeback_io_excep_en),
    .io_excep_pc(writeback_io_excep_pc),
    .io_excep_etype(writeback_io_excep_etype),
    .io_wb2if_seq_pc(writeback_io_wb2if_seq_pc),
    .io_wb2if_valid(writeback_io_wb2if_valid),
    .io_recov(writeback_io_recov),
    .io_flush_tlb(writeback_io_flush_tlb),
    .io_flush_cache(writeback_io_flush_cache)
  );
  Regs regs ( // @[playground/src/noop/cpu.scala 104:29]
    .clock(regs_clock),
    .reset(regs_reset),
    .io_rs1_id(regs_io_rs1_id),
    .io_rs1_data(regs_io_rs1_data),
    .io_rs2_id(regs_io_rs2_id),
    .io_rs2_data(regs_io_rs2_data),
    .io_dst_id(regs_io_dst_id),
    .io_dst_data(regs_io_dst_data),
    .io_dst_en(regs_io_dst_en)
  );
  Csrs csrs ( // @[playground/src/noop/cpu.scala 105:29]
    .clock(csrs_clock),
    .reset(csrs_reset),
    .io_rs_id(csrs_io_rs_id),
    .io_rs_data(csrs_io_rs_data),
    .io_rs_is_err(csrs_io_rs_is_err),
    .io_rd_id(csrs_io_rd_id),
    .io_rd_data(csrs_io_rd_data),
    .io_rd_en(csrs_io_rd_en),
    .io_excep_cause(csrs_io_excep_cause),
    .io_excep_tval(csrs_io_excep_tval),
    .io_excep_en(csrs_io_excep_en),
    .io_excep_pc(csrs_io_excep_pc),
    .io_excep_etype(csrs_io_excep_etype),
    .io_mmuState_priv(csrs_io_mmuState_priv),
    .io_mmuState_mstatus(csrs_io_mmuState_mstatus),
    .io_mmuState_satp(csrs_io_mmuState_satp),
    .io_idState_priv(csrs_io_idState_priv),
    .io_reg2if_seq_pc(csrs_io_reg2if_seq_pc),
    .io_reg2if_valid(csrs_io_reg2if_valid),
    .io_intr_out_en(csrs_io_intr_out_en),
    .io_intr_out_cause(csrs_io_intr_out_cause),
    .io_clint_raise(csrs_io_clint_raise),
    .io_clint_clear(csrs_io_clint_clear),
    .io_plic_m_raise(csrs_io_plic_m_raise),
    .io_plic_m_clear(csrs_io_plic_m_clear),
    .io_plic_s_raise(csrs_io_plic_s_raise),
    .io_plic_s_clear(csrs_io_plic_s_clear),
    .io_updateNextPc_seq_pc(csrs_io_updateNextPc_seq_pc),
    .io_updateNextPc_valid(csrs_io_updateNextPc_valid),
    .io_intr_msip_raise(csrs_io_intr_msip_raise),
    .io_intr_msip_clear(csrs_io_intr_msip_clear)
  );
  InstCache icache ( // @[playground/src/noop/cpu.scala 106:29]
    .clock(icache_clock),
    .reset(icache_reset),
    .io_instAxi_ra_ready(icache_io_instAxi_ra_ready),
    .io_instAxi_ra_valid(icache_io_instAxi_ra_valid),
    .io_instAxi_ra_bits_addr(icache_io_instAxi_ra_bits_addr),
    .io_instAxi_rd_valid(icache_io_instAxi_rd_valid),
    .io_instAxi_rd_bits_data(icache_io_instAxi_rd_bits_data),
    .io_instAxi_rd_bits_last(icache_io_instAxi_rd_bits_last),
    .io_icRead_addr(icache_io_icRead_addr),
    .io_icRead_inst(icache_io_icRead_inst),
    .io_icRead_arvalid(icache_io_icRead_arvalid),
    .io_icRead_ready(icache_io_icRead_ready),
    .io_icRead_rvalid(icache_io_icRead_rvalid),
    .io_flush(icache_io_flush)
  );
  DataCache dcache ( // @[playground/src/noop/cpu.scala 107:29]
    .clock(dcache_clock),
    .reset(dcache_reset),
    .io_dataAxi_wa_ready(dcache_io_dataAxi_wa_ready),
    .io_dataAxi_wa_valid(dcache_io_dataAxi_wa_valid),
    .io_dataAxi_wa_bits_addr(dcache_io_dataAxi_wa_bits_addr),
    .io_dataAxi_wd_ready(dcache_io_dataAxi_wd_ready),
    .io_dataAxi_wd_valid(dcache_io_dataAxi_wd_valid),
    .io_dataAxi_wd_bits_data(dcache_io_dataAxi_wd_bits_data),
    .io_dataAxi_wd_bits_last(dcache_io_dataAxi_wd_bits_last),
    .io_dataAxi_ra_ready(dcache_io_dataAxi_ra_ready),
    .io_dataAxi_ra_valid(dcache_io_dataAxi_ra_valid),
    .io_dataAxi_ra_bits_addr(dcache_io_dataAxi_ra_bits_addr),
    .io_dataAxi_rd_valid(dcache_io_dataAxi_rd_valid),
    .io_dataAxi_rd_bits_data(dcache_io_dataAxi_rd_bits_data),
    .io_dataAxi_rd_bits_last(dcache_io_dataAxi_rd_bits_last),
    .io_dcRW_addr(dcache_io_dcRW_addr),
    .io_dcRW_rdata(dcache_io_dcRW_rdata),
    .io_dcRW_rvalid(dcache_io_dcRW_rvalid),
    .io_dcRW_wdata(dcache_io_dcRW_wdata),
    .io_dcRW_dc_mode(dcache_io_dcRW_dc_mode),
    .io_dcRW_amo(dcache_io_dcRW_amo),
    .io_dcRW_ready(dcache_io_dcRW_ready),
    .io_flush(dcache_io_flush),
    .io_flush_out(dcache_io_flush_out)
  );
  ToAXI mem2Axi ( // @[playground/src/noop/cpu.scala 109:29]
    .clock(mem2Axi_clock),
    .reset(mem2Axi_reset),
    .io_dataIO_addr(mem2Axi_io_dataIO_addr),
    .io_dataIO_rdata(mem2Axi_io_dataIO_rdata),
    .io_dataIO_rvalid(mem2Axi_io_dataIO_rvalid),
    .io_dataIO_wdata(mem2Axi_io_dataIO_wdata),
    .io_dataIO_dc_mode(mem2Axi_io_dataIO_dc_mode),
    .io_dataIO_ready(mem2Axi_io_dataIO_ready),
    .io_outAxi_wa_ready(mem2Axi_io_outAxi_wa_ready),
    .io_outAxi_wa_valid(mem2Axi_io_outAxi_wa_valid),
    .io_outAxi_wa_bits_id(mem2Axi_io_outAxi_wa_bits_id),
    .io_outAxi_wa_bits_addr(mem2Axi_io_outAxi_wa_bits_addr),
    .io_outAxi_wa_bits_len(mem2Axi_io_outAxi_wa_bits_len),
    .io_outAxi_wa_bits_size(mem2Axi_io_outAxi_wa_bits_size),
    .io_outAxi_wa_bits_burst(mem2Axi_io_outAxi_wa_bits_burst),
    .io_outAxi_wd_ready(mem2Axi_io_outAxi_wd_ready),
    .io_outAxi_wd_valid(mem2Axi_io_outAxi_wd_valid),
    .io_outAxi_wd_bits_data(mem2Axi_io_outAxi_wd_bits_data),
    .io_outAxi_wd_bits_strb(mem2Axi_io_outAxi_wd_bits_strb),
    .io_outAxi_wd_bits_last(mem2Axi_io_outAxi_wd_bits_last),
    .io_outAxi_wr_ready(mem2Axi_io_outAxi_wr_ready),
    .io_outAxi_wr_valid(mem2Axi_io_outAxi_wr_valid),
    .io_outAxi_wr_bits_id(mem2Axi_io_outAxi_wr_bits_id),
    .io_outAxi_wr_bits_resp(mem2Axi_io_outAxi_wr_bits_resp),
    .io_outAxi_ra_ready(mem2Axi_io_outAxi_ra_ready),
    .io_outAxi_ra_valid(mem2Axi_io_outAxi_ra_valid),
    .io_outAxi_ra_bits_id(mem2Axi_io_outAxi_ra_bits_id),
    .io_outAxi_ra_bits_addr(mem2Axi_io_outAxi_ra_bits_addr),
    .io_outAxi_ra_bits_len(mem2Axi_io_outAxi_ra_bits_len),
    .io_outAxi_ra_bits_size(mem2Axi_io_outAxi_ra_bits_size),
    .io_outAxi_ra_bits_burst(mem2Axi_io_outAxi_ra_bits_burst),
    .io_outAxi_rd_ready(mem2Axi_io_outAxi_rd_ready),
    .io_outAxi_rd_valid(mem2Axi_io_outAxi_rd_valid),
    .io_outAxi_rd_bits_id(mem2Axi_io_outAxi_rd_bits_id),
    .io_outAxi_rd_bits_data(mem2Axi_io_outAxi_rd_bits_data),
    .io_outAxi_rd_bits_resp(mem2Axi_io_outAxi_rd_bits_resp),
    .io_outAxi_rd_bits_last(mem2Axi_io_outAxi_rd_bits_last)
  );
  ToAXI flash2Axi ( // @[playground/src/noop/cpu.scala 110:29]
    .clock(flash2Axi_clock),
    .reset(flash2Axi_reset),
    .io_dataIO_addr(flash2Axi_io_dataIO_addr),
    .io_dataIO_rdata(flash2Axi_io_dataIO_rdata),
    .io_dataIO_rvalid(flash2Axi_io_dataIO_rvalid),
    .io_dataIO_wdata(flash2Axi_io_dataIO_wdata),
    .io_dataIO_dc_mode(flash2Axi_io_dataIO_dc_mode),
    .io_dataIO_ready(flash2Axi_io_dataIO_ready),
    .io_outAxi_wa_ready(flash2Axi_io_outAxi_wa_ready),
    .io_outAxi_wa_valid(flash2Axi_io_outAxi_wa_valid),
    .io_outAxi_wa_bits_id(flash2Axi_io_outAxi_wa_bits_id),
    .io_outAxi_wa_bits_addr(flash2Axi_io_outAxi_wa_bits_addr),
    .io_outAxi_wa_bits_len(flash2Axi_io_outAxi_wa_bits_len),
    .io_outAxi_wa_bits_size(flash2Axi_io_outAxi_wa_bits_size),
    .io_outAxi_wa_bits_burst(flash2Axi_io_outAxi_wa_bits_burst),
    .io_outAxi_wd_ready(flash2Axi_io_outAxi_wd_ready),
    .io_outAxi_wd_valid(flash2Axi_io_outAxi_wd_valid),
    .io_outAxi_wd_bits_data(flash2Axi_io_outAxi_wd_bits_data),
    .io_outAxi_wd_bits_strb(flash2Axi_io_outAxi_wd_bits_strb),
    .io_outAxi_wd_bits_last(flash2Axi_io_outAxi_wd_bits_last),
    .io_outAxi_wr_ready(flash2Axi_io_outAxi_wr_ready),
    .io_outAxi_wr_valid(flash2Axi_io_outAxi_wr_valid),
    .io_outAxi_wr_bits_id(flash2Axi_io_outAxi_wr_bits_id),
    .io_outAxi_wr_bits_resp(flash2Axi_io_outAxi_wr_bits_resp),
    .io_outAxi_ra_ready(flash2Axi_io_outAxi_ra_ready),
    .io_outAxi_ra_valid(flash2Axi_io_outAxi_ra_valid),
    .io_outAxi_ra_bits_id(flash2Axi_io_outAxi_ra_bits_id),
    .io_outAxi_ra_bits_addr(flash2Axi_io_outAxi_ra_bits_addr),
    .io_outAxi_ra_bits_len(flash2Axi_io_outAxi_ra_bits_len),
    .io_outAxi_ra_bits_size(flash2Axi_io_outAxi_ra_bits_size),
    .io_outAxi_ra_bits_burst(flash2Axi_io_outAxi_ra_bits_burst),
    .io_outAxi_rd_ready(flash2Axi_io_outAxi_rd_ready),
    .io_outAxi_rd_valid(flash2Axi_io_outAxi_rd_valid),
    .io_outAxi_rd_bits_id(flash2Axi_io_outAxi_rd_bits_id),
    .io_outAxi_rd_bits_data(flash2Axi_io_outAxi_rd_bits_data),
    .io_outAxi_rd_bits_resp(flash2Axi_io_outAxi_rd_bits_resp),
    .io_outAxi_rd_bits_last(flash2Axi_io_outAxi_rd_bits_last)
  );
  CrossBar crossBar ( // @[playground/src/noop/cpu.scala 112:29]
    .clock(crossBar_clock),
    .reset(crossBar_reset),
    .io_icAxi_ra_ready(crossBar_io_icAxi_ra_ready),
    .io_icAxi_ra_valid(crossBar_io_icAxi_ra_valid),
    .io_icAxi_ra_bits_addr(crossBar_io_icAxi_ra_bits_addr),
    .io_icAxi_rd_valid(crossBar_io_icAxi_rd_valid),
    .io_icAxi_rd_bits_data(crossBar_io_icAxi_rd_bits_data),
    .io_icAxi_rd_bits_last(crossBar_io_icAxi_rd_bits_last),
    .io_flashAxi_wa_ready(crossBar_io_flashAxi_wa_ready),
    .io_flashAxi_wa_valid(crossBar_io_flashAxi_wa_valid),
    .io_flashAxi_wa_bits_id(crossBar_io_flashAxi_wa_bits_id),
    .io_flashAxi_wa_bits_addr(crossBar_io_flashAxi_wa_bits_addr),
    .io_flashAxi_wa_bits_len(crossBar_io_flashAxi_wa_bits_len),
    .io_flashAxi_wa_bits_size(crossBar_io_flashAxi_wa_bits_size),
    .io_flashAxi_wa_bits_burst(crossBar_io_flashAxi_wa_bits_burst),
    .io_flashAxi_wd_ready(crossBar_io_flashAxi_wd_ready),
    .io_flashAxi_wd_valid(crossBar_io_flashAxi_wd_valid),
    .io_flashAxi_wd_bits_data(crossBar_io_flashAxi_wd_bits_data),
    .io_flashAxi_wd_bits_strb(crossBar_io_flashAxi_wd_bits_strb),
    .io_flashAxi_wd_bits_last(crossBar_io_flashAxi_wd_bits_last),
    .io_flashAxi_wr_ready(crossBar_io_flashAxi_wr_ready),
    .io_flashAxi_wr_valid(crossBar_io_flashAxi_wr_valid),
    .io_flashAxi_wr_bits_id(crossBar_io_flashAxi_wr_bits_id),
    .io_flashAxi_wr_bits_resp(crossBar_io_flashAxi_wr_bits_resp),
    .io_flashAxi_ra_ready(crossBar_io_flashAxi_ra_ready),
    .io_flashAxi_ra_valid(crossBar_io_flashAxi_ra_valid),
    .io_flashAxi_ra_bits_id(crossBar_io_flashAxi_ra_bits_id),
    .io_flashAxi_ra_bits_addr(crossBar_io_flashAxi_ra_bits_addr),
    .io_flashAxi_ra_bits_len(crossBar_io_flashAxi_ra_bits_len),
    .io_flashAxi_ra_bits_size(crossBar_io_flashAxi_ra_bits_size),
    .io_flashAxi_ra_bits_burst(crossBar_io_flashAxi_ra_bits_burst),
    .io_flashAxi_rd_ready(crossBar_io_flashAxi_rd_ready),
    .io_flashAxi_rd_valid(crossBar_io_flashAxi_rd_valid),
    .io_flashAxi_rd_bits_id(crossBar_io_flashAxi_rd_bits_id),
    .io_flashAxi_rd_bits_data(crossBar_io_flashAxi_rd_bits_data),
    .io_flashAxi_rd_bits_resp(crossBar_io_flashAxi_rd_bits_resp),
    .io_flashAxi_rd_bits_last(crossBar_io_flashAxi_rd_bits_last),
    .io_memAxi_wa_ready(crossBar_io_memAxi_wa_ready),
    .io_memAxi_wa_valid(crossBar_io_memAxi_wa_valid),
    .io_memAxi_wa_bits_addr(crossBar_io_memAxi_wa_bits_addr),
    .io_memAxi_wd_ready(crossBar_io_memAxi_wd_ready),
    .io_memAxi_wd_valid(crossBar_io_memAxi_wd_valid),
    .io_memAxi_wd_bits_data(crossBar_io_memAxi_wd_bits_data),
    .io_memAxi_wd_bits_last(crossBar_io_memAxi_wd_bits_last),
    .io_memAxi_ra_ready(crossBar_io_memAxi_ra_ready),
    .io_memAxi_ra_valid(crossBar_io_memAxi_ra_valid),
    .io_memAxi_ra_bits_addr(crossBar_io_memAxi_ra_bits_addr),
    .io_memAxi_rd_valid(crossBar_io_memAxi_rd_valid),
    .io_memAxi_rd_bits_data(crossBar_io_memAxi_rd_bits_data),
    .io_memAxi_rd_bits_last(crossBar_io_memAxi_rd_bits_last),
    .io_mmioAxi_wa_ready(crossBar_io_mmioAxi_wa_ready),
    .io_mmioAxi_wa_valid(crossBar_io_mmioAxi_wa_valid),
    .io_mmioAxi_wa_bits_id(crossBar_io_mmioAxi_wa_bits_id),
    .io_mmioAxi_wa_bits_addr(crossBar_io_mmioAxi_wa_bits_addr),
    .io_mmioAxi_wa_bits_len(crossBar_io_mmioAxi_wa_bits_len),
    .io_mmioAxi_wa_bits_size(crossBar_io_mmioAxi_wa_bits_size),
    .io_mmioAxi_wa_bits_burst(crossBar_io_mmioAxi_wa_bits_burst),
    .io_mmioAxi_wd_ready(crossBar_io_mmioAxi_wd_ready),
    .io_mmioAxi_wd_valid(crossBar_io_mmioAxi_wd_valid),
    .io_mmioAxi_wd_bits_data(crossBar_io_mmioAxi_wd_bits_data),
    .io_mmioAxi_wd_bits_strb(crossBar_io_mmioAxi_wd_bits_strb),
    .io_mmioAxi_wd_bits_last(crossBar_io_mmioAxi_wd_bits_last),
    .io_mmioAxi_wr_ready(crossBar_io_mmioAxi_wr_ready),
    .io_mmioAxi_wr_valid(crossBar_io_mmioAxi_wr_valid),
    .io_mmioAxi_wr_bits_id(crossBar_io_mmioAxi_wr_bits_id),
    .io_mmioAxi_wr_bits_resp(crossBar_io_mmioAxi_wr_bits_resp),
    .io_mmioAxi_ra_ready(crossBar_io_mmioAxi_ra_ready),
    .io_mmioAxi_ra_valid(crossBar_io_mmioAxi_ra_valid),
    .io_mmioAxi_ra_bits_id(crossBar_io_mmioAxi_ra_bits_id),
    .io_mmioAxi_ra_bits_addr(crossBar_io_mmioAxi_ra_bits_addr),
    .io_mmioAxi_ra_bits_len(crossBar_io_mmioAxi_ra_bits_len),
    .io_mmioAxi_ra_bits_size(crossBar_io_mmioAxi_ra_bits_size),
    .io_mmioAxi_ra_bits_burst(crossBar_io_mmioAxi_ra_bits_burst),
    .io_mmioAxi_rd_ready(crossBar_io_mmioAxi_rd_ready),
    .io_mmioAxi_rd_valid(crossBar_io_mmioAxi_rd_valid),
    .io_mmioAxi_rd_bits_id(crossBar_io_mmioAxi_rd_bits_id),
    .io_mmioAxi_rd_bits_data(crossBar_io_mmioAxi_rd_bits_data),
    .io_mmioAxi_rd_bits_resp(crossBar_io_mmioAxi_rd_bits_resp),
    .io_mmioAxi_rd_bits_last(crossBar_io_mmioAxi_rd_bits_last),
    .io_outAxi_wa_ready(crossBar_io_outAxi_wa_ready),
    .io_outAxi_wa_valid(crossBar_io_outAxi_wa_valid),
    .io_outAxi_wa_bits_id(crossBar_io_outAxi_wa_bits_id),
    .io_outAxi_wa_bits_addr(crossBar_io_outAxi_wa_bits_addr),
    .io_outAxi_wa_bits_len(crossBar_io_outAxi_wa_bits_len),
    .io_outAxi_wa_bits_size(crossBar_io_outAxi_wa_bits_size),
    .io_outAxi_wa_bits_burst(crossBar_io_outAxi_wa_bits_burst),
    .io_outAxi_wd_ready(crossBar_io_outAxi_wd_ready),
    .io_outAxi_wd_valid(crossBar_io_outAxi_wd_valid),
    .io_outAxi_wd_bits_data(crossBar_io_outAxi_wd_bits_data),
    .io_outAxi_wd_bits_strb(crossBar_io_outAxi_wd_bits_strb),
    .io_outAxi_wd_bits_last(crossBar_io_outAxi_wd_bits_last),
    .io_outAxi_wr_ready(crossBar_io_outAxi_wr_ready),
    .io_outAxi_wr_valid(crossBar_io_outAxi_wr_valid),
    .io_outAxi_wr_bits_id(crossBar_io_outAxi_wr_bits_id),
    .io_outAxi_wr_bits_resp(crossBar_io_outAxi_wr_bits_resp),
    .io_outAxi_ra_ready(crossBar_io_outAxi_ra_ready),
    .io_outAxi_ra_valid(crossBar_io_outAxi_ra_valid),
    .io_outAxi_ra_bits_id(crossBar_io_outAxi_ra_bits_id),
    .io_outAxi_ra_bits_addr(crossBar_io_outAxi_ra_bits_addr),
    .io_outAxi_ra_bits_len(crossBar_io_outAxi_ra_bits_len),
    .io_outAxi_ra_bits_size(crossBar_io_outAxi_ra_bits_size),
    .io_outAxi_ra_bits_burst(crossBar_io_outAxi_ra_bits_burst),
    .io_outAxi_rd_ready(crossBar_io_outAxi_rd_ready),
    .io_outAxi_rd_valid(crossBar_io_outAxi_rd_valid),
    .io_outAxi_rd_bits_id(crossBar_io_outAxi_rd_bits_id),
    .io_outAxi_rd_bits_data(crossBar_io_outAxi_rd_bits_data),
    .io_outAxi_rd_bits_resp(crossBar_io_outAxi_rd_bits_resp),
    .io_outAxi_rd_bits_last(crossBar_io_outAxi_rd_bits_last),
    .io_selectMem(crossBar_io_selectMem)
  );
  FetchCrossBar fetchCrossbar ( // @[playground/src/noop/cpu.scala 113:31]
    .clock(fetchCrossbar_clock),
    .reset(fetchCrossbar_reset),
    .io_instIO_addr(fetchCrossbar_io_instIO_addr),
    .io_instIO_inst(fetchCrossbar_io_instIO_inst),
    .io_instIO_arvalid(fetchCrossbar_io_instIO_arvalid),
    .io_instIO_rvalid(fetchCrossbar_io_instIO_rvalid),
    .io_icRead_addr(fetchCrossbar_io_icRead_addr),
    .io_icRead_inst(fetchCrossbar_io_icRead_inst),
    .io_icRead_arvalid(fetchCrossbar_io_icRead_arvalid),
    .io_icRead_rvalid(fetchCrossbar_io_icRead_rvalid),
    .io_flashRead_addr(fetchCrossbar_io_flashRead_addr),
    .io_flashRead_rdata(fetchCrossbar_io_flashRead_rdata),
    .io_flashRead_rvalid(fetchCrossbar_io_flashRead_rvalid),
    .io_flashRead_dc_mode(fetchCrossbar_io_flashRead_dc_mode)
  );
  Splite64to32 split64to32 ( // @[playground/src/noop/cpu.scala 114:29]
    .clock(split64to32_clock),
    .reset(split64to32_reset),
    .io_data_in_addr(split64to32_io_data_in_addr),
    .io_data_in_rdata(split64to32_io_data_in_rdata),
    .io_data_in_rvalid(split64to32_io_data_in_rvalid),
    .io_data_in_dc_mode(split64to32_io_data_in_dc_mode),
    .io_data_out_addr(split64to32_io_data_out_addr),
    .io_data_out_rdata(split64to32_io_data_out_rdata),
    .io_data_out_rvalid(split64to32_io_data_out_rvalid),
    .io_data_out_dc_mode(split64to32_io_data_out_dc_mode),
    .io_data_out_ready(split64to32_io_data_out_ready)
  );
  MemCrossBar memCrossbar ( // @[playground/src/noop/cpu.scala 115:29]
    .clock(memCrossbar_clock),
    .reset(memCrossbar_reset),
    .io_dataRW_addr(memCrossbar_io_dataRW_addr),
    .io_dataRW_rdata(memCrossbar_io_dataRW_rdata),
    .io_dataRW_rvalid(memCrossbar_io_dataRW_rvalid),
    .io_dataRW_wdata(memCrossbar_io_dataRW_wdata),
    .io_dataRW_dc_mode(memCrossbar_io_dataRW_dc_mode),
    .io_dataRW_amo(memCrossbar_io_dataRW_amo),
    .io_dataRW_ready(memCrossbar_io_dataRW_ready),
    .io_mmio_addr(memCrossbar_io_mmio_addr),
    .io_mmio_rdata(memCrossbar_io_mmio_rdata),
    .io_mmio_rvalid(memCrossbar_io_mmio_rvalid),
    .io_mmio_wdata(memCrossbar_io_mmio_wdata),
    .io_mmio_dc_mode(memCrossbar_io_mmio_dc_mode),
    .io_mmio_ready(memCrossbar_io_mmio_ready),
    .io_dcRW_addr(memCrossbar_io_dcRW_addr),
    .io_dcRW_rdata(memCrossbar_io_dcRW_rdata),
    .io_dcRW_rvalid(memCrossbar_io_dcRW_rvalid),
    .io_dcRW_wdata(memCrossbar_io_dcRW_wdata),
    .io_dcRW_dc_mode(memCrossbar_io_dcRW_dc_mode),
    .io_dcRW_amo(memCrossbar_io_dcRW_amo),
    .io_dcRW_ready(memCrossbar_io_dcRW_ready),
    .io_clintIO_addr(memCrossbar_io_clintIO_addr),
    .io_clintIO_rdata(memCrossbar_io_clintIO_rdata),
    .io_clintIO_wdata(memCrossbar_io_clintIO_wdata),
    .io_clintIO_wvalid(memCrossbar_io_clintIO_wvalid),
    .io_plicIO_addr(memCrossbar_io_plicIO_addr),
    .io_plicIO_rdata(memCrossbar_io_plicIO_rdata),
    .io_plicIO_wdata(memCrossbar_io_plicIO_wdata),
    .io_plicIO_wvalid(memCrossbar_io_plicIO_wvalid),
    .io_plicIO_arvalid(memCrossbar_io_plicIO_arvalid)
  );
  TLB tlb_if ( // @[playground/src/noop/cpu.scala 116:30]
    .clock(tlb_if_clock),
    .reset(tlb_if_reset),
    .io_va2pa_vaddr(tlb_if_io_va2pa_vaddr),
    .io_va2pa_vvalid(tlb_if_io_va2pa_vvalid),
    .io_va2pa_ready(tlb_if_io_va2pa_ready),
    .io_va2pa_paddr(tlb_if_io_va2pa_paddr),
    .io_va2pa_pvalid(tlb_if_io_va2pa_pvalid),
    .io_va2pa_tlb_excep_cause(tlb_if_io_va2pa_tlb_excep_cause),
    .io_va2pa_tlb_excep_tval(tlb_if_io_va2pa_tlb_excep_tval),
    .io_va2pa_tlb_excep_en(tlb_if_io_va2pa_tlb_excep_en),
    .io_mmuState_priv(tlb_if_io_mmuState_priv),
    .io_mmuState_mstatus(tlb_if_io_mmuState_mstatus),
    .io_mmuState_satp(tlb_if_io_mmuState_satp),
    .io_flush(tlb_if_io_flush),
    .io_dcacheRW_addr(tlb_if_io_dcacheRW_addr),
    .io_dcacheRW_rdata(tlb_if_io_dcacheRW_rdata),
    .io_dcacheRW_rvalid(tlb_if_io_dcacheRW_rvalid),
    .io_dcacheRW_wdata(tlb_if_io_dcacheRW_wdata),
    .io_dcacheRW_dc_mode(tlb_if_io_dcacheRW_dc_mode),
    .io_dcacheRW_ready(tlb_if_io_dcacheRW_ready)
  );
  TLB_1 tlb_mem ( // @[playground/src/noop/cpu.scala 117:30]
    .clock(tlb_mem_clock),
    .reset(tlb_mem_reset),
    .io_va2pa_vaddr(tlb_mem_io_va2pa_vaddr),
    .io_va2pa_vvalid(tlb_mem_io_va2pa_vvalid),
    .io_va2pa_m_type(tlb_mem_io_va2pa_m_type),
    .io_va2pa_ready(tlb_mem_io_va2pa_ready),
    .io_va2pa_paddr(tlb_mem_io_va2pa_paddr),
    .io_va2pa_pvalid(tlb_mem_io_va2pa_pvalid),
    .io_va2pa_tlb_excep_cause(tlb_mem_io_va2pa_tlb_excep_cause),
    .io_va2pa_tlb_excep_tval(tlb_mem_io_va2pa_tlb_excep_tval),
    .io_va2pa_tlb_excep_en(tlb_mem_io_va2pa_tlb_excep_en),
    .io_mmuState_priv(tlb_mem_io_mmuState_priv),
    .io_mmuState_mstatus(tlb_mem_io_mmuState_mstatus),
    .io_mmuState_satp(tlb_mem_io_mmuState_satp),
    .io_flush(tlb_mem_io_flush),
    .io_dcacheRW_addr(tlb_mem_io_dcacheRW_addr),
    .io_dcacheRW_rdata(tlb_mem_io_dcacheRW_rdata),
    .io_dcacheRW_rvalid(tlb_mem_io_dcacheRW_rvalid),
    .io_dcacheRW_wdata(tlb_mem_io_dcacheRW_wdata),
    .io_dcacheRW_dc_mode(tlb_mem_io_dcacheRW_dc_mode),
    .io_dcacheRW_ready(tlb_mem_io_dcacheRW_ready)
  );
  DcacheSelector dcSelector ( // @[playground/src/noop/cpu.scala 118:29]
    .clock(dcSelector_clock),
    .reset(dcSelector_reset),
    .io_tlb_if2dc_addr(dcSelector_io_tlb_if2dc_addr),
    .io_tlb_if2dc_rdata(dcSelector_io_tlb_if2dc_rdata),
    .io_tlb_if2dc_rvalid(dcSelector_io_tlb_if2dc_rvalid),
    .io_tlb_if2dc_wdata(dcSelector_io_tlb_if2dc_wdata),
    .io_tlb_if2dc_dc_mode(dcSelector_io_tlb_if2dc_dc_mode),
    .io_tlb_if2dc_ready(dcSelector_io_tlb_if2dc_ready),
    .io_tlb_mem2dc_addr(dcSelector_io_tlb_mem2dc_addr),
    .io_tlb_mem2dc_rdata(dcSelector_io_tlb_mem2dc_rdata),
    .io_tlb_mem2dc_rvalid(dcSelector_io_tlb_mem2dc_rvalid),
    .io_tlb_mem2dc_wdata(dcSelector_io_tlb_mem2dc_wdata),
    .io_tlb_mem2dc_dc_mode(dcSelector_io_tlb_mem2dc_dc_mode),
    .io_tlb_mem2dc_ready(dcSelector_io_tlb_mem2dc_ready),
    .io_mem2dc_addr(dcSelector_io_mem2dc_addr),
    .io_mem2dc_rdata(dcSelector_io_mem2dc_rdata),
    .io_mem2dc_rvalid(dcSelector_io_mem2dc_rvalid),
    .io_mem2dc_wdata(dcSelector_io_mem2dc_wdata),
    .io_mem2dc_dc_mode(dcSelector_io_mem2dc_dc_mode),
    .io_mem2dc_amo(dcSelector_io_mem2dc_amo),
    .io_mem2dc_ready(dcSelector_io_mem2dc_ready),
    .io_dma2dc_addr(dcSelector_io_dma2dc_addr),
    .io_dma2dc_rdata(dcSelector_io_dma2dc_rdata),
    .io_dma2dc_rvalid(dcSelector_io_dma2dc_rvalid),
    .io_dma2dc_wdata(dcSelector_io_dma2dc_wdata),
    .io_dma2dc_dc_mode(dcSelector_io_dma2dc_dc_mode),
    .io_dma2dc_ready(dcSelector_io_dma2dc_ready),
    .io_select_addr(dcSelector_io_select_addr),
    .io_select_rdata(dcSelector_io_select_rdata),
    .io_select_rvalid(dcSelector_io_select_rvalid),
    .io_select_wdata(dcSelector_io_select_wdata),
    .io_select_dc_mode(dcSelector_io_select_dc_mode),
    .io_select_amo(dcSelector_io_select_amo),
    .io_select_ready(dcSelector_io_select_ready)
  );
  CLINT clint ( // @[playground/src/noop/cpu.scala 119:29]
    .clock(clint_clock),
    .reset(clint_reset),
    .io_rw_addr(clint_io_rw_addr),
    .io_rw_rdata(clint_io_rw_rdata),
    .io_rw_wdata(clint_io_rw_wdata),
    .io_rw_wvalid(clint_io_rw_wvalid),
    .io_intr_raise(clint_io_intr_raise),
    .io_intr_clear(clint_io_intr_clear),
    .io_intr_msip_raise(clint_io_intr_msip_raise),
    .io_intr_msip_clear(clint_io_intr_msip_clear)
  );
  Plic plic ( // @[playground/src/noop/cpu.scala 120:29]
    .clock(plic_clock),
    .reset(plic_reset),
    .io_intr_in1(plic_io_intr_in1),
    .io_intr_out_m_raise(plic_io_intr_out_m_raise),
    .io_intr_out_m_clear(plic_io_intr_out_m_clear),
    .io_intr_out_s_raise(plic_io_intr_out_s_raise),
    .io_intr_out_s_clear(plic_io_intr_out_s_clear),
    .io_rw_addr(plic_io_rw_addr),
    .io_rw_rdata(plic_io_rw_rdata),
    .io_rw_wdata(plic_io_rw_wdata),
    .io_rw_wvalid(plic_io_rw_wvalid),
    .io_rw_arvalid(plic_io_rw_arvalid)
  );
  DmaBridge dmaBridge ( // @[playground/src/noop/cpu.scala 121:29]
    .clock(dmaBridge_clock),
    .reset(dmaBridge_reset),
    .io_dmaAxi_awready(dmaBridge_io_dmaAxi_awready),
    .io_dmaAxi_awvalid(dmaBridge_io_dmaAxi_awvalid),
    .io_dmaAxi_awaddr(dmaBridge_io_dmaAxi_awaddr),
    .io_dmaAxi_awid(dmaBridge_io_dmaAxi_awid),
    .io_dmaAxi_awlen(dmaBridge_io_dmaAxi_awlen),
    .io_dmaAxi_awsize(dmaBridge_io_dmaAxi_awsize),
    .io_dmaAxi_wready(dmaBridge_io_dmaAxi_wready),
    .io_dmaAxi_wvalid(dmaBridge_io_dmaAxi_wvalid),
    .io_dmaAxi_wdata(dmaBridge_io_dmaAxi_wdata),
    .io_dmaAxi_wstrb(dmaBridge_io_dmaAxi_wstrb),
    .io_dmaAxi_bready(dmaBridge_io_dmaAxi_bready),
    .io_dmaAxi_bvalid(dmaBridge_io_dmaAxi_bvalid),
    .io_dmaAxi_bid(dmaBridge_io_dmaAxi_bid),
    .io_dmaAxi_arready(dmaBridge_io_dmaAxi_arready),
    .io_dmaAxi_arvalid(dmaBridge_io_dmaAxi_arvalid),
    .io_dmaAxi_araddr(dmaBridge_io_dmaAxi_araddr),
    .io_dmaAxi_arid(dmaBridge_io_dmaAxi_arid),
    .io_dmaAxi_arlen(dmaBridge_io_dmaAxi_arlen),
    .io_dmaAxi_arsize(dmaBridge_io_dmaAxi_arsize),
    .io_dmaAxi_rready(dmaBridge_io_dmaAxi_rready),
    .io_dmaAxi_rvalid(dmaBridge_io_dmaAxi_rvalid),
    .io_dmaAxi_rdata(dmaBridge_io_dmaAxi_rdata),
    .io_dmaAxi_rlast(dmaBridge_io_dmaAxi_rlast),
    .io_dmaAxi_rid(dmaBridge_io_dmaAxi_rid),
    .io_dcRW_addr(dmaBridge_io_dcRW_addr),
    .io_dcRW_rdata(dmaBridge_io_dcRW_rdata),
    .io_dcRW_rvalid(dmaBridge_io_dcRW_rvalid),
    .io_dcRW_wdata(dmaBridge_io_dcRW_wdata),
    .io_dcRW_dc_mode(dmaBridge_io_dcRW_dc_mode),
    .io_dcRW_ready(dmaBridge_io_dcRW_ready)
  );
  assign io_master_awvalid = crossBar_io_outAxi_wa_valid; // @[playground/src/noop/cpu.scala 189:23]
  assign io_master_awaddr = crossBar_io_outAxi_wa_bits_addr; // @[playground/src/noop/cpu.scala 190:23]
  assign io_master_awid = crossBar_io_outAxi_wa_bits_id; // @[playground/src/noop/cpu.scala 191:23]
  assign io_master_awlen = crossBar_io_outAxi_wa_bits_len; // @[playground/src/noop/cpu.scala 192:23]
  assign io_master_awsize = crossBar_io_outAxi_wa_bits_size; // @[playground/src/noop/cpu.scala 193:23]
  assign io_master_awburst = crossBar_io_outAxi_wa_bits_burst; // @[playground/src/noop/cpu.scala 194:23]
  assign io_master_wvalid = crossBar_io_outAxi_wd_valid; // @[playground/src/noop/cpu.scala 197:23]
  assign io_master_wdata = crossBar_io_outAxi_wd_bits_data; // @[playground/src/noop/cpu.scala 198:23]
  assign io_master_wstrb = crossBar_io_outAxi_wd_bits_strb; // @[playground/src/noop/cpu.scala 199:23]
  assign io_master_wlast = crossBar_io_outAxi_wd_bits_last; // @[playground/src/noop/cpu.scala 200:23]
  assign io_master_bready = crossBar_io_outAxi_wr_ready; // @[playground/src/noop/cpu.scala 202:23]
  assign io_master_arvalid = crossBar_io_outAxi_ra_valid; // @[playground/src/noop/cpu.scala 208:23]
  assign io_master_araddr = crossBar_io_outAxi_ra_bits_addr; // @[playground/src/noop/cpu.scala 209:23]
  assign io_master_arid = crossBar_io_outAxi_ra_bits_id; // @[playground/src/noop/cpu.scala 210:23]
  assign io_master_arlen = crossBar_io_outAxi_ra_bits_len; // @[playground/src/noop/cpu.scala 211:23]
  assign io_master_arsize = crossBar_io_outAxi_ra_bits_size; // @[playground/src/noop/cpu.scala 212:23]
  assign io_master_arburst = crossBar_io_outAxi_ra_bits_burst; // @[playground/src/noop/cpu.scala 213:23]
  assign io_master_rready = crossBar_io_outAxi_rd_ready; // @[playground/src/noop/cpu.scala 215:23]
  assign io_slave_awready = dmaBridge_io_dmaAxi_awready; // @[playground/src/noop/cpu.scala 185:14]
  assign io_slave_wready = dmaBridge_io_dmaAxi_wready; // @[playground/src/noop/cpu.scala 185:14]
  assign io_slave_bvalid = dmaBridge_io_dmaAxi_bvalid; // @[playground/src/noop/cpu.scala 185:14]
  assign io_slave_bresp = 2'h0; // @[playground/src/noop/cpu.scala 185:14]
  assign io_slave_bid = dmaBridge_io_dmaAxi_bid; // @[playground/src/noop/cpu.scala 185:14]
  assign io_slave_arready = dmaBridge_io_dmaAxi_arready; // @[playground/src/noop/cpu.scala 185:14]
  assign io_slave_rvalid = dmaBridge_io_dmaAxi_rvalid; // @[playground/src/noop/cpu.scala 185:14]
  assign io_slave_rresp = 2'h0; // @[playground/src/noop/cpu.scala 185:14]
  assign io_slave_rdata = dmaBridge_io_dmaAxi_rdata; // @[playground/src/noop/cpu.scala 185:14]
  assign io_slave_rlast = dmaBridge_io_dmaAxi_rlast; // @[playground/src/noop/cpu.scala 185:14]
  assign io_slave_rid = dmaBridge_io_dmaAxi_rid; // @[playground/src/noop/cpu.scala 185:14]
  assign fetch_clock = clock;
  assign fetch_reset = reset;
  assign fetch_io_instRead_inst = fetchCrossbar_io_instIO_inst; // @[playground/src/noop/cpu.scala 123:25]
  assign fetch_io_instRead_rvalid = fetchCrossbar_io_instIO_rvalid; // @[playground/src/noop/cpu.scala 123:25]
  assign fetch_io_va2pa_paddr = tlb_if_io_va2pa_paddr; // @[playground/src/noop/cpu.scala 124:25]
  assign fetch_io_va2pa_pvalid = tlb_if_io_va2pa_pvalid; // @[playground/src/noop/cpu.scala 124:25]
  assign fetch_io_va2pa_tlb_excep_cause = tlb_if_io_va2pa_tlb_excep_cause; // @[playground/src/noop/cpu.scala 124:25]
  assign fetch_io_va2pa_tlb_excep_tval = tlb_if_io_va2pa_tlb_excep_tval; // @[playground/src/noop/cpu.scala 124:25]
  assign fetch_io_va2pa_tlb_excep_en = tlb_if_io_va2pa_tlb_excep_en; // @[playground/src/noop/cpu.scala 124:25]
  assign fetch_io_reg2if_seq_pc = csrs_io_reg2if_seq_pc; // @[playground/src/noop/cpu.scala 125:25]
  assign fetch_io_reg2if_valid = csrs_io_reg2if_valid; // @[playground/src/noop/cpu.scala 125:25]
  assign fetch_io_wb2if_seq_pc = writeback_io_wb2if_seq_pc; // @[playground/src/noop/cpu.scala 126:25]
  assign fetch_io_wb2if_valid = writeback_io_wb2if_valid; // @[playground/src/noop/cpu.scala 126:25]
  assign fetch_io_recov = writeback_io_recov; // @[playground/src/noop/cpu.scala 130:25]
  assign fetch_io_intr_in_en = csrs_io_intr_out_en; // @[playground/src/noop/cpu.scala 127:25]
  assign fetch_io_intr_in_cause = csrs_io_intr_out_cause; // @[playground/src/noop/cpu.scala 127:25]
  assign fetch_io_branchFail_seq_pc = execute_io_ex2if_seq_pc; // @[playground/src/noop/cpu.scala 128:25]
  assign fetch_io_branchFail_valid = execute_io_ex2if_valid; // @[playground/src/noop/cpu.scala 128:25]
  assign fetch_io_if2id_drop = decode_io_if2id_drop; // @[playground/src/noop/cpu.scala 129:25]
  assign fetch_io_if2id_stall = decode_io_if2id_stall; // @[playground/src/noop/cpu.scala 129:25]
  assign fetch_io_if2id_ready = decode_io_if2id_ready; // @[playground/src/noop/cpu.scala 129:25]
  assign decode_clock = clock;
  assign decode_reset = reset;
  assign decode_io_if2id_inst = fetch_io_if2id_inst; // @[playground/src/noop/cpu.scala 129:25]
  assign decode_io_if2id_pc = fetch_io_if2id_pc; // @[playground/src/noop/cpu.scala 129:25]
  assign decode_io_if2id_excep_cause = fetch_io_if2id_excep_cause; // @[playground/src/noop/cpu.scala 129:25]
  assign decode_io_if2id_excep_tval = fetch_io_if2id_excep_tval; // @[playground/src/noop/cpu.scala 129:25]
  assign decode_io_if2id_excep_en = fetch_io_if2id_excep_en; // @[playground/src/noop/cpu.scala 129:25]
  assign decode_io_if2id_excep_pc = fetch_io_if2id_excep_pc; // @[playground/src/noop/cpu.scala 129:25]
  assign decode_io_if2id_recov = fetch_io_if2id_recov; // @[playground/src/noop/cpu.scala 129:25]
  assign decode_io_if2id_valid = fetch_io_if2id_valid; // @[playground/src/noop/cpu.scala 129:25]
  assign decode_io_id2df_drop = forwading_io_id2df_drop; // @[playground/src/noop/cpu.scala 132:25]
  assign decode_io_id2df_stall = forwading_io_id2df_stall; // @[playground/src/noop/cpu.scala 132:25]
  assign decode_io_id2df_ready = forwading_io_id2df_ready; // @[playground/src/noop/cpu.scala 132:25]
  assign decode_io_idState_priv = csrs_io_idState_priv; // @[playground/src/noop/cpu.scala 133:25]
  assign forwading_clock = clock;
  assign forwading_reset = reset;
  assign forwading_io_id2df_inst = decode_io_id2df_inst; // @[playground/src/noop/cpu.scala 132:25]
  assign forwading_io_id2df_pc = decode_io_id2df_pc; // @[playground/src/noop/cpu.scala 132:25]
  assign forwading_io_id2df_excep_cause = decode_io_id2df_excep_cause; // @[playground/src/noop/cpu.scala 132:25]
  assign forwading_io_id2df_excep_tval = decode_io_id2df_excep_tval; // @[playground/src/noop/cpu.scala 132:25]
  assign forwading_io_id2df_excep_en = decode_io_id2df_excep_en; // @[playground/src/noop/cpu.scala 132:25]
  assign forwading_io_id2df_excep_pc = decode_io_id2df_excep_pc; // @[playground/src/noop/cpu.scala 132:25]
  assign forwading_io_id2df_excep_etype = decode_io_id2df_excep_etype; // @[playground/src/noop/cpu.scala 132:25]
  assign forwading_io_id2df_ctrl_aluOp = decode_io_id2df_ctrl_aluOp; // @[playground/src/noop/cpu.scala 132:25]
  assign forwading_io_id2df_ctrl_aluWidth = decode_io_id2df_ctrl_aluWidth; // @[playground/src/noop/cpu.scala 132:25]
  assign forwading_io_id2df_ctrl_dcMode = decode_io_id2df_ctrl_dcMode; // @[playground/src/noop/cpu.scala 132:25]
  assign forwading_io_id2df_ctrl_writeRegEn = decode_io_id2df_ctrl_writeRegEn; // @[playground/src/noop/cpu.scala 132:25]
  assign forwading_io_id2df_ctrl_writeCSREn = decode_io_id2df_ctrl_writeCSREn; // @[playground/src/noop/cpu.scala 132:25]
  assign forwading_io_id2df_ctrl_brType = decode_io_id2df_ctrl_brType; // @[playground/src/noop/cpu.scala 132:25]
  assign forwading_io_id2df_rs1 = decode_io_id2df_rs1; // @[playground/src/noop/cpu.scala 132:25]
  assign forwading_io_id2df_rrs1 = decode_io_id2df_rrs1; // @[playground/src/noop/cpu.scala 132:25]
  assign forwading_io_id2df_rs1_d = decode_io_id2df_rs1_d; // @[playground/src/noop/cpu.scala 132:25]
  assign forwading_io_id2df_rs2 = decode_io_id2df_rs2; // @[playground/src/noop/cpu.scala 132:25]
  assign forwading_io_id2df_rrs2 = decode_io_id2df_rrs2; // @[playground/src/noop/cpu.scala 132:25]
  assign forwading_io_id2df_rs2_d = decode_io_id2df_rs2_d; // @[playground/src/noop/cpu.scala 132:25]
  assign forwading_io_id2df_dst = decode_io_id2df_dst; // @[playground/src/noop/cpu.scala 132:25]
  assign forwading_io_id2df_dst_d = decode_io_id2df_dst_d; // @[playground/src/noop/cpu.scala 132:25]
  assign forwading_io_id2df_jmp_type = decode_io_id2df_jmp_type; // @[playground/src/noop/cpu.scala 132:25]
  assign forwading_io_id2df_special = decode_io_id2df_special; // @[playground/src/noop/cpu.scala 132:25]
  assign forwading_io_id2df_swap = decode_io_id2df_swap; // @[playground/src/noop/cpu.scala 132:25]
  assign forwading_io_id2df_indi = decode_io_id2df_indi; // @[playground/src/noop/cpu.scala 132:25]
  assign forwading_io_id2df_recov = decode_io_id2df_recov; // @[playground/src/noop/cpu.scala 132:25]
  assign forwading_io_id2df_valid = decode_io_id2df_valid; // @[playground/src/noop/cpu.scala 132:25]
  assign forwading_io_df2rr_drop = readregs_io_df2rr_drop; // @[playground/src/noop/cpu.scala 134:25]
  assign forwading_io_df2rr_stall = readregs_io_df2rr_stall; // @[playground/src/noop/cpu.scala 134:25]
  assign forwading_io_df2rr_ready = readregs_io_df2rr_ready; // @[playground/src/noop/cpu.scala 134:25]
  assign forwading_io_d_rr_id = readregs_io_d_rr_id; // @[playground/src/noop/cpu.scala 135:25]
  assign forwading_io_d_rr_data = readregs_io_d_rr_data; // @[playground/src/noop/cpu.scala 135:25]
  assign forwading_io_d_rr_state = readregs_io_d_rr_state; // @[playground/src/noop/cpu.scala 135:25]
  assign forwading_io_d_ex_id = execute_io_d_ex_id; // @[playground/src/noop/cpu.scala 136:25]
  assign forwading_io_d_ex_data = execute_io_d_ex_data; // @[playground/src/noop/cpu.scala 136:25]
  assign forwading_io_d_ex_state = execute_io_d_ex_state; // @[playground/src/noop/cpu.scala 136:25]
  assign forwading_io_d_mem1_id = memory_io_d_mem1_id; // @[playground/src/noop/cpu.scala 137:25]
  assign forwading_io_d_mem1_data = memory_io_d_mem1_data; // @[playground/src/noop/cpu.scala 137:25]
  assign forwading_io_d_mem1_state = memory_io_d_mem1_state; // @[playground/src/noop/cpu.scala 137:25]
  assign forwading_io_d_mem2_id = memory_io_d_mem2_id; // @[playground/src/noop/cpu.scala 138:25]
  assign forwading_io_d_mem2_data = memory_io_d_mem2_data; // @[playground/src/noop/cpu.scala 138:25]
  assign forwading_io_d_mem2_state = memory_io_d_mem2_state; // @[playground/src/noop/cpu.scala 138:25]
  assign forwading_io_d_mem3_id = memory_io_d_mem3_id; // @[playground/src/noop/cpu.scala 139:25]
  assign forwading_io_d_mem3_data = memory_io_d_mem3_data; // @[playground/src/noop/cpu.scala 139:25]
  assign forwading_io_d_mem3_state = memory_io_d_mem3_state; // @[playground/src/noop/cpu.scala 139:25]
  assign readregs_clock = clock;
  assign readregs_reset = reset;
  assign readregs_io_df2rr_inst = forwading_io_df2rr_inst; // @[playground/src/noop/cpu.scala 134:25]
  assign readregs_io_df2rr_pc = forwading_io_df2rr_pc; // @[playground/src/noop/cpu.scala 134:25]
  assign readregs_io_df2rr_excep_cause = forwading_io_df2rr_excep_cause; // @[playground/src/noop/cpu.scala 134:25]
  assign readregs_io_df2rr_excep_tval = forwading_io_df2rr_excep_tval; // @[playground/src/noop/cpu.scala 134:25]
  assign readregs_io_df2rr_excep_en = forwading_io_df2rr_excep_en; // @[playground/src/noop/cpu.scala 134:25]
  assign readregs_io_df2rr_excep_pc = forwading_io_df2rr_excep_pc; // @[playground/src/noop/cpu.scala 134:25]
  assign readregs_io_df2rr_excep_etype = forwading_io_df2rr_excep_etype; // @[playground/src/noop/cpu.scala 134:25]
  assign readregs_io_df2rr_ctrl_aluOp = forwading_io_df2rr_ctrl_aluOp; // @[playground/src/noop/cpu.scala 134:25]
  assign readregs_io_df2rr_ctrl_aluWidth = forwading_io_df2rr_ctrl_aluWidth; // @[playground/src/noop/cpu.scala 134:25]
  assign readregs_io_df2rr_ctrl_dcMode = forwading_io_df2rr_ctrl_dcMode; // @[playground/src/noop/cpu.scala 134:25]
  assign readregs_io_df2rr_ctrl_writeRegEn = forwading_io_df2rr_ctrl_writeRegEn; // @[playground/src/noop/cpu.scala 134:25]
  assign readregs_io_df2rr_ctrl_writeCSREn = forwading_io_df2rr_ctrl_writeCSREn; // @[playground/src/noop/cpu.scala 134:25]
  assign readregs_io_df2rr_ctrl_brType = forwading_io_df2rr_ctrl_brType; // @[playground/src/noop/cpu.scala 134:25]
  assign readregs_io_df2rr_rs1 = forwading_io_df2rr_rs1; // @[playground/src/noop/cpu.scala 134:25]
  assign readregs_io_df2rr_rrs1 = forwading_io_df2rr_rrs1; // @[playground/src/noop/cpu.scala 134:25]
  assign readregs_io_df2rr_rs1_d = forwading_io_df2rr_rs1_d; // @[playground/src/noop/cpu.scala 134:25]
  assign readregs_io_df2rr_rs2 = forwading_io_df2rr_rs2; // @[playground/src/noop/cpu.scala 134:25]
  assign readregs_io_df2rr_rrs2 = forwading_io_df2rr_rrs2; // @[playground/src/noop/cpu.scala 134:25]
  assign readregs_io_df2rr_rs2_d = forwading_io_df2rr_rs2_d; // @[playground/src/noop/cpu.scala 134:25]
  assign readregs_io_df2rr_dst = forwading_io_df2rr_dst; // @[playground/src/noop/cpu.scala 134:25]
  assign readregs_io_df2rr_dst_d = forwading_io_df2rr_dst_d; // @[playground/src/noop/cpu.scala 134:25]
  assign readregs_io_df2rr_jmp_type = forwading_io_df2rr_jmp_type; // @[playground/src/noop/cpu.scala 134:25]
  assign readregs_io_df2rr_special = forwading_io_df2rr_special; // @[playground/src/noop/cpu.scala 134:25]
  assign readregs_io_df2rr_swap = forwading_io_df2rr_swap; // @[playground/src/noop/cpu.scala 134:25]
  assign readregs_io_df2rr_indi = forwading_io_df2rr_indi; // @[playground/src/noop/cpu.scala 134:25]
  assign readregs_io_df2rr_recov = forwading_io_df2rr_recov; // @[playground/src/noop/cpu.scala 134:25]
  assign readregs_io_df2rr_valid = forwading_io_df2rr_valid; // @[playground/src/noop/cpu.scala 134:25]
  assign readregs_io_rr2ex_drop = execute_io_rr2ex_drop; // @[playground/src/noop/cpu.scala 140:25]
  assign readregs_io_rr2ex_stall = execute_io_rr2ex_stall; // @[playground/src/noop/cpu.scala 140:25]
  assign readregs_io_rr2ex_ready = execute_io_rr2ex_ready; // @[playground/src/noop/cpu.scala 140:25]
  assign readregs_io_rs1Read_data = regs_io_rs1_data; // @[playground/src/noop/cpu.scala 141:25]
  assign readregs_io_rs2Read_data = regs_io_rs2_data; // @[playground/src/noop/cpu.scala 142:25]
  assign readregs_io_csrRead_data = csrs_io_rs_data; // @[playground/src/noop/cpu.scala 143:25]
  assign readregs_io_csrRead_is_err = csrs_io_rs_is_err; // @[playground/src/noop/cpu.scala 143:25]
  assign execute_clock = clock;
  assign execute_reset = reset;
  assign execute_io_rr2ex_inst = readregs_io_rr2ex_inst; // @[playground/src/noop/cpu.scala 140:25]
  assign execute_io_rr2ex_pc = readregs_io_rr2ex_pc; // @[playground/src/noop/cpu.scala 140:25]
  assign execute_io_rr2ex_excep_cause = readregs_io_rr2ex_excep_cause; // @[playground/src/noop/cpu.scala 140:25]
  assign execute_io_rr2ex_excep_tval = readregs_io_rr2ex_excep_tval; // @[playground/src/noop/cpu.scala 140:25]
  assign execute_io_rr2ex_excep_en = readregs_io_rr2ex_excep_en; // @[playground/src/noop/cpu.scala 140:25]
  assign execute_io_rr2ex_excep_pc = readregs_io_rr2ex_excep_pc; // @[playground/src/noop/cpu.scala 140:25]
  assign execute_io_rr2ex_excep_etype = readregs_io_rr2ex_excep_etype; // @[playground/src/noop/cpu.scala 140:25]
  assign execute_io_rr2ex_ctrl_aluOp = readregs_io_rr2ex_ctrl_aluOp; // @[playground/src/noop/cpu.scala 140:25]
  assign execute_io_rr2ex_ctrl_aluWidth = readregs_io_rr2ex_ctrl_aluWidth; // @[playground/src/noop/cpu.scala 140:25]
  assign execute_io_rr2ex_ctrl_dcMode = readregs_io_rr2ex_ctrl_dcMode; // @[playground/src/noop/cpu.scala 140:25]
  assign execute_io_rr2ex_ctrl_writeRegEn = readregs_io_rr2ex_ctrl_writeRegEn; // @[playground/src/noop/cpu.scala 140:25]
  assign execute_io_rr2ex_ctrl_writeCSREn = readregs_io_rr2ex_ctrl_writeCSREn; // @[playground/src/noop/cpu.scala 140:25]
  assign execute_io_rr2ex_ctrl_brType = readregs_io_rr2ex_ctrl_brType; // @[playground/src/noop/cpu.scala 140:25]
  assign execute_io_rr2ex_rs1_d = readregs_io_rr2ex_rs1_d; // @[playground/src/noop/cpu.scala 140:25]
  assign execute_io_rr2ex_rs2 = readregs_io_rr2ex_rs2; // @[playground/src/noop/cpu.scala 140:25]
  assign execute_io_rr2ex_rs2_d = readregs_io_rr2ex_rs2_d; // @[playground/src/noop/cpu.scala 140:25]
  assign execute_io_rr2ex_dst = readregs_io_rr2ex_dst; // @[playground/src/noop/cpu.scala 140:25]
  assign execute_io_rr2ex_dst_d = readregs_io_rr2ex_dst_d; // @[playground/src/noop/cpu.scala 140:25]
  assign execute_io_rr2ex_rcsr_id = readregs_io_rr2ex_rcsr_id; // @[playground/src/noop/cpu.scala 140:25]
  assign execute_io_rr2ex_jmp_type = readregs_io_rr2ex_jmp_type; // @[playground/src/noop/cpu.scala 140:25]
  assign execute_io_rr2ex_special = readregs_io_rr2ex_special; // @[playground/src/noop/cpu.scala 140:25]
  assign execute_io_rr2ex_indi = readregs_io_rr2ex_indi; // @[playground/src/noop/cpu.scala 140:25]
  assign execute_io_rr2ex_recov = readregs_io_rr2ex_recov; // @[playground/src/noop/cpu.scala 140:25]
  assign execute_io_rr2ex_valid = readregs_io_rr2ex_valid; // @[playground/src/noop/cpu.scala 140:25]
  assign execute_io_ex2mem_drop = memory_io_ex2mem_drop; // @[playground/src/noop/cpu.scala 145:25]
  assign execute_io_ex2mem_stall = memory_io_ex2mem_stall; // @[playground/src/noop/cpu.scala 145:25]
  assign execute_io_ex2mem_ready = memory_io_ex2mem_ready; // @[playground/src/noop/cpu.scala 145:25]
  assign execute_io_updateNextPc_seq_pc = csrs_io_updateNextPc_seq_pc; // @[playground/src/noop/cpu.scala 146:29]
  assign execute_io_updateNextPc_valid = csrs_io_updateNextPc_valid; // @[playground/src/noop/cpu.scala 146:29]
  assign memory_clock = clock;
  assign memory_reset = reset;
  assign memory_io_ex2mem_inst = execute_io_ex2mem_inst; // @[playground/src/noop/cpu.scala 145:25]
  assign memory_io_ex2mem_pc = execute_io_ex2mem_pc; // @[playground/src/noop/cpu.scala 145:25]
  assign memory_io_ex2mem_excep_cause = execute_io_ex2mem_excep_cause; // @[playground/src/noop/cpu.scala 145:25]
  assign memory_io_ex2mem_excep_tval = execute_io_ex2mem_excep_tval; // @[playground/src/noop/cpu.scala 145:25]
  assign memory_io_ex2mem_excep_en = execute_io_ex2mem_excep_en; // @[playground/src/noop/cpu.scala 145:25]
  assign memory_io_ex2mem_excep_pc = execute_io_ex2mem_excep_pc; // @[playground/src/noop/cpu.scala 145:25]
  assign memory_io_ex2mem_excep_etype = execute_io_ex2mem_excep_etype; // @[playground/src/noop/cpu.scala 145:25]
  assign memory_io_ex2mem_ctrl_dcMode = execute_io_ex2mem_ctrl_dcMode; // @[playground/src/noop/cpu.scala 145:25]
  assign memory_io_ex2mem_ctrl_writeRegEn = execute_io_ex2mem_ctrl_writeRegEn; // @[playground/src/noop/cpu.scala 145:25]
  assign memory_io_ex2mem_ctrl_writeCSREn = execute_io_ex2mem_ctrl_writeCSREn; // @[playground/src/noop/cpu.scala 145:25]
  assign memory_io_ex2mem_mem_addr = execute_io_ex2mem_mem_addr; // @[playground/src/noop/cpu.scala 145:25]
  assign memory_io_ex2mem_mem_data = execute_io_ex2mem_mem_data; // @[playground/src/noop/cpu.scala 145:25]
  assign memory_io_ex2mem_csr_id = execute_io_ex2mem_csr_id; // @[playground/src/noop/cpu.scala 145:25]
  assign memory_io_ex2mem_csr_d = execute_io_ex2mem_csr_d; // @[playground/src/noop/cpu.scala 145:25]
  assign memory_io_ex2mem_dst = execute_io_ex2mem_dst; // @[playground/src/noop/cpu.scala 145:25]
  assign memory_io_ex2mem_dst_d = execute_io_ex2mem_dst_d; // @[playground/src/noop/cpu.scala 145:25]
  assign memory_io_ex2mem_rcsr_id = execute_io_ex2mem_rcsr_id; // @[playground/src/noop/cpu.scala 145:25]
  assign memory_io_ex2mem_special = execute_io_ex2mem_special; // @[playground/src/noop/cpu.scala 145:25]
  assign memory_io_ex2mem_indi = execute_io_ex2mem_indi; // @[playground/src/noop/cpu.scala 145:25]
  assign memory_io_ex2mem_recov = execute_io_ex2mem_recov; // @[playground/src/noop/cpu.scala 145:25]
  assign memory_io_ex2mem_valid = execute_io_ex2mem_valid; // @[playground/src/noop/cpu.scala 145:25]
  assign memory_io_mem2rb_drop = writeback_io_mem2rb_drop; // @[playground/src/noop/cpu.scala 147:25]
  assign memory_io_mem2rb_stall = writeback_io_mem2rb_stall; // @[playground/src/noop/cpu.scala 147:25]
  assign memory_io_mem2rb_ready = writeback_io_mem2rb_ready; // @[playground/src/noop/cpu.scala 147:25]
  assign memory_io_dataRW_rdata = memCrossbar_io_dataRW_rdata; // @[playground/src/noop/cpu.scala 148:25]
  assign memory_io_dataRW_rvalid = memCrossbar_io_dataRW_rvalid; // @[playground/src/noop/cpu.scala 148:25]
  assign memory_io_dataRW_ready = memCrossbar_io_dataRW_ready; // @[playground/src/noop/cpu.scala 148:25]
  assign memory_io_va2pa_paddr = tlb_mem_io_va2pa_paddr; // @[playground/src/noop/cpu.scala 149:25]
  assign memory_io_va2pa_pvalid = tlb_mem_io_va2pa_pvalid; // @[playground/src/noop/cpu.scala 149:25]
  assign memory_io_va2pa_tlb_excep_cause = tlb_mem_io_va2pa_tlb_excep_cause; // @[playground/src/noop/cpu.scala 149:25]
  assign memory_io_va2pa_tlb_excep_tval = tlb_mem_io_va2pa_tlb_excep_tval; // @[playground/src/noop/cpu.scala 149:25]
  assign memory_io_va2pa_tlb_excep_en = tlb_mem_io_va2pa_tlb_excep_en; // @[playground/src/noop/cpu.scala 149:25]
  assign writeback_clock = clock;
  assign writeback_reset = reset;
  assign writeback_io_mem2rb_inst = memory_io_mem2rb_inst; // @[playground/src/noop/cpu.scala 147:25]
  assign writeback_io_mem2rb_pc = memory_io_mem2rb_pc; // @[playground/src/noop/cpu.scala 147:25]
  assign writeback_io_mem2rb_excep_cause = memory_io_mem2rb_excep_cause; // @[playground/src/noop/cpu.scala 147:25]
  assign writeback_io_mem2rb_excep_tval = memory_io_mem2rb_excep_tval; // @[playground/src/noop/cpu.scala 147:25]
  assign writeback_io_mem2rb_excep_en = memory_io_mem2rb_excep_en; // @[playground/src/noop/cpu.scala 147:25]
  assign writeback_io_mem2rb_excep_pc = memory_io_mem2rb_excep_pc; // @[playground/src/noop/cpu.scala 147:25]
  assign writeback_io_mem2rb_excep_etype = memory_io_mem2rb_excep_etype; // @[playground/src/noop/cpu.scala 147:25]
  assign writeback_io_mem2rb_csr_id = memory_io_mem2rb_csr_id; // @[playground/src/noop/cpu.scala 147:25]
  assign writeback_io_mem2rb_csr_d = memory_io_mem2rb_csr_d; // @[playground/src/noop/cpu.scala 147:25]
  assign writeback_io_mem2rb_csr_en = memory_io_mem2rb_csr_en; // @[playground/src/noop/cpu.scala 147:25]
  assign writeback_io_mem2rb_dst = memory_io_mem2rb_dst; // @[playground/src/noop/cpu.scala 147:25]
  assign writeback_io_mem2rb_dst_d = memory_io_mem2rb_dst_d; // @[playground/src/noop/cpu.scala 147:25]
  assign writeback_io_mem2rb_dst_en = memory_io_mem2rb_dst_en; // @[playground/src/noop/cpu.scala 147:25]
  assign writeback_io_mem2rb_rcsr_id = memory_io_mem2rb_rcsr_id; // @[playground/src/noop/cpu.scala 147:25]
  assign writeback_io_mem2rb_special = memory_io_mem2rb_special; // @[playground/src/noop/cpu.scala 147:25]
  assign writeback_io_mem2rb_is_mmio = memory_io_mem2rb_is_mmio; // @[playground/src/noop/cpu.scala 147:25]
  assign writeback_io_mem2rb_recov = memory_io_mem2rb_recov; // @[playground/src/noop/cpu.scala 147:25]
  assign writeback_io_mem2rb_valid = memory_io_mem2rb_valid; // @[playground/src/noop/cpu.scala 147:25]
  assign regs_clock = clock;
  assign regs_reset = reset;
  assign regs_io_rs1_id = readregs_io_rs1Read_id; // @[playground/src/noop/cpu.scala 141:25]
  assign regs_io_rs2_id = readregs_io_rs2Read_id; // @[playground/src/noop/cpu.scala 142:25]
  assign regs_io_dst_id = writeback_io_wReg_id; // @[playground/src/noop/cpu.scala 151:25]
  assign regs_io_dst_data = writeback_io_wReg_data; // @[playground/src/noop/cpu.scala 151:25]
  assign regs_io_dst_en = writeback_io_wReg_en; // @[playground/src/noop/cpu.scala 151:25]
  assign csrs_clock = clock;
  assign csrs_reset = reset;
  assign csrs_io_rs_id = readregs_io_csrRead_id; // @[playground/src/noop/cpu.scala 143:25]
  assign csrs_io_rd_id = writeback_io_wCsr_id; // @[playground/src/noop/cpu.scala 152:25]
  assign csrs_io_rd_data = writeback_io_wCsr_data; // @[playground/src/noop/cpu.scala 152:25]
  assign csrs_io_rd_en = writeback_io_wCsr_en; // @[playground/src/noop/cpu.scala 152:25]
  assign csrs_io_excep_cause = writeback_io_excep_cause; // @[playground/src/noop/cpu.scala 153:25]
  assign csrs_io_excep_tval = writeback_io_excep_tval; // @[playground/src/noop/cpu.scala 153:25]
  assign csrs_io_excep_en = writeback_io_excep_en; // @[playground/src/noop/cpu.scala 153:25]
  assign csrs_io_excep_pc = writeback_io_excep_pc; // @[playground/src/noop/cpu.scala 153:25]
  assign csrs_io_excep_etype = writeback_io_excep_etype; // @[playground/src/noop/cpu.scala 153:25]
  assign csrs_io_clint_raise = clint_io_intr_raise; // @[playground/src/noop/cpu.scala 154:25]
  assign csrs_io_clint_clear = clint_io_intr_clear; // @[playground/src/noop/cpu.scala 154:25]
  assign csrs_io_plic_m_raise = plic_io_intr_out_m_raise; // @[playground/src/noop/cpu.scala 181:25]
  assign csrs_io_plic_m_clear = plic_io_intr_out_m_clear; // @[playground/src/noop/cpu.scala 181:25]
  assign csrs_io_plic_s_raise = plic_io_intr_out_s_raise; // @[playground/src/noop/cpu.scala 182:25]
  assign csrs_io_plic_s_clear = plic_io_intr_out_s_clear; // @[playground/src/noop/cpu.scala 182:25]
  assign csrs_io_intr_msip_raise = clint_io_intr_msip_raise; // @[playground/src/noop/cpu.scala 155:25]
  assign csrs_io_intr_msip_clear = clint_io_intr_msip_clear; // @[playground/src/noop/cpu.scala 155:25]
  assign icache_clock = clock;
  assign icache_reset = reset;
  assign icache_io_instAxi_ra_ready = crossBar_io_icAxi_ra_ready; // @[playground/src/noop/cpu.scala 174:25]
  assign icache_io_instAxi_rd_valid = crossBar_io_icAxi_rd_valid; // @[playground/src/noop/cpu.scala 174:25]
  assign icache_io_instAxi_rd_bits_data = crossBar_io_icAxi_rd_bits_data; // @[playground/src/noop/cpu.scala 174:25]
  assign icache_io_instAxi_rd_bits_last = crossBar_io_icAxi_rd_bits_last; // @[playground/src/noop/cpu.scala 174:25]
  assign icache_io_icRead_addr = fetchCrossbar_io_icRead_addr; // @[playground/src/noop/cpu.scala 162:33]
  assign icache_io_icRead_arvalid = fetchCrossbar_io_icRead_arvalid; // @[playground/src/noop/cpu.scala 162:33]
  assign icache_io_flush = writeback_io_flush_cache; // @[playground/src/noop/cpu.scala 157:25]
  assign dcache_clock = clock;
  assign dcache_reset = reset;
  assign dcache_io_dataAxi_wa_ready = crossBar_io_memAxi_wa_ready; // @[playground/src/noop/cpu.scala 175:25]
  assign dcache_io_dataAxi_wd_ready = crossBar_io_memAxi_wd_ready; // @[playground/src/noop/cpu.scala 175:25]
  assign dcache_io_dataAxi_ra_ready = crossBar_io_memAxi_ra_ready; // @[playground/src/noop/cpu.scala 175:25]
  assign dcache_io_dataAxi_rd_valid = crossBar_io_memAxi_rd_valid; // @[playground/src/noop/cpu.scala 175:25]
  assign dcache_io_dataAxi_rd_bits_data = crossBar_io_memAxi_rd_bits_data; // @[playground/src/noop/cpu.scala 175:25]
  assign dcache_io_dataAxi_rd_bits_last = crossBar_io_memAxi_rd_bits_last; // @[playground/src/noop/cpu.scala 175:25]
  assign dcache_io_dcRW_addr = dcSelector_io_select_addr; // @[playground/src/noop/cpu.scala 168:33]
  assign dcache_io_dcRW_wdata = dcSelector_io_select_wdata; // @[playground/src/noop/cpu.scala 168:33]
  assign dcache_io_dcRW_dc_mode = dcSelector_io_select_dc_mode; // @[playground/src/noop/cpu.scala 168:33]
  assign dcache_io_dcRW_amo = dcSelector_io_select_amo; // @[playground/src/noop/cpu.scala 168:33]
  assign dcache_io_flush = writeback_io_flush_cache; // @[playground/src/noop/cpu.scala 158:25]
  assign mem2Axi_clock = clock;
  assign mem2Axi_reset = reset;
  assign mem2Axi_io_dataIO_addr = memCrossbar_io_mmio_addr; // @[playground/src/noop/cpu.scala 166:33]
  assign mem2Axi_io_dataIO_wdata = memCrossbar_io_mmio_wdata; // @[playground/src/noop/cpu.scala 166:33]
  assign mem2Axi_io_dataIO_dc_mode = memCrossbar_io_mmio_dc_mode; // @[playground/src/noop/cpu.scala 166:33]
  assign mem2Axi_io_outAxi_wa_ready = crossBar_io_mmioAxi_wa_ready; // @[playground/src/noop/cpu.scala 176:25]
  assign mem2Axi_io_outAxi_wd_ready = crossBar_io_mmioAxi_wd_ready; // @[playground/src/noop/cpu.scala 176:25]
  assign mem2Axi_io_outAxi_wr_valid = crossBar_io_mmioAxi_wr_valid; // @[playground/src/noop/cpu.scala 176:25]
  assign mem2Axi_io_outAxi_wr_bits_id = crossBar_io_mmioAxi_wr_bits_id; // @[playground/src/noop/cpu.scala 176:25]
  assign mem2Axi_io_outAxi_wr_bits_resp = crossBar_io_mmioAxi_wr_bits_resp; // @[playground/src/noop/cpu.scala 176:25]
  assign mem2Axi_io_outAxi_ra_ready = crossBar_io_mmioAxi_ra_ready; // @[playground/src/noop/cpu.scala 176:25]
  assign mem2Axi_io_outAxi_rd_valid = crossBar_io_mmioAxi_rd_valid; // @[playground/src/noop/cpu.scala 176:25]
  assign mem2Axi_io_outAxi_rd_bits_id = crossBar_io_mmioAxi_rd_bits_id; // @[playground/src/noop/cpu.scala 176:25]
  assign mem2Axi_io_outAxi_rd_bits_data = crossBar_io_mmioAxi_rd_bits_data; // @[playground/src/noop/cpu.scala 176:25]
  assign mem2Axi_io_outAxi_rd_bits_resp = crossBar_io_mmioAxi_rd_bits_resp; // @[playground/src/noop/cpu.scala 176:25]
  assign mem2Axi_io_outAxi_rd_bits_last = crossBar_io_mmioAxi_rd_bits_last; // @[playground/src/noop/cpu.scala 176:25]
  assign flash2Axi_clock = clock;
  assign flash2Axi_reset = reset;
  assign flash2Axi_io_dataIO_addr = split64to32_io_data_out_addr; // @[playground/src/noop/cpu.scala 164:33]
  assign flash2Axi_io_dataIO_wdata = 64'h0; // @[playground/src/noop/cpu.scala 164:33]
  assign flash2Axi_io_dataIO_dc_mode = split64to32_io_data_out_dc_mode; // @[playground/src/noop/cpu.scala 164:33]
  assign flash2Axi_io_outAxi_wa_ready = crossBar_io_flashAxi_wa_ready; // @[playground/src/noop/cpu.scala 177:26]
  assign flash2Axi_io_outAxi_wd_ready = crossBar_io_flashAxi_wd_ready; // @[playground/src/noop/cpu.scala 177:26]
  assign flash2Axi_io_outAxi_wr_valid = crossBar_io_flashAxi_wr_valid; // @[playground/src/noop/cpu.scala 177:26]
  assign flash2Axi_io_outAxi_wr_bits_id = crossBar_io_flashAxi_wr_bits_id; // @[playground/src/noop/cpu.scala 177:26]
  assign flash2Axi_io_outAxi_wr_bits_resp = crossBar_io_flashAxi_wr_bits_resp; // @[playground/src/noop/cpu.scala 177:26]
  assign flash2Axi_io_outAxi_ra_ready = crossBar_io_flashAxi_ra_ready; // @[playground/src/noop/cpu.scala 177:26]
  assign flash2Axi_io_outAxi_rd_valid = crossBar_io_flashAxi_rd_valid; // @[playground/src/noop/cpu.scala 177:26]
  assign flash2Axi_io_outAxi_rd_bits_id = crossBar_io_flashAxi_rd_bits_id; // @[playground/src/noop/cpu.scala 177:26]
  assign flash2Axi_io_outAxi_rd_bits_data = crossBar_io_flashAxi_rd_bits_data; // @[playground/src/noop/cpu.scala 177:26]
  assign flash2Axi_io_outAxi_rd_bits_resp = crossBar_io_flashAxi_rd_bits_resp; // @[playground/src/noop/cpu.scala 177:26]
  assign flash2Axi_io_outAxi_rd_bits_last = crossBar_io_flashAxi_rd_bits_last; // @[playground/src/noop/cpu.scala 177:26]
  assign crossBar_clock = clock;
  assign crossBar_reset = reset;
  assign crossBar_io_icAxi_ra_valid = icache_io_instAxi_ra_valid; // @[playground/src/noop/cpu.scala 174:25]
  assign crossBar_io_icAxi_ra_bits_addr = icache_io_instAxi_ra_bits_addr; // @[playground/src/noop/cpu.scala 174:25]
  assign crossBar_io_flashAxi_wa_valid = flash2Axi_io_outAxi_wa_valid; // @[playground/src/noop/cpu.scala 177:26]
  assign crossBar_io_flashAxi_wa_bits_id = flash2Axi_io_outAxi_wa_bits_id; // @[playground/src/noop/cpu.scala 177:26]
  assign crossBar_io_flashAxi_wa_bits_addr = flash2Axi_io_outAxi_wa_bits_addr; // @[playground/src/noop/cpu.scala 177:26]
  assign crossBar_io_flashAxi_wa_bits_len = flash2Axi_io_outAxi_wa_bits_len; // @[playground/src/noop/cpu.scala 177:26]
  assign crossBar_io_flashAxi_wa_bits_size = flash2Axi_io_outAxi_wa_bits_size; // @[playground/src/noop/cpu.scala 177:26]
  assign crossBar_io_flashAxi_wa_bits_burst = flash2Axi_io_outAxi_wa_bits_burst; // @[playground/src/noop/cpu.scala 177:26]
  assign crossBar_io_flashAxi_wd_valid = flash2Axi_io_outAxi_wd_valid; // @[playground/src/noop/cpu.scala 177:26]
  assign crossBar_io_flashAxi_wd_bits_data = flash2Axi_io_outAxi_wd_bits_data; // @[playground/src/noop/cpu.scala 177:26]
  assign crossBar_io_flashAxi_wd_bits_strb = flash2Axi_io_outAxi_wd_bits_strb; // @[playground/src/noop/cpu.scala 177:26]
  assign crossBar_io_flashAxi_wd_bits_last = flash2Axi_io_outAxi_wd_bits_last; // @[playground/src/noop/cpu.scala 177:26]
  assign crossBar_io_flashAxi_wr_ready = flash2Axi_io_outAxi_wr_ready; // @[playground/src/noop/cpu.scala 177:26]
  assign crossBar_io_flashAxi_ra_valid = flash2Axi_io_outAxi_ra_valid; // @[playground/src/noop/cpu.scala 177:26]
  assign crossBar_io_flashAxi_ra_bits_id = flash2Axi_io_outAxi_ra_bits_id; // @[playground/src/noop/cpu.scala 177:26]
  assign crossBar_io_flashAxi_ra_bits_addr = flash2Axi_io_outAxi_ra_bits_addr; // @[playground/src/noop/cpu.scala 177:26]
  assign crossBar_io_flashAxi_ra_bits_len = flash2Axi_io_outAxi_ra_bits_len; // @[playground/src/noop/cpu.scala 177:26]
  assign crossBar_io_flashAxi_ra_bits_size = flash2Axi_io_outAxi_ra_bits_size; // @[playground/src/noop/cpu.scala 177:26]
  assign crossBar_io_flashAxi_ra_bits_burst = flash2Axi_io_outAxi_ra_bits_burst; // @[playground/src/noop/cpu.scala 177:26]
  assign crossBar_io_flashAxi_rd_ready = flash2Axi_io_outAxi_rd_ready; // @[playground/src/noop/cpu.scala 177:26]
  assign crossBar_io_memAxi_wa_valid = dcache_io_dataAxi_wa_valid; // @[playground/src/noop/cpu.scala 175:25]
  assign crossBar_io_memAxi_wa_bits_addr = dcache_io_dataAxi_wa_bits_addr; // @[playground/src/noop/cpu.scala 175:25]
  assign crossBar_io_memAxi_wd_valid = dcache_io_dataAxi_wd_valid; // @[playground/src/noop/cpu.scala 175:25]
  assign crossBar_io_memAxi_wd_bits_data = dcache_io_dataAxi_wd_bits_data; // @[playground/src/noop/cpu.scala 175:25]
  assign crossBar_io_memAxi_wd_bits_last = dcache_io_dataAxi_wd_bits_last; // @[playground/src/noop/cpu.scala 175:25]
  assign crossBar_io_memAxi_ra_valid = dcache_io_dataAxi_ra_valid; // @[playground/src/noop/cpu.scala 175:25]
  assign crossBar_io_memAxi_ra_bits_addr = dcache_io_dataAxi_ra_bits_addr; // @[playground/src/noop/cpu.scala 175:25]
  assign crossBar_io_mmioAxi_wa_valid = mem2Axi_io_outAxi_wa_valid; // @[playground/src/noop/cpu.scala 176:25]
  assign crossBar_io_mmioAxi_wa_bits_id = mem2Axi_io_outAxi_wa_bits_id; // @[playground/src/noop/cpu.scala 176:25]
  assign crossBar_io_mmioAxi_wa_bits_addr = mem2Axi_io_outAxi_wa_bits_addr; // @[playground/src/noop/cpu.scala 176:25]
  assign crossBar_io_mmioAxi_wa_bits_len = mem2Axi_io_outAxi_wa_bits_len; // @[playground/src/noop/cpu.scala 176:25]
  assign crossBar_io_mmioAxi_wa_bits_size = mem2Axi_io_outAxi_wa_bits_size; // @[playground/src/noop/cpu.scala 176:25]
  assign crossBar_io_mmioAxi_wa_bits_burst = mem2Axi_io_outAxi_wa_bits_burst; // @[playground/src/noop/cpu.scala 176:25]
  assign crossBar_io_mmioAxi_wd_valid = mem2Axi_io_outAxi_wd_valid; // @[playground/src/noop/cpu.scala 176:25]
  assign crossBar_io_mmioAxi_wd_bits_data = mem2Axi_io_outAxi_wd_bits_data; // @[playground/src/noop/cpu.scala 176:25]
  assign crossBar_io_mmioAxi_wd_bits_strb = mem2Axi_io_outAxi_wd_bits_strb; // @[playground/src/noop/cpu.scala 176:25]
  assign crossBar_io_mmioAxi_wd_bits_last = mem2Axi_io_outAxi_wd_bits_last; // @[playground/src/noop/cpu.scala 176:25]
  assign crossBar_io_mmioAxi_wr_ready = mem2Axi_io_outAxi_wr_ready; // @[playground/src/noop/cpu.scala 176:25]
  assign crossBar_io_mmioAxi_ra_valid = mem2Axi_io_outAxi_ra_valid; // @[playground/src/noop/cpu.scala 176:25]
  assign crossBar_io_mmioAxi_ra_bits_id = mem2Axi_io_outAxi_ra_bits_id; // @[playground/src/noop/cpu.scala 176:25]
  assign crossBar_io_mmioAxi_ra_bits_addr = mem2Axi_io_outAxi_ra_bits_addr; // @[playground/src/noop/cpu.scala 176:25]
  assign crossBar_io_mmioAxi_ra_bits_len = mem2Axi_io_outAxi_ra_bits_len; // @[playground/src/noop/cpu.scala 176:25]
  assign crossBar_io_mmioAxi_ra_bits_size = mem2Axi_io_outAxi_ra_bits_size; // @[playground/src/noop/cpu.scala 176:25]
  assign crossBar_io_mmioAxi_ra_bits_burst = mem2Axi_io_outAxi_ra_bits_burst; // @[playground/src/noop/cpu.scala 176:25]
  assign crossBar_io_mmioAxi_rd_ready = mem2Axi_io_outAxi_rd_ready; // @[playground/src/noop/cpu.scala 176:25]
  assign crossBar_io_outAxi_wa_ready = io_master_awready; // @[playground/src/noop/cpu.scala 188:36]
  assign crossBar_io_outAxi_wd_ready = io_master_wready; // @[playground/src/noop/cpu.scala 196:35]
  assign crossBar_io_outAxi_wr_valid = io_master_bvalid; // @[playground/src/noop/cpu.scala 203:40]
  assign crossBar_io_outAxi_wr_bits_id = io_master_bid; // @[playground/src/noop/cpu.scala 205:40]
  assign crossBar_io_outAxi_wr_bits_resp = io_master_bresp; // @[playground/src/noop/cpu.scala 204:40]
  assign crossBar_io_outAxi_ra_ready = io_master_arready; // @[playground/src/noop/cpu.scala 207:34]
  assign crossBar_io_outAxi_rd_valid = io_master_rvalid; // @[playground/src/noop/cpu.scala 216:35]
  assign crossBar_io_outAxi_rd_bits_id = io_master_rid; // @[playground/src/noop/cpu.scala 220:40]
  assign crossBar_io_outAxi_rd_bits_data = io_master_rdata; // @[playground/src/noop/cpu.scala 218:40]
  assign crossBar_io_outAxi_rd_bits_resp = io_master_rresp; // @[playground/src/noop/cpu.scala 217:40]
  assign crossBar_io_outAxi_rd_bits_last = io_master_rlast; // @[playground/src/noop/cpu.scala 219:40]
  assign crossBar_io_selectMem = dcache_io_flush_out; // @[playground/src/noop/cpu.scala 178:27]
  assign fetchCrossbar_clock = clock;
  assign fetchCrossbar_reset = reset;
  assign fetchCrossbar_io_instIO_addr = fetch_io_instRead_addr; // @[playground/src/noop/cpu.scala 123:25]
  assign fetchCrossbar_io_instIO_arvalid = fetch_io_instRead_arvalid; // @[playground/src/noop/cpu.scala 123:25]
  assign fetchCrossbar_io_icRead_inst = icache_io_icRead_inst; // @[playground/src/noop/cpu.scala 162:33]
  assign fetchCrossbar_io_icRead_rvalid = icache_io_icRead_rvalid; // @[playground/src/noop/cpu.scala 162:33]
  assign fetchCrossbar_io_flashRead_rdata = split64to32_io_data_in_rdata; // @[playground/src/noop/cpu.scala 163:33]
  assign fetchCrossbar_io_flashRead_rvalid = split64to32_io_data_in_rvalid; // @[playground/src/noop/cpu.scala 163:33]
  assign split64to32_clock = clock;
  assign split64to32_reset = reset;
  assign split64to32_io_data_in_addr = fetchCrossbar_io_flashRead_addr; // @[playground/src/noop/cpu.scala 163:33]
  assign split64to32_io_data_in_dc_mode = fetchCrossbar_io_flashRead_dc_mode; // @[playground/src/noop/cpu.scala 163:33]
  assign split64to32_io_data_out_rdata = flash2Axi_io_dataIO_rdata; // @[playground/src/noop/cpu.scala 164:33]
  assign split64to32_io_data_out_rvalid = flash2Axi_io_dataIO_rvalid; // @[playground/src/noop/cpu.scala 164:33]
  assign split64to32_io_data_out_ready = flash2Axi_io_dataIO_ready; // @[playground/src/noop/cpu.scala 164:33]
  assign memCrossbar_clock = clock;
  assign memCrossbar_reset = reset;
  assign memCrossbar_io_dataRW_addr = memory_io_dataRW_addr; // @[playground/src/noop/cpu.scala 148:25]
  assign memCrossbar_io_dataRW_wdata = memory_io_dataRW_wdata; // @[playground/src/noop/cpu.scala 148:25]
  assign memCrossbar_io_dataRW_dc_mode = memory_io_dataRW_dc_mode; // @[playground/src/noop/cpu.scala 148:25]
  assign memCrossbar_io_dataRW_amo = memory_io_dataRW_amo; // @[playground/src/noop/cpu.scala 148:25]
  assign memCrossbar_io_mmio_rdata = mem2Axi_io_dataIO_rdata; // @[playground/src/noop/cpu.scala 166:33]
  assign memCrossbar_io_mmio_rvalid = mem2Axi_io_dataIO_rvalid; // @[playground/src/noop/cpu.scala 166:33]
  assign memCrossbar_io_mmio_ready = mem2Axi_io_dataIO_ready; // @[playground/src/noop/cpu.scala 166:33]
  assign memCrossbar_io_dcRW_rdata = dcSelector_io_mem2dc_rdata; // @[playground/src/noop/cpu.scala 165:33]
  assign memCrossbar_io_dcRW_rvalid = dcSelector_io_mem2dc_rvalid; // @[playground/src/noop/cpu.scala 165:33]
  assign memCrossbar_io_dcRW_ready = dcSelector_io_mem2dc_ready; // @[playground/src/noop/cpu.scala 165:33]
  assign memCrossbar_io_clintIO_rdata = clint_io_rw_rdata; // @[playground/src/noop/cpu.scala 167:33]
  assign memCrossbar_io_plicIO_rdata = plic_io_rw_rdata; // @[playground/src/noop/cpu.scala 183:25]
  assign tlb_if_clock = clock;
  assign tlb_if_reset = reset;
  assign tlb_if_io_va2pa_vaddr = fetch_io_va2pa_vaddr; // @[playground/src/noop/cpu.scala 124:25]
  assign tlb_if_io_va2pa_vvalid = fetch_io_va2pa_vvalid; // @[playground/src/noop/cpu.scala 124:25]
  assign tlb_if_io_mmuState_priv = csrs_io_mmuState_priv; // @[playground/src/noop/cpu.scala 170:33]
  assign tlb_if_io_mmuState_mstatus = csrs_io_mmuState_mstatus; // @[playground/src/noop/cpu.scala 170:33]
  assign tlb_if_io_mmuState_satp = csrs_io_mmuState_satp; // @[playground/src/noop/cpu.scala 170:33]
  assign tlb_if_io_flush = writeback_io_flush_tlb; // @[playground/src/noop/cpu.scala 159:25]
  assign tlb_if_io_dcacheRW_rdata = dcSelector_io_tlb_if2dc_rdata; // @[playground/src/noop/cpu.scala 169:33]
  assign tlb_if_io_dcacheRW_rvalid = dcSelector_io_tlb_if2dc_rvalid; // @[playground/src/noop/cpu.scala 169:33]
  assign tlb_if_io_dcacheRW_ready = dcSelector_io_tlb_if2dc_ready; // @[playground/src/noop/cpu.scala 169:33]
  assign tlb_mem_clock = clock;
  assign tlb_mem_reset = reset;
  assign tlb_mem_io_va2pa_vaddr = memory_io_va2pa_vaddr; // @[playground/src/noop/cpu.scala 149:25]
  assign tlb_mem_io_va2pa_vvalid = memory_io_va2pa_vvalid; // @[playground/src/noop/cpu.scala 149:25]
  assign tlb_mem_io_va2pa_m_type = memory_io_va2pa_m_type; // @[playground/src/noop/cpu.scala 149:25]
  assign tlb_mem_io_mmuState_priv = csrs_io_mmuState_priv; // @[playground/src/noop/cpu.scala 172:33]
  assign tlb_mem_io_mmuState_mstatus = csrs_io_mmuState_mstatus; // @[playground/src/noop/cpu.scala 172:33]
  assign tlb_mem_io_mmuState_satp = csrs_io_mmuState_satp; // @[playground/src/noop/cpu.scala 172:33]
  assign tlb_mem_io_flush = writeback_io_flush_tlb; // @[playground/src/noop/cpu.scala 160:25]
  assign tlb_mem_io_dcacheRW_rdata = dcSelector_io_tlb_mem2dc_rdata; // @[playground/src/noop/cpu.scala 171:33]
  assign tlb_mem_io_dcacheRW_rvalid = dcSelector_io_tlb_mem2dc_rvalid; // @[playground/src/noop/cpu.scala 171:33]
  assign tlb_mem_io_dcacheRW_ready = dcSelector_io_tlb_mem2dc_ready; // @[playground/src/noop/cpu.scala 171:33]
  assign dcSelector_clock = clock;
  assign dcSelector_reset = reset;
  assign dcSelector_io_tlb_if2dc_addr = tlb_if_io_dcacheRW_addr; // @[playground/src/noop/cpu.scala 169:33]
  assign dcSelector_io_tlb_if2dc_wdata = tlb_if_io_dcacheRW_wdata; // @[playground/src/noop/cpu.scala 169:33]
  assign dcSelector_io_tlb_if2dc_dc_mode = tlb_if_io_dcacheRW_dc_mode; // @[playground/src/noop/cpu.scala 169:33]
  assign dcSelector_io_tlb_mem2dc_addr = tlb_mem_io_dcacheRW_addr; // @[playground/src/noop/cpu.scala 171:33]
  assign dcSelector_io_tlb_mem2dc_wdata = tlb_mem_io_dcacheRW_wdata; // @[playground/src/noop/cpu.scala 171:33]
  assign dcSelector_io_tlb_mem2dc_dc_mode = tlb_mem_io_dcacheRW_dc_mode; // @[playground/src/noop/cpu.scala 171:33]
  assign dcSelector_io_mem2dc_addr = memCrossbar_io_dcRW_addr; // @[playground/src/noop/cpu.scala 165:33]
  assign dcSelector_io_mem2dc_wdata = memCrossbar_io_dcRW_wdata; // @[playground/src/noop/cpu.scala 165:33]
  assign dcSelector_io_mem2dc_dc_mode = memCrossbar_io_dcRW_dc_mode; // @[playground/src/noop/cpu.scala 165:33]
  assign dcSelector_io_mem2dc_amo = memCrossbar_io_dcRW_amo; // @[playground/src/noop/cpu.scala 165:33]
  assign dcSelector_io_dma2dc_addr = dmaBridge_io_dcRW_addr; // @[playground/src/noop/cpu.scala 186:23]
  assign dcSelector_io_dma2dc_wdata = dmaBridge_io_dcRW_wdata; // @[playground/src/noop/cpu.scala 186:23]
  assign dcSelector_io_dma2dc_dc_mode = dmaBridge_io_dcRW_dc_mode; // @[playground/src/noop/cpu.scala 186:23]
  assign dcSelector_io_select_rdata = dcache_io_dcRW_rdata; // @[playground/src/noop/cpu.scala 168:33]
  assign dcSelector_io_select_rvalid = dcache_io_dcRW_rvalid; // @[playground/src/noop/cpu.scala 168:33]
  assign dcSelector_io_select_ready = dcache_io_dcRW_ready; // @[playground/src/noop/cpu.scala 168:33]
  assign clint_clock = clock;
  assign clint_reset = reset;
  assign clint_io_rw_addr = memCrossbar_io_clintIO_addr; // @[playground/src/noop/cpu.scala 167:33]
  assign clint_io_rw_wdata = memCrossbar_io_clintIO_wdata; // @[playground/src/noop/cpu.scala 167:33]
  assign clint_io_rw_wvalid = memCrossbar_io_clintIO_wvalid; // @[playground/src/noop/cpu.scala 167:33]
  assign plic_clock = clock;
  assign plic_reset = reset;
  assign plic_io_intr_in1 = io_interrupt; // @[playground/src/noop/cpu.scala 180:25]
  assign plic_io_rw_addr = memCrossbar_io_plicIO_addr; // @[playground/src/noop/cpu.scala 183:25]
  assign plic_io_rw_wdata = memCrossbar_io_plicIO_wdata; // @[playground/src/noop/cpu.scala 183:25]
  assign plic_io_rw_wvalid = memCrossbar_io_plicIO_wvalid; // @[playground/src/noop/cpu.scala 183:25]
  assign plic_io_rw_arvalid = memCrossbar_io_plicIO_arvalid; // @[playground/src/noop/cpu.scala 183:25]
  assign dmaBridge_clock = clock;
  assign dmaBridge_reset = reset;
  assign dmaBridge_io_dmaAxi_awvalid = io_slave_awvalid; // @[playground/src/noop/cpu.scala 185:14]
  assign dmaBridge_io_dmaAxi_awaddr = io_slave_awaddr; // @[playground/src/noop/cpu.scala 185:14]
  assign dmaBridge_io_dmaAxi_awid = io_slave_awid; // @[playground/src/noop/cpu.scala 185:14]
  assign dmaBridge_io_dmaAxi_awlen = io_slave_awlen; // @[playground/src/noop/cpu.scala 185:14]
  assign dmaBridge_io_dmaAxi_awsize = io_slave_awsize; // @[playground/src/noop/cpu.scala 185:14]
  assign dmaBridge_io_dmaAxi_wvalid = io_slave_wvalid; // @[playground/src/noop/cpu.scala 185:14]
  assign dmaBridge_io_dmaAxi_wdata = io_slave_wdata; // @[playground/src/noop/cpu.scala 185:14]
  assign dmaBridge_io_dmaAxi_wstrb = io_slave_wstrb; // @[playground/src/noop/cpu.scala 185:14]
  assign dmaBridge_io_dmaAxi_bready = io_slave_bready; // @[playground/src/noop/cpu.scala 185:14]
  assign dmaBridge_io_dmaAxi_arvalid = io_slave_arvalid; // @[playground/src/noop/cpu.scala 185:14]
  assign dmaBridge_io_dmaAxi_araddr = io_slave_araddr; // @[playground/src/noop/cpu.scala 185:14]
  assign dmaBridge_io_dmaAxi_arid = io_slave_arid; // @[playground/src/noop/cpu.scala 185:14]
  assign dmaBridge_io_dmaAxi_arlen = io_slave_arlen; // @[playground/src/noop/cpu.scala 185:14]
  assign dmaBridge_io_dmaAxi_arsize = io_slave_arsize; // @[playground/src/noop/cpu.scala 185:14]
  assign dmaBridge_io_dmaAxi_rready = io_slave_rready; // @[playground/src/noop/cpu.scala 185:14]
  assign dmaBridge_io_dcRW_rdata = dcSelector_io_dma2dc_rdata; // @[playground/src/noop/cpu.scala 186:23]
  assign dmaBridge_io_dcRW_rvalid = dcSelector_io_dma2dc_rvalid; // @[playground/src/noop/cpu.scala 186:23]
  assign dmaBridge_io_dcRW_ready = dcSelector_io_dma2dc_ready; // @[playground/src/noop/cpu.scala 186:23]
endmodule
module SimMEM(
  input         clock,
  input         reset,
  output        io_memAxi_wa_ready, // @[playground/src/sim/sim_mem.scala 16:16]
  input         io_memAxi_wa_valid, // @[playground/src/sim/sim_mem.scala 16:16]
  input  [3:0]  io_memAxi_wa_bits_id, // @[playground/src/sim/sim_mem.scala 16:16]
  input  [31:0] io_memAxi_wa_bits_addr, // @[playground/src/sim/sim_mem.scala 16:16]
  input  [7:0]  io_memAxi_wa_bits_len, // @[playground/src/sim/sim_mem.scala 16:16]
  input  [2:0]  io_memAxi_wa_bits_size, // @[playground/src/sim/sim_mem.scala 16:16]
  input  [1:0]  io_memAxi_wa_bits_burst, // @[playground/src/sim/sim_mem.scala 16:16]
  output        io_memAxi_wd_ready, // @[playground/src/sim/sim_mem.scala 16:16]
  input         io_memAxi_wd_valid, // @[playground/src/sim/sim_mem.scala 16:16]
  input  [63:0] io_memAxi_wd_bits_data, // @[playground/src/sim/sim_mem.scala 16:16]
  input  [7:0]  io_memAxi_wd_bits_strb, // @[playground/src/sim/sim_mem.scala 16:16]
  input         io_memAxi_wd_bits_last, // @[playground/src/sim/sim_mem.scala 16:16]
  input         io_memAxi_wr_ready, // @[playground/src/sim/sim_mem.scala 16:16]
  output        io_memAxi_wr_valid, // @[playground/src/sim/sim_mem.scala 16:16]
  output [3:0]  io_memAxi_wr_bits_id, // @[playground/src/sim/sim_mem.scala 16:16]
  output [1:0]  io_memAxi_wr_bits_resp, // @[playground/src/sim/sim_mem.scala 16:16]
  output        io_memAxi_ra_ready, // @[playground/src/sim/sim_mem.scala 16:16]
  input         io_memAxi_ra_valid, // @[playground/src/sim/sim_mem.scala 16:16]
  input  [3:0]  io_memAxi_ra_bits_id, // @[playground/src/sim/sim_mem.scala 16:16]
  input  [31:0] io_memAxi_ra_bits_addr, // @[playground/src/sim/sim_mem.scala 16:16]
  input  [7:0]  io_memAxi_ra_bits_len, // @[playground/src/sim/sim_mem.scala 16:16]
  input  [2:0]  io_memAxi_ra_bits_size, // @[playground/src/sim/sim_mem.scala 16:16]
  input  [1:0]  io_memAxi_ra_bits_burst, // @[playground/src/sim/sim_mem.scala 16:16]
  input         io_memAxi_rd_ready, // @[playground/src/sim/sim_mem.scala 16:16]
  output        io_memAxi_rd_valid, // @[playground/src/sim/sim_mem.scala 16:16]
  output [3:0]  io_memAxi_rd_bits_id, // @[playground/src/sim/sim_mem.scala 16:16]
  output [63:0] io_memAxi_rd_bits_data, // @[playground/src/sim/sim_mem.scala 16:16]
  output [1:0]  io_memAxi_rd_bits_resp, // @[playground/src/sim/sim_mem.scala 16:16]
  output        io_memAxi_rd_bits_last // @[playground/src/sim/sim_mem.scala 16:16]
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
`endif // RANDOMIZE_REG_INIT
  reg /* sparse */ [7:0] ram [0:268435455]; // @[playground/src/sim/sim_mem.scala 18:18]
  wire  ram_rdata_MPORT_en; // @[playground/src/sim/sim_mem.scala 18:18]
  wire [27:0] ram_rdata_MPORT_addr; // @[playground/src/sim/sim_mem.scala 18:18]
  wire [7:0] ram_rdata_MPORT_data; // @[playground/src/sim/sim_mem.scala 18:18]
  wire  ram_rdata_MPORT_1_en; // @[playground/src/sim/sim_mem.scala 18:18]
  wire [27:0] ram_rdata_MPORT_1_addr; // @[playground/src/sim/sim_mem.scala 18:18]
  wire [7:0] ram_rdata_MPORT_1_data; // @[playground/src/sim/sim_mem.scala 18:18]
  wire  ram_rdata_MPORT_2_en; // @[playground/src/sim/sim_mem.scala 18:18]
  wire [27:0] ram_rdata_MPORT_2_addr; // @[playground/src/sim/sim_mem.scala 18:18]
  wire [7:0] ram_rdata_MPORT_2_data; // @[playground/src/sim/sim_mem.scala 18:18]
  wire  ram_rdata_MPORT_3_en; // @[playground/src/sim/sim_mem.scala 18:18]
  wire [27:0] ram_rdata_MPORT_3_addr; // @[playground/src/sim/sim_mem.scala 18:18]
  wire [7:0] ram_rdata_MPORT_3_data; // @[playground/src/sim/sim_mem.scala 18:18]
  wire  ram_rdata_MPORT_4_en; // @[playground/src/sim/sim_mem.scala 18:18]
  wire [27:0] ram_rdata_MPORT_4_addr; // @[playground/src/sim/sim_mem.scala 18:18]
  wire [7:0] ram_rdata_MPORT_4_data; // @[playground/src/sim/sim_mem.scala 18:18]
  wire  ram_rdata_MPORT_5_en; // @[playground/src/sim/sim_mem.scala 18:18]
  wire [27:0] ram_rdata_MPORT_5_addr; // @[playground/src/sim/sim_mem.scala 18:18]
  wire [7:0] ram_rdata_MPORT_5_data; // @[playground/src/sim/sim_mem.scala 18:18]
  wire  ram_rdata_MPORT_6_en; // @[playground/src/sim/sim_mem.scala 18:18]
  wire [27:0] ram_rdata_MPORT_6_addr; // @[playground/src/sim/sim_mem.scala 18:18]
  wire [7:0] ram_rdata_MPORT_6_data; // @[playground/src/sim/sim_mem.scala 18:18]
  wire  ram_rdata_MPORT_7_en; // @[playground/src/sim/sim_mem.scala 18:18]
  wire [27:0] ram_rdata_MPORT_7_addr; // @[playground/src/sim/sim_mem.scala 18:18]
  wire [7:0] ram_rdata_MPORT_7_data; // @[playground/src/sim/sim_mem.scala 18:18]
  wire  ram_MPORT_1_en; // @[playground/src/sim/sim_mem.scala 18:18]
  wire [27:0] ram_MPORT_1_addr; // @[playground/src/sim/sim_mem.scala 18:18]
  wire [7:0] ram_MPORT_1_data; // @[playground/src/sim/sim_mem.scala 18:18]
  wire  ram_MPORT_3_en; // @[playground/src/sim/sim_mem.scala 18:18]
  wire [27:0] ram_MPORT_3_addr; // @[playground/src/sim/sim_mem.scala 18:18]
  wire [7:0] ram_MPORT_3_data; // @[playground/src/sim/sim_mem.scala 18:18]
  wire  ram_MPORT_5_en; // @[playground/src/sim/sim_mem.scala 18:18]
  wire [27:0] ram_MPORT_5_addr; // @[playground/src/sim/sim_mem.scala 18:18]
  wire [7:0] ram_MPORT_5_data; // @[playground/src/sim/sim_mem.scala 18:18]
  wire  ram_MPORT_7_en; // @[playground/src/sim/sim_mem.scala 18:18]
  wire [27:0] ram_MPORT_7_addr; // @[playground/src/sim/sim_mem.scala 18:18]
  wire [7:0] ram_MPORT_7_data; // @[playground/src/sim/sim_mem.scala 18:18]
  wire  ram_MPORT_9_en; // @[playground/src/sim/sim_mem.scala 18:18]
  wire [27:0] ram_MPORT_9_addr; // @[playground/src/sim/sim_mem.scala 18:18]
  wire [7:0] ram_MPORT_9_data; // @[playground/src/sim/sim_mem.scala 18:18]
  wire  ram_MPORT_11_en; // @[playground/src/sim/sim_mem.scala 18:18]
  wire [27:0] ram_MPORT_11_addr; // @[playground/src/sim/sim_mem.scala 18:18]
  wire [7:0] ram_MPORT_11_data; // @[playground/src/sim/sim_mem.scala 18:18]
  wire  ram_MPORT_13_en; // @[playground/src/sim/sim_mem.scala 18:18]
  wire [27:0] ram_MPORT_13_addr; // @[playground/src/sim/sim_mem.scala 18:18]
  wire [7:0] ram_MPORT_13_data; // @[playground/src/sim/sim_mem.scala 18:18]
  wire  ram_MPORT_15_en; // @[playground/src/sim/sim_mem.scala 18:18]
  wire [27:0] ram_MPORT_15_addr; // @[playground/src/sim/sim_mem.scala 18:18]
  wire [7:0] ram_MPORT_15_data; // @[playground/src/sim/sim_mem.scala 18:18]
  wire [7:0] ram_MPORT_data; // @[playground/src/sim/sim_mem.scala 18:18]
  wire [27:0] ram_MPORT_addr; // @[playground/src/sim/sim_mem.scala 18:18]
  wire  ram_MPORT_mask; // @[playground/src/sim/sim_mem.scala 18:18]
  wire  ram_MPORT_en; // @[playground/src/sim/sim_mem.scala 18:18]
  wire [7:0] ram_MPORT_2_data; // @[playground/src/sim/sim_mem.scala 18:18]
  wire [27:0] ram_MPORT_2_addr; // @[playground/src/sim/sim_mem.scala 18:18]
  wire  ram_MPORT_2_mask; // @[playground/src/sim/sim_mem.scala 18:18]
  wire  ram_MPORT_2_en; // @[playground/src/sim/sim_mem.scala 18:18]
  wire [7:0] ram_MPORT_4_data; // @[playground/src/sim/sim_mem.scala 18:18]
  wire [27:0] ram_MPORT_4_addr; // @[playground/src/sim/sim_mem.scala 18:18]
  wire  ram_MPORT_4_mask; // @[playground/src/sim/sim_mem.scala 18:18]
  wire  ram_MPORT_4_en; // @[playground/src/sim/sim_mem.scala 18:18]
  wire [7:0] ram_MPORT_6_data; // @[playground/src/sim/sim_mem.scala 18:18]
  wire [27:0] ram_MPORT_6_addr; // @[playground/src/sim/sim_mem.scala 18:18]
  wire  ram_MPORT_6_mask; // @[playground/src/sim/sim_mem.scala 18:18]
  wire  ram_MPORT_6_en; // @[playground/src/sim/sim_mem.scala 18:18]
  wire [7:0] ram_MPORT_8_data; // @[playground/src/sim/sim_mem.scala 18:18]
  wire [27:0] ram_MPORT_8_addr; // @[playground/src/sim/sim_mem.scala 18:18]
  wire  ram_MPORT_8_mask; // @[playground/src/sim/sim_mem.scala 18:18]
  wire  ram_MPORT_8_en; // @[playground/src/sim/sim_mem.scala 18:18]
  wire [7:0] ram_MPORT_10_data; // @[playground/src/sim/sim_mem.scala 18:18]
  wire [27:0] ram_MPORT_10_addr; // @[playground/src/sim/sim_mem.scala 18:18]
  wire  ram_MPORT_10_mask; // @[playground/src/sim/sim_mem.scala 18:18]
  wire  ram_MPORT_10_en; // @[playground/src/sim/sim_mem.scala 18:18]
  wire [7:0] ram_MPORT_12_data; // @[playground/src/sim/sim_mem.scala 18:18]
  wire [27:0] ram_MPORT_12_addr; // @[playground/src/sim/sim_mem.scala 18:18]
  wire  ram_MPORT_12_mask; // @[playground/src/sim/sim_mem.scala 18:18]
  wire  ram_MPORT_12_en; // @[playground/src/sim/sim_mem.scala 18:18]
  wire [7:0] ram_MPORT_14_data; // @[playground/src/sim/sim_mem.scala 18:18]
  wire [27:0] ram_MPORT_14_addr; // @[playground/src/sim/sim_mem.scala 18:18]
  wire  ram_MPORT_14_mask; // @[playground/src/sim/sim_mem.scala 18:18]
  wire  ram_MPORT_14_en; // @[playground/src/sim/sim_mem.scala 18:18]
  reg [7:0] burstLen; // @[playground/src/sim/sim_mem.scala 20:27]
  reg [7:0] offset; // @[playground/src/sim/sim_mem.scala 21:26]
  reg  waReady; // @[playground/src/sim/sim_mem.scala 23:26]
  reg  wdReady; // @[playground/src/sim/sim_mem.scala 24:26]
  reg [31:0] waStart; // @[playground/src/sim/sim_mem.scala 25:26]
  wire [11:0] _waddr_T = offset * 4'h8; // @[playground/src/sim/sim_mem.scala 27:37]
  wire [31:0] _GEN_116 = {{20'd0}, _waddr_T}; // @[playground/src/sim/sim_mem.scala 27:28]
  wire [31:0] _waddr_T_2 = waStart + _GEN_116; // @[playground/src/sim/sim_mem.scala 27:28]
  wire [31:0] waddr = _waddr_T_2 & 32'hfffffff; // @[playground/src/sim/sim_mem.scala 27:44]
  reg  raReady; // @[playground/src/sim/sim_mem.scala 29:26]
  reg [31:0] raStart; // @[playground/src/sim/sim_mem.scala 30:26]
  reg  rdValid; // @[playground/src/sim/sim_mem.scala 31:26]
  wire [31:0] _rdata_T_2 = raStart + _GEN_116; // @[playground/src/sim/sim_mem.scala 32:65]
  wire [31:0] _rdata_T_4 = _rdata_T_2 + 32'h7; // @[playground/src/sim/sim_mem.scala 32:80]
  wire [31:0] _rdata_T_5 = _rdata_T_4 & 32'hfffffff; // @[playground/src/sim/sim_mem.scala 32:86]
  wire [31:0] _rdata_T_11 = _rdata_T_2 + 32'h6; // @[playground/src/sim/sim_mem.scala 32:80]
  wire [31:0] _rdata_T_12 = _rdata_T_11 & 32'hfffffff; // @[playground/src/sim/sim_mem.scala 32:86]
  wire [31:0] _rdata_T_18 = _rdata_T_2 + 32'h5; // @[playground/src/sim/sim_mem.scala 32:80]
  wire [31:0] _rdata_T_19 = _rdata_T_18 & 32'hfffffff; // @[playground/src/sim/sim_mem.scala 32:86]
  wire [31:0] _rdata_T_25 = _rdata_T_2 + 32'h4; // @[playground/src/sim/sim_mem.scala 32:80]
  wire [31:0] _rdata_T_26 = _rdata_T_25 & 32'hfffffff; // @[playground/src/sim/sim_mem.scala 32:86]
  wire [31:0] _rdata_T_32 = _rdata_T_2 + 32'h3; // @[playground/src/sim/sim_mem.scala 32:80]
  wire [31:0] _rdata_T_33 = _rdata_T_32 & 32'hfffffff; // @[playground/src/sim/sim_mem.scala 32:86]
  wire [31:0] _rdata_T_39 = _rdata_T_2 + 32'h2; // @[playground/src/sim/sim_mem.scala 32:80]
  wire [31:0] _rdata_T_40 = _rdata_T_39 & 32'hfffffff; // @[playground/src/sim/sim_mem.scala 32:86]
  wire [31:0] _rdata_T_46 = _rdata_T_2 + 32'h1; // @[playground/src/sim/sim_mem.scala 32:80]
  wire [31:0] _rdata_T_47 = _rdata_T_46 & 32'hfffffff; // @[playground/src/sim/sim_mem.scala 32:86]
  wire [32:0] _rdata_T_52 = {{1'd0}, _rdata_T_2}; // @[playground/src/sim/sim_mem.scala 32:80]
  wire [31:0] _rdata_T_54 = _rdata_T_52[31:0] & 32'hfffffff; // @[playground/src/sim/sim_mem.scala 32:86]
  wire [31:0] rdata_lo = {ram_rdata_MPORT_4_data,ram_rdata_MPORT_5_data,ram_rdata_MPORT_6_data,ram_rdata_MPORT_7_data}; // @[playground/src/sim/sim_mem.scala 32:22]
  wire [31:0] rdata_hi = {ram_rdata_MPORT_data,ram_rdata_MPORT_1_data,ram_rdata_MPORT_2_data,ram_rdata_MPORT_3_data}; // @[playground/src/sim/sim_mem.scala 32:22]
  reg [1:0] state; // @[playground/src/sim/sim_mem.scala 34:24]
  wire  isLast = offset >= burstLen; // @[playground/src/sim/sim_mem.scala 36:27]
  wire  _T = 2'h0 == state; // @[playground/src/sim/sim_mem.scala 38:18]
  wire  _GEN_4 = io_memAxi_wa_valid & waReady | wdReady; // @[playground/src/sim/sim_mem.scala 43:48 48:25 24:26]
  wire  _GEN_9 = io_memAxi_ra_valid & raReady | rdValid; // @[playground/src/sim/sim_mem.scala 50:48 55:25 31:26]
  wire [32:0] _T_4 = {{1'd0}, waddr}; // @[playground/src/sim/sim_mem.scala 62:35]
  wire [31:0] _T_15 = waddr + 32'h1; // @[playground/src/sim/sim_mem.scala 62:35]
  wire [31:0] _T_25 = waddr + 32'h2; // @[playground/src/sim/sim_mem.scala 62:35]
  wire [31:0] _T_35 = waddr + 32'h3; // @[playground/src/sim/sim_mem.scala 62:35]
  wire [31:0] _T_45 = waddr + 32'h4; // @[playground/src/sim/sim_mem.scala 62:35]
  wire [31:0] _T_55 = waddr + 32'h5; // @[playground/src/sim/sim_mem.scala 62:35]
  wire [31:0] _T_65 = waddr + 32'h6; // @[playground/src/sim/sim_mem.scala 62:35]
  wire [31:0] _T_75 = waddr + 32'h7; // @[playground/src/sim/sim_mem.scala 62:35]
  wire [7:0] _offset_T_1 = offset + 8'h1; // @[playground/src/sim/sim_mem.scala 65:34]
  wire  _GEN_10 = io_memAxi_wd_bits_last ? 1'h0 : wdReady; // @[playground/src/sim/sim_mem.scala 24:26 66:45 67:29]
  wire [1:0] _GEN_11 = io_memAxi_wd_bits_last ? 2'h0 : state; // @[playground/src/sim/sim_mem.scala 34:24 66:45 68:29]
  wire [1:0] _GEN_42 = isLast ? 2'h0 : state; // @[playground/src/sim/sim_mem.scala 34:24 78:29 79:27]
  wire [7:0] _GEN_43 = rdValid & io_memAxi_rd_ready ? _offset_T_1 : offset; // @[playground/src/sim/sim_mem.scala 75:48 76:25 21:26]
  wire  _GEN_44 = rdValid & io_memAxi_rd_ready ? 1'h0 : 1'h1; // @[playground/src/sim/sim_mem.scala 74:21 75:48 77:25]
  wire [1:0] _GEN_45 = rdValid & io_memAxi_rd_ready ? _GEN_42 : state; // @[playground/src/sim/sim_mem.scala 34:24 75:48]
  wire  _GEN_51 = 2'h1 == state & io_memAxi_wd_valid; // @[playground/src/sim/sim_mem.scala 18:18 38:18]
  assign ram_rdata_MPORT_en = 1'h1;
  assign ram_rdata_MPORT_addr = _rdata_T_5[27:0];
  assign ram_rdata_MPORT_data = ram[ram_rdata_MPORT_addr]; // @[playground/src/sim/sim_mem.scala 18:18]
  assign ram_rdata_MPORT_1_en = 1'h1;
  assign ram_rdata_MPORT_1_addr = _rdata_T_12[27:0];
  assign ram_rdata_MPORT_1_data = ram[ram_rdata_MPORT_1_addr]; // @[playground/src/sim/sim_mem.scala 18:18]
  assign ram_rdata_MPORT_2_en = 1'h1;
  assign ram_rdata_MPORT_2_addr = _rdata_T_19[27:0];
  assign ram_rdata_MPORT_2_data = ram[ram_rdata_MPORT_2_addr]; // @[playground/src/sim/sim_mem.scala 18:18]
  assign ram_rdata_MPORT_3_en = 1'h1;
  assign ram_rdata_MPORT_3_addr = _rdata_T_26[27:0];
  assign ram_rdata_MPORT_3_data = ram[ram_rdata_MPORT_3_addr]; // @[playground/src/sim/sim_mem.scala 18:18]
  assign ram_rdata_MPORT_4_en = 1'h1;
  assign ram_rdata_MPORT_4_addr = _rdata_T_33[27:0];
  assign ram_rdata_MPORT_4_data = ram[ram_rdata_MPORT_4_addr]; // @[playground/src/sim/sim_mem.scala 18:18]
  assign ram_rdata_MPORT_5_en = 1'h1;
  assign ram_rdata_MPORT_5_addr = _rdata_T_40[27:0];
  assign ram_rdata_MPORT_5_data = ram[ram_rdata_MPORT_5_addr]; // @[playground/src/sim/sim_mem.scala 18:18]
  assign ram_rdata_MPORT_6_en = 1'h1;
  assign ram_rdata_MPORT_6_addr = _rdata_T_47[27:0];
  assign ram_rdata_MPORT_6_data = ram[ram_rdata_MPORT_6_addr]; // @[playground/src/sim/sim_mem.scala 18:18]
  assign ram_rdata_MPORT_7_en = 1'h1;
  assign ram_rdata_MPORT_7_addr = _rdata_T_54[27:0];
  assign ram_rdata_MPORT_7_data = ram[ram_rdata_MPORT_7_addr]; // @[playground/src/sim/sim_mem.scala 18:18]
  assign ram_MPORT_1_en = _T ? 1'h0 : _GEN_51;
  assign ram_MPORT_1_addr = _T_4[27:0];
  assign ram_MPORT_1_data = ram[ram_MPORT_1_addr]; // @[playground/src/sim/sim_mem.scala 18:18]
  assign ram_MPORT_3_en = _T ? 1'h0 : _GEN_51;
  assign ram_MPORT_3_addr = _T_15[27:0];
  assign ram_MPORT_3_data = ram[ram_MPORT_3_addr]; // @[playground/src/sim/sim_mem.scala 18:18]
  assign ram_MPORT_5_en = _T ? 1'h0 : _GEN_51;
  assign ram_MPORT_5_addr = _T_25[27:0];
  assign ram_MPORT_5_data = ram[ram_MPORT_5_addr]; // @[playground/src/sim/sim_mem.scala 18:18]
  assign ram_MPORT_7_en = _T ? 1'h0 : _GEN_51;
  assign ram_MPORT_7_addr = _T_35[27:0];
  assign ram_MPORT_7_data = ram[ram_MPORT_7_addr]; // @[playground/src/sim/sim_mem.scala 18:18]
  assign ram_MPORT_9_en = _T ? 1'h0 : _GEN_51;
  assign ram_MPORT_9_addr = _T_45[27:0];
  assign ram_MPORT_9_data = ram[ram_MPORT_9_addr]; // @[playground/src/sim/sim_mem.scala 18:18]
  assign ram_MPORT_11_en = _T ? 1'h0 : _GEN_51;
  assign ram_MPORT_11_addr = _T_55[27:0];
  assign ram_MPORT_11_data = ram[ram_MPORT_11_addr]; // @[playground/src/sim/sim_mem.scala 18:18]
  assign ram_MPORT_13_en = _T ? 1'h0 : _GEN_51;
  assign ram_MPORT_13_addr = _T_65[27:0];
  assign ram_MPORT_13_data = ram[ram_MPORT_13_addr]; // @[playground/src/sim/sim_mem.scala 18:18]
  assign ram_MPORT_15_en = _T ? 1'h0 : _GEN_51;
  assign ram_MPORT_15_addr = _T_75[27:0];
  assign ram_MPORT_15_data = ram[ram_MPORT_15_addr]; // @[playground/src/sim/sim_mem.scala 18:18]
  assign ram_MPORT_data = io_memAxi_wd_bits_strb[0] ? io_memAxi_wd_bits_data[7:0] : ram_MPORT_1_data;
  assign ram_MPORT_addr = _T_4[27:0];
  assign ram_MPORT_mask = 1'h1;
  assign ram_MPORT_en = _T ? 1'h0 : _GEN_51;
  assign ram_MPORT_2_data = io_memAxi_wd_bits_strb[1] ? io_memAxi_wd_bits_data[15:8] : ram_MPORT_3_data;
  assign ram_MPORT_2_addr = _T_15[27:0];
  assign ram_MPORT_2_mask = 1'h1;
  assign ram_MPORT_2_en = _T ? 1'h0 : _GEN_51;
  assign ram_MPORT_4_data = io_memAxi_wd_bits_strb[2] ? io_memAxi_wd_bits_data[23:16] : ram_MPORT_5_data;
  assign ram_MPORT_4_addr = _T_25[27:0];
  assign ram_MPORT_4_mask = 1'h1;
  assign ram_MPORT_4_en = _T ? 1'h0 : _GEN_51;
  assign ram_MPORT_6_data = io_memAxi_wd_bits_strb[3] ? io_memAxi_wd_bits_data[31:24] : ram_MPORT_7_data;
  assign ram_MPORT_6_addr = _T_35[27:0];
  assign ram_MPORT_6_mask = 1'h1;
  assign ram_MPORT_6_en = _T ? 1'h0 : _GEN_51;
  assign ram_MPORT_8_data = io_memAxi_wd_bits_strb[4] ? io_memAxi_wd_bits_data[39:32] : ram_MPORT_9_data;
  assign ram_MPORT_8_addr = _T_45[27:0];
  assign ram_MPORT_8_mask = 1'h1;
  assign ram_MPORT_8_en = _T ? 1'h0 : _GEN_51;
  assign ram_MPORT_10_data = io_memAxi_wd_bits_strb[5] ? io_memAxi_wd_bits_data[47:40] : ram_MPORT_11_data;
  assign ram_MPORT_10_addr = _T_55[27:0];
  assign ram_MPORT_10_mask = 1'h1;
  assign ram_MPORT_10_en = _T ? 1'h0 : _GEN_51;
  assign ram_MPORT_12_data = io_memAxi_wd_bits_strb[6] ? io_memAxi_wd_bits_data[55:48] : ram_MPORT_13_data;
  assign ram_MPORT_12_addr = _T_65[27:0];
  assign ram_MPORT_12_mask = 1'h1;
  assign ram_MPORT_12_en = _T ? 1'h0 : _GEN_51;
  assign ram_MPORT_14_data = io_memAxi_wd_bits_strb[7] ? io_memAxi_wd_bits_data[63:56] : ram_MPORT_15_data;
  assign ram_MPORT_14_addr = _T_75[27:0];
  assign ram_MPORT_14_mask = 1'h1;
  assign ram_MPORT_14_en = _T ? 1'h0 : _GEN_51;
  assign io_memAxi_wa_ready = waReady; // @[playground/src/sim/sim_mem.scala 89:24]
  assign io_memAxi_wd_ready = wdReady; // @[playground/src/sim/sim_mem.scala 90:24]
  assign io_memAxi_wr_valid = 1'h1; // @[playground/src/sim/sim_mem.scala 87:24]
  assign io_memAxi_wr_bits_id = 4'h0; // @[playground/src/axi/axi.scala 58:{38,38}]
  assign io_memAxi_wr_bits_resp = 2'h0; // @[playground/src/sim/sim_mem.scala 88:28]
  assign io_memAxi_ra_ready = raReady; // @[playground/src/sim/sim_mem.scala 91:24]
  assign io_memAxi_rd_valid = rdValid; // @[playground/src/sim/sim_mem.scala 92:24]
  assign io_memAxi_rd_bits_id = 4'h0; // @[playground/src/axi/axi.scala 68:{38,38}]
  assign io_memAxi_rd_bits_data = {rdata_hi,rdata_lo}; // @[playground/src/sim/sim_mem.scala 32:22]
  assign io_memAxi_rd_bits_resp = 2'h0; // @[playground/src/axi/axi.scala 68:{38,38}]
  assign io_memAxi_rd_bits_last = offset >= burstLen; // @[playground/src/sim/sim_mem.scala 36:27]
  always @(posedge clock) begin
    if (ram_MPORT_en & ram_MPORT_mask) begin
      ram[ram_MPORT_addr] <= ram_MPORT_data; // @[playground/src/sim/sim_mem.scala 18:18]
    end
    if (ram_MPORT_2_en & ram_MPORT_2_mask) begin
      ram[ram_MPORT_2_addr] <= ram_MPORT_2_data; // @[playground/src/sim/sim_mem.scala 18:18]
    end
    if (ram_MPORT_4_en & ram_MPORT_4_mask) begin
      ram[ram_MPORT_4_addr] <= ram_MPORT_4_data; // @[playground/src/sim/sim_mem.scala 18:18]
    end
    if (ram_MPORT_6_en & ram_MPORT_6_mask) begin
      ram[ram_MPORT_6_addr] <= ram_MPORT_6_data; // @[playground/src/sim/sim_mem.scala 18:18]
    end
    if (ram_MPORT_8_en & ram_MPORT_8_mask) begin
      ram[ram_MPORT_8_addr] <= ram_MPORT_8_data; // @[playground/src/sim/sim_mem.scala 18:18]
    end
    if (ram_MPORT_10_en & ram_MPORT_10_mask) begin
      ram[ram_MPORT_10_addr] <= ram_MPORT_10_data; // @[playground/src/sim/sim_mem.scala 18:18]
    end
    if (ram_MPORT_12_en & ram_MPORT_12_mask) begin
      ram[ram_MPORT_12_addr] <= ram_MPORT_12_data; // @[playground/src/sim/sim_mem.scala 18:18]
    end
    if (ram_MPORT_14_en & ram_MPORT_14_mask) begin
      ram[ram_MPORT_14_addr] <= ram_MPORT_14_data; // @[playground/src/sim/sim_mem.scala 18:18]
    end
    if (reset) begin // @[playground/src/sim/sim_mem.scala 20:27]
      burstLen <= 8'h0; // @[playground/src/sim/sim_mem.scala 20:27]
    end else if (2'h0 == state) begin // @[playground/src/sim/sim_mem.scala 38:18]
      if (io_memAxi_ra_valid & raReady) begin // @[playground/src/sim/sim_mem.scala 50:48]
        burstLen <= io_memAxi_ra_bits_len; // @[playground/src/sim/sim_mem.scala 53:26]
      end else if (io_memAxi_wa_valid & waReady) begin // @[playground/src/sim/sim_mem.scala 43:48]
        burstLen <= io_memAxi_wa_bits_len; // @[playground/src/sim/sim_mem.scala 46:26]
      end
    end
    if (reset) begin // @[playground/src/sim/sim_mem.scala 21:26]
      offset <= 8'h0; // @[playground/src/sim/sim_mem.scala 21:26]
    end else if (2'h0 == state) begin // @[playground/src/sim/sim_mem.scala 38:18]
      offset <= 8'h0; // @[playground/src/sim/sim_mem.scala 42:21]
    end else if (2'h1 == state) begin // @[playground/src/sim/sim_mem.scala 38:18]
      if (io_memAxi_wd_valid) begin // @[playground/src/sim/sim_mem.scala 60:37]
        offset <= _offset_T_1; // @[playground/src/sim/sim_mem.scala 65:24]
      end
    end else if (2'h3 == state) begin // @[playground/src/sim/sim_mem.scala 38:18]
      offset <= _GEN_43;
    end
    if (reset) begin // @[playground/src/sim/sim_mem.scala 23:26]
      waReady <= 1'h0; // @[playground/src/sim/sim_mem.scala 23:26]
    end else if (2'h0 == state) begin // @[playground/src/sim/sim_mem.scala 38:18]
      if (io_memAxi_wa_valid & waReady) begin // @[playground/src/sim/sim_mem.scala 43:48]
        waReady <= 1'h0; // @[playground/src/sim/sim_mem.scala 47:25]
      end else begin
        waReady <= 1'h1; // @[playground/src/sim/sim_mem.scala 40:21]
      end
    end
    if (reset) begin // @[playground/src/sim/sim_mem.scala 24:26]
      wdReady <= 1'h0; // @[playground/src/sim/sim_mem.scala 24:26]
    end else if (2'h0 == state) begin // @[playground/src/sim/sim_mem.scala 38:18]
      wdReady <= _GEN_4;
    end else if (2'h1 == state) begin // @[playground/src/sim/sim_mem.scala 38:18]
      if (io_memAxi_wd_valid) begin // @[playground/src/sim/sim_mem.scala 60:37]
        wdReady <= _GEN_10;
      end
    end
    if (reset) begin // @[playground/src/sim/sim_mem.scala 25:26]
      waStart <= 32'h0; // @[playground/src/sim/sim_mem.scala 25:26]
    end else if (2'h0 == state) begin // @[playground/src/sim/sim_mem.scala 38:18]
      if (io_memAxi_wa_valid & waReady) begin // @[playground/src/sim/sim_mem.scala 43:48]
        waStart <= io_memAxi_wa_bits_addr; // @[playground/src/sim/sim_mem.scala 45:27]
      end
    end
    if (reset) begin // @[playground/src/sim/sim_mem.scala 29:26]
      raReady <= 1'h0; // @[playground/src/sim/sim_mem.scala 29:26]
    end else if (2'h0 == state) begin // @[playground/src/sim/sim_mem.scala 38:18]
      if (io_memAxi_ra_valid & raReady) begin // @[playground/src/sim/sim_mem.scala 50:48]
        raReady <= 1'h0; // @[playground/src/sim/sim_mem.scala 54:25]
      end else begin
        raReady <= 1'h1; // @[playground/src/sim/sim_mem.scala 41:21]
      end
    end
    if (reset) begin // @[playground/src/sim/sim_mem.scala 30:26]
      raStart <= 32'h0; // @[playground/src/sim/sim_mem.scala 30:26]
    end else if (2'h0 == state) begin // @[playground/src/sim/sim_mem.scala 38:18]
      if (io_memAxi_ra_valid & raReady) begin // @[playground/src/sim/sim_mem.scala 50:48]
        raStart <= io_memAxi_ra_bits_addr; // @[playground/src/sim/sim_mem.scala 52:27]
      end
    end
    if (reset) begin // @[playground/src/sim/sim_mem.scala 31:26]
      rdValid <= 1'h0; // @[playground/src/sim/sim_mem.scala 31:26]
    end else if (2'h0 == state) begin // @[playground/src/sim/sim_mem.scala 38:18]
      rdValid <= _GEN_9;
    end else if (!(2'h1 == state)) begin // @[playground/src/sim/sim_mem.scala 38:18]
      if (2'h3 == state) begin // @[playground/src/sim/sim_mem.scala 38:18]
        rdValid <= _GEN_44;
      end
    end
    if (reset) begin // @[playground/src/sim/sim_mem.scala 34:24]
      state <= 2'h0; // @[playground/src/sim/sim_mem.scala 34:24]
    end else if (2'h0 == state) begin // @[playground/src/sim/sim_mem.scala 38:18]
      if (io_memAxi_ra_valid & raReady) begin // @[playground/src/sim/sim_mem.scala 50:48]
        state <= 2'h3; // @[playground/src/sim/sim_mem.scala 51:25]
      end else if (io_memAxi_wa_valid & waReady) begin // @[playground/src/sim/sim_mem.scala 43:48]
        state <= 2'h1; // @[playground/src/sim/sim_mem.scala 44:25]
      end
    end else if (2'h1 == state) begin // @[playground/src/sim/sim_mem.scala 38:18]
      if (io_memAxi_wd_valid) begin // @[playground/src/sim/sim_mem.scala 60:37]
        state <= _GEN_11;
      end
    end else if (2'h3 == state) begin // @[playground/src/sim/sim_mem.scala 38:18]
      state <= _GEN_45;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 268435456; initvar = initvar+1)
    ram[initvar] = _RAND_0[7:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  burstLen = _RAND_1[7:0];
  _RAND_2 = {1{`RANDOM}};
  offset = _RAND_2[7:0];
  _RAND_3 = {1{`RANDOM}};
  waReady = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  wdReady = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  waStart = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  raReady = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  raStart = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  rdValid = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  state = _RAND_9[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module SimMMIO(
  input         clock,
  input         reset,
  output        io_mmioAxi_wa_ready, // @[playground/src/sim/sim_mmio.scala 45:16]
  input         io_mmioAxi_wa_valid, // @[playground/src/sim/sim_mmio.scala 45:16]
  input  [31:0] io_mmioAxi_wa_bits_addr, // @[playground/src/sim/sim_mmio.scala 45:16]
  output        io_mmioAxi_wd_ready, // @[playground/src/sim/sim_mmio.scala 45:16]
  input         io_mmioAxi_wd_valid, // @[playground/src/sim/sim_mmio.scala 45:16]
  input  [63:0] io_mmioAxi_wd_bits_data, // @[playground/src/sim/sim_mmio.scala 45:16]
  input  [7:0]  io_mmioAxi_wd_bits_strb, // @[playground/src/sim/sim_mmio.scala 45:16]
  input         io_mmioAxi_wd_bits_last, // @[playground/src/sim/sim_mmio.scala 45:16]
  output        io_mmioAxi_ra_ready, // @[playground/src/sim/sim_mmio.scala 45:16]
  input         io_mmioAxi_ra_valid, // @[playground/src/sim/sim_mmio.scala 45:16]
  input  [31:0] io_mmioAxi_ra_bits_addr, // @[playground/src/sim/sim_mmio.scala 45:16]
  input         io_mmioAxi_rd_ready, // @[playground/src/sim/sim_mmio.scala 45:16]
  output        io_mmioAxi_rd_valid, // @[playground/src/sim/sim_mmio.scala 45:16]
  output [63:0] io_mmioAxi_rd_bits_data, // @[playground/src/sim/sim_mmio.scala 45:16]
  output        io_mmioAxi_rd_bits_last // @[playground/src/sim/sim_mmio.scala 45:16]
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [63:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
`endif // RANDOMIZE_REG_INIT
  wire [6:0] sdcard_addr; // @[playground/src/sim/sim_mmio.scala 46:24]
  wire  sdcard_wen; // @[playground/src/sim/sim_mmio.scala 46:24]
  wire [63:0] sdcard_wdata; // @[playground/src/sim/sim_mmio.scala 46:24]
  wire  sdcard_clock; // @[playground/src/sim/sim_mmio.scala 46:24]
  wire  sdcard_cen; // @[playground/src/sim/sim_mmio.scala 46:24]
  wire [63:0] sdcard_rdata; // @[playground/src/sim/sim_mmio.scala 46:24]
  reg [7:0] disk [0:67108863]; // @[playground/src/sim/sim_mmio.scala 55:19]
  wire  disk_disk_rdata_MPORT_en; // @[playground/src/sim/sim_mmio.scala 55:19]
  wire [25:0] disk_disk_rdata_MPORT_addr; // @[playground/src/sim/sim_mmio.scala 55:19]
  wire [7:0] disk_disk_rdata_MPORT_data; // @[playground/src/sim/sim_mmio.scala 55:19]
  wire  disk_disk_rdata_MPORT_1_en; // @[playground/src/sim/sim_mmio.scala 55:19]
  wire [25:0] disk_disk_rdata_MPORT_1_addr; // @[playground/src/sim/sim_mmio.scala 55:19]
  wire [7:0] disk_disk_rdata_MPORT_1_data; // @[playground/src/sim/sim_mmio.scala 55:19]
  wire  disk_disk_rdata_MPORT_2_en; // @[playground/src/sim/sim_mmio.scala 55:19]
  wire [25:0] disk_disk_rdata_MPORT_2_addr; // @[playground/src/sim/sim_mmio.scala 55:19]
  wire [7:0] disk_disk_rdata_MPORT_2_data; // @[playground/src/sim/sim_mmio.scala 55:19]
  wire  disk_disk_rdata_MPORT_3_en; // @[playground/src/sim/sim_mmio.scala 55:19]
  wire [25:0] disk_disk_rdata_MPORT_3_addr; // @[playground/src/sim/sim_mmio.scala 55:19]
  wire [7:0] disk_disk_rdata_MPORT_3_data; // @[playground/src/sim/sim_mmio.scala 55:19]
  wire  disk_disk_rdata_MPORT_4_en; // @[playground/src/sim/sim_mmio.scala 55:19]
  wire [25:0] disk_disk_rdata_MPORT_4_addr; // @[playground/src/sim/sim_mmio.scala 55:19]
  wire [7:0] disk_disk_rdata_MPORT_4_data; // @[playground/src/sim/sim_mmio.scala 55:19]
  wire  disk_disk_rdata_MPORT_5_en; // @[playground/src/sim/sim_mmio.scala 55:19]
  wire [25:0] disk_disk_rdata_MPORT_5_addr; // @[playground/src/sim/sim_mmio.scala 55:19]
  wire [7:0] disk_disk_rdata_MPORT_5_data; // @[playground/src/sim/sim_mmio.scala 55:19]
  wire  disk_disk_rdata_MPORT_6_en; // @[playground/src/sim/sim_mmio.scala 55:19]
  wire [25:0] disk_disk_rdata_MPORT_6_addr; // @[playground/src/sim/sim_mmio.scala 55:19]
  wire [7:0] disk_disk_rdata_MPORT_6_data; // @[playground/src/sim/sim_mmio.scala 55:19]
  wire  disk_disk_rdata_MPORT_7_en; // @[playground/src/sim/sim_mmio.scala 55:19]
  wire [25:0] disk_disk_rdata_MPORT_7_addr; // @[playground/src/sim/sim_mmio.scala 55:19]
  wire [7:0] disk_disk_rdata_MPORT_7_data; // @[playground/src/sim/sim_mmio.scala 55:19]
  wire [7:0] disk_MPORT_4_data; // @[playground/src/sim/sim_mmio.scala 55:19]
  wire [25:0] disk_MPORT_4_addr; // @[playground/src/sim/sim_mmio.scala 55:19]
  wire  disk_MPORT_4_mask; // @[playground/src/sim/sim_mmio.scala 55:19]
  wire  disk_MPORT_4_en; // @[playground/src/sim/sim_mmio.scala 55:19]
  wire [7:0] disk_MPORT_5_data; // @[playground/src/sim/sim_mmio.scala 55:19]
  wire [25:0] disk_MPORT_5_addr; // @[playground/src/sim/sim_mmio.scala 55:19]
  wire  disk_MPORT_5_mask; // @[playground/src/sim/sim_mmio.scala 55:19]
  wire  disk_MPORT_5_en; // @[playground/src/sim/sim_mmio.scala 55:19]
  wire [7:0] disk_MPORT_6_data; // @[playground/src/sim/sim_mmio.scala 55:19]
  wire [25:0] disk_MPORT_6_addr; // @[playground/src/sim/sim_mmio.scala 55:19]
  wire  disk_MPORT_6_mask; // @[playground/src/sim/sim_mmio.scala 55:19]
  wire  disk_MPORT_6_en; // @[playground/src/sim/sim_mmio.scala 55:19]
  wire [7:0] disk_MPORT_7_data; // @[playground/src/sim/sim_mmio.scala 55:19]
  wire [25:0] disk_MPORT_7_addr; // @[playground/src/sim/sim_mmio.scala 55:19]
  wire  disk_MPORT_7_mask; // @[playground/src/sim/sim_mmio.scala 55:19]
  wire  disk_MPORT_7_en; // @[playground/src/sim/sim_mmio.scala 55:19]
  wire [7:0] disk_MPORT_8_data; // @[playground/src/sim/sim_mmio.scala 55:19]
  wire [25:0] disk_MPORT_8_addr; // @[playground/src/sim/sim_mmio.scala 55:19]
  wire  disk_MPORT_8_mask; // @[playground/src/sim/sim_mmio.scala 55:19]
  wire  disk_MPORT_8_en; // @[playground/src/sim/sim_mmio.scala 55:19]
  wire [7:0] disk_MPORT_9_data; // @[playground/src/sim/sim_mmio.scala 55:19]
  wire [25:0] disk_MPORT_9_addr; // @[playground/src/sim/sim_mmio.scala 55:19]
  wire  disk_MPORT_9_mask; // @[playground/src/sim/sim_mmio.scala 55:19]
  wire  disk_MPORT_9_en; // @[playground/src/sim/sim_mmio.scala 55:19]
  wire [7:0] disk_MPORT_10_data; // @[playground/src/sim/sim_mmio.scala 55:19]
  wire [25:0] disk_MPORT_10_addr; // @[playground/src/sim/sim_mmio.scala 55:19]
  wire  disk_MPORT_10_mask; // @[playground/src/sim/sim_mmio.scala 55:19]
  wire  disk_MPORT_10_en; // @[playground/src/sim/sim_mmio.scala 55:19]
  wire [7:0] disk_MPORT_11_data; // @[playground/src/sim/sim_mmio.scala 55:19]
  wire [25:0] disk_MPORT_11_addr; // @[playground/src/sim/sim_mmio.scala 55:19]
  wire  disk_MPORT_11_mask; // @[playground/src/sim/sim_mmio.scala 55:19]
  wire  disk_MPORT_11_en; // @[playground/src/sim/sim_mmio.scala 55:19]
  reg /* sparse */ [7:0] flash [0:268435455]; // @[playground/src/sim/sim_mmio.scala 56:20]
  wire  flash_flash_rdata_MPORT_en; // @[playground/src/sim/sim_mmio.scala 56:20]
  wire [27:0] flash_flash_rdata_MPORT_addr; // @[playground/src/sim/sim_mmio.scala 56:20]
  wire [7:0] flash_flash_rdata_MPORT_data; // @[playground/src/sim/sim_mmio.scala 56:20]
  wire  flash_flash_rdata_MPORT_1_en; // @[playground/src/sim/sim_mmio.scala 56:20]
  wire [27:0] flash_flash_rdata_MPORT_1_addr; // @[playground/src/sim/sim_mmio.scala 56:20]
  wire [7:0] flash_flash_rdata_MPORT_1_data; // @[playground/src/sim/sim_mmio.scala 56:20]
  wire  flash_flash_rdata_MPORT_2_en; // @[playground/src/sim/sim_mmio.scala 56:20]
  wire [27:0] flash_flash_rdata_MPORT_2_addr; // @[playground/src/sim/sim_mmio.scala 56:20]
  wire [7:0] flash_flash_rdata_MPORT_2_data; // @[playground/src/sim/sim_mmio.scala 56:20]
  wire  flash_flash_rdata_MPORT_3_en; // @[playground/src/sim/sim_mmio.scala 56:20]
  wire [27:0] flash_flash_rdata_MPORT_3_addr; // @[playground/src/sim/sim_mmio.scala 56:20]
  wire [7:0] flash_flash_rdata_MPORT_3_data; // @[playground/src/sim/sim_mmio.scala 56:20]
  wire  flash_flash_rdata_MPORT_4_en; // @[playground/src/sim/sim_mmio.scala 56:20]
  wire [27:0] flash_flash_rdata_MPORT_4_addr; // @[playground/src/sim/sim_mmio.scala 56:20]
  wire [7:0] flash_flash_rdata_MPORT_4_data; // @[playground/src/sim/sim_mmio.scala 56:20]
  wire  flash_flash_rdata_MPORT_5_en; // @[playground/src/sim/sim_mmio.scala 56:20]
  wire [27:0] flash_flash_rdata_MPORT_5_addr; // @[playground/src/sim/sim_mmio.scala 56:20]
  wire [7:0] flash_flash_rdata_MPORT_5_data; // @[playground/src/sim/sim_mmio.scala 56:20]
  wire  flash_flash_rdata_MPORT_6_en; // @[playground/src/sim/sim_mmio.scala 56:20]
  wire [27:0] flash_flash_rdata_MPORT_6_addr; // @[playground/src/sim/sim_mmio.scala 56:20]
  wire [7:0] flash_flash_rdata_MPORT_6_data; // @[playground/src/sim/sim_mmio.scala 56:20]
  wire  flash_flash_rdata_MPORT_7_en; // @[playground/src/sim/sim_mmio.scala 56:20]
  wire [27:0] flash_flash_rdata_MPORT_7_addr; // @[playground/src/sim/sim_mmio.scala 56:20]
  wire [7:0] flash_flash_rdata_MPORT_7_data; // @[playground/src/sim/sim_mmio.scala 56:20]
  reg [7:0] uart_0; // @[playground/src/sim/sim_mmio.scala 50:23]
  reg [7:0] uart_1; // @[playground/src/sim/sim_mmio.scala 50:23]
  reg [7:0] uart_2; // @[playground/src/sim/sim_mmio.scala 50:23]
  reg [7:0] uart_3; // @[playground/src/sim/sim_mmio.scala 50:23]
  reg [7:0] uart_4; // @[playground/src/sim/sim_mmio.scala 50:23]
  reg [7:0] uart_5; // @[playground/src/sim/sim_mmio.scala 50:23]
  reg [7:0] uart_6; // @[playground/src/sim/sim_mmio.scala 50:23]
  reg [7:0] uart_7; // @[playground/src/sim/sim_mmio.scala 50:23]
  reg [63:0] mtime; // @[playground/src/sim/sim_mmio.scala 51:24]
  reg [63:0] mtimecmp; // @[playground/src/sim/sim_mmio.scala 52:27]
  reg  waready; // @[playground/src/sim/sim_mmio.scala 58:27]
  reg  wdready; // @[playground/src/sim/sim_mmio.scala 59:27]
  reg [31:0] waddr; // @[playground/src/sim/sim_mmio.scala 60:26]
  reg  raready; // @[playground/src/sim/sim_mmio.scala 64:26]
  reg  rdvalid; // @[playground/src/sim/sim_mmio.scala 65:26]
  reg [63:0] rdata; // @[playground/src/sim/sim_mmio.scala 67:26]
  reg [7:0] offset; // @[playground/src/sim/sim_mmio.scala 69:26]
  wire [63:0] _mtime_T_1 = mtime + 64'h14; // @[playground/src/sim/sim_mmio.scala 76:24]
  reg [2:0] state; // @[playground/src/sim/sim_mmio.scala 78:24]
  wire  islast = offset == 8'h0; // @[playground/src/sim/sim_mmio.scala 79:27]
  wire [7:0] _inputwd_T_3 = io_mmioAxi_wd_bits_strb[7] ? io_mmioAxi_wd_bits_data[63:56] : 8'h0; // @[playground/src/sim/sim_mmio.scala 81:55]
  wire [7:0] _inputwd_T_7 = io_mmioAxi_wd_bits_strb[6] ? io_mmioAxi_wd_bits_data[55:48] : 8'h0; // @[playground/src/sim/sim_mmio.scala 81:55]
  wire [7:0] _inputwd_T_11 = io_mmioAxi_wd_bits_strb[5] ? io_mmioAxi_wd_bits_data[47:40] : 8'h0; // @[playground/src/sim/sim_mmio.scala 81:55]
  wire [7:0] _inputwd_T_15 = io_mmioAxi_wd_bits_strb[4] ? io_mmioAxi_wd_bits_data[39:32] : 8'h0; // @[playground/src/sim/sim_mmio.scala 81:55]
  wire [7:0] _inputwd_T_19 = io_mmioAxi_wd_bits_strb[3] ? io_mmioAxi_wd_bits_data[31:24] : 8'h0; // @[playground/src/sim/sim_mmio.scala 81:55]
  wire [7:0] _inputwd_T_23 = io_mmioAxi_wd_bits_strb[2] ? io_mmioAxi_wd_bits_data[23:16] : 8'h0; // @[playground/src/sim/sim_mmio.scala 81:55]
  wire [7:0] _inputwd_T_27 = io_mmioAxi_wd_bits_strb[1] ? io_mmioAxi_wd_bits_data[15:8] : 8'h0; // @[playground/src/sim/sim_mmio.scala 81:55]
  wire [7:0] _inputwd_T_31 = io_mmioAxi_wd_bits_strb[0] ? io_mmioAxi_wd_bits_data[7:0] : 8'h0; // @[playground/src/sim/sim_mmio.scala 81:55]
  wire [63:0] inputwd = {_inputwd_T_3,_inputwd_T_7,_inputwd_T_11,_inputwd_T_15,_inputwd_T_19,_inputwd_T_23,_inputwd_T_27
    ,_inputwd_T_31}; // @[playground/src/sim/sim_mmio.scala 81:22]
  wire [31:0] _disk_rdata_T_1 = io_mmioAxi_ra_bits_addr + 32'h7; // @[playground/src/sim/sim_mmio.scala 82:87]
  wire [31:0] _disk_rdata_T_2 = _disk_rdata_T_1 & 32'h3ffffff; // @[playground/src/sim/sim_mmio.scala 82:93]
  wire [31:0] _disk_rdata_T_5 = io_mmioAxi_ra_bits_addr + 32'h6; // @[playground/src/sim/sim_mmio.scala 82:87]
  wire [31:0] _disk_rdata_T_6 = _disk_rdata_T_5 & 32'h3ffffff; // @[playground/src/sim/sim_mmio.scala 82:93]
  wire [31:0] _disk_rdata_T_9 = io_mmioAxi_ra_bits_addr + 32'h5; // @[playground/src/sim/sim_mmio.scala 82:87]
  wire [31:0] _disk_rdata_T_10 = _disk_rdata_T_9 & 32'h3ffffff; // @[playground/src/sim/sim_mmio.scala 82:93]
  wire [31:0] _disk_rdata_T_13 = io_mmioAxi_ra_bits_addr + 32'h4; // @[playground/src/sim/sim_mmio.scala 82:87]
  wire [31:0] _disk_rdata_T_14 = _disk_rdata_T_13 & 32'h3ffffff; // @[playground/src/sim/sim_mmio.scala 82:93]
  wire [31:0] _disk_rdata_T_17 = io_mmioAxi_ra_bits_addr + 32'h3; // @[playground/src/sim/sim_mmio.scala 82:87]
  wire [31:0] _disk_rdata_T_18 = _disk_rdata_T_17 & 32'h3ffffff; // @[playground/src/sim/sim_mmio.scala 82:93]
  wire [31:0] _disk_rdata_T_21 = io_mmioAxi_ra_bits_addr + 32'h2; // @[playground/src/sim/sim_mmio.scala 82:87]
  wire [31:0] _disk_rdata_T_22 = _disk_rdata_T_21 & 32'h3ffffff; // @[playground/src/sim/sim_mmio.scala 82:93]
  wire [31:0] _disk_rdata_T_25 = io_mmioAxi_ra_bits_addr + 32'h1; // @[playground/src/sim/sim_mmio.scala 82:87]
  wire [31:0] _disk_rdata_T_26 = _disk_rdata_T_25 & 32'h3ffffff; // @[playground/src/sim/sim_mmio.scala 82:93]
  wire [32:0] _disk_rdata_T_28 = {{1'd0}, io_mmioAxi_ra_bits_addr}; // @[playground/src/sim/sim_mmio.scala 82:87]
  wire [31:0] _disk_rdata_T_30 = _disk_rdata_T_28[31:0] & 32'h3ffffff; // @[playground/src/sim/sim_mmio.scala 82:93]
  wire [63:0] disk_rdata = {disk_disk_rdata_MPORT_data,disk_disk_rdata_MPORT_1_data,disk_disk_rdata_MPORT_2_data,
    disk_disk_rdata_MPORT_3_data,disk_disk_rdata_MPORT_4_data,disk_disk_rdata_MPORT_5_data,disk_disk_rdata_MPORT_6_data,
    disk_disk_rdata_MPORT_7_data}; // @[playground/src/sim/sim_mmio.scala 82:27]
  wire [31:0] _flash_rdata_T = io_mmioAxi_ra_bits_addr & 32'hffffff8; // @[playground/src/sim/sim_mmio.scala 83:89]
  wire [31:0] _flash_rdata_T_2 = _flash_rdata_T + 32'h7; // @[playground/src/sim/sim_mmio.scala 83:104]
  wire [31:0] _flash_rdata_T_6 = _flash_rdata_T + 32'h6; // @[playground/src/sim/sim_mmio.scala 83:104]
  wire [31:0] _flash_rdata_T_10 = _flash_rdata_T + 32'h5; // @[playground/src/sim/sim_mmio.scala 83:104]
  wire [31:0] _flash_rdata_T_14 = _flash_rdata_T + 32'h4; // @[playground/src/sim/sim_mmio.scala 83:104]
  wire [31:0] _flash_rdata_T_18 = _flash_rdata_T + 32'h3; // @[playground/src/sim/sim_mmio.scala 83:104]
  wire [31:0] _flash_rdata_T_22 = _flash_rdata_T + 32'h2; // @[playground/src/sim/sim_mmio.scala 83:104]
  wire [31:0] _flash_rdata_T_26 = _flash_rdata_T + 32'h1; // @[playground/src/sim/sim_mmio.scala 83:104]
  wire [32:0] _flash_rdata_T_29 = {{1'd0}, _flash_rdata_T}; // @[playground/src/sim/sim_mmio.scala 83:104]
  wire [63:0] flash_rdata = {flash_flash_rdata_MPORT_data,flash_flash_rdata_MPORT_1_data,flash_flash_rdata_MPORT_2_data,
    flash_flash_rdata_MPORT_3_data,flash_flash_rdata_MPORT_4_data,flash_flash_rdata_MPORT_5_data,
    flash_flash_rdata_MPORT_6_data,flash_flash_rdata_MPORT_7_data}; // @[playground/src/sim/sim_mmio.scala 83:28]
  wire  _T_1 = 3'h0 == state; // @[playground/src/sim/sim_mmio.scala 85:18]
  wire  _T_3 = io_mmioAxi_ra_valid & raready; // @[playground/src/sim/sim_mmio.scala 96:38]
  wire  _T_8 = io_mmioAxi_ra_bits_addr >= 32'h10000000 & io_mmioAxi_ra_bits_addr <= 32'h10000007; // @[playground/src/sim/sim_mmio.scala 100:64]
  wire [31:0] _rdata_T_1 = io_mmioAxi_ra_bits_addr - 32'h10000000; // @[playground/src/sim/sim_mmio.scala 101:61]
  wire [6:0] _rdata_T_4 = io_mmioAxi_ra_bits_addr[2:0] * 4'h8; // @[playground/src/sim/sim_mmio.scala 101:112]
  wire [7:0] _GEN_6 = 3'h1 == _rdata_T_1[2:0] ? uart_1 : uart_0; // @[playground/src/sim/sim_mmio.scala 101:{79,79}]
  wire [7:0] _GEN_7 = 3'h2 == _rdata_T_1[2:0] ? uart_2 : _GEN_6; // @[playground/src/sim/sim_mmio.scala 101:{79,79}]
  wire [7:0] _GEN_8 = 3'h3 == _rdata_T_1[2:0] ? uart_3 : _GEN_7; // @[playground/src/sim/sim_mmio.scala 101:{79,79}]
  wire [7:0] _GEN_9 = 3'h4 == _rdata_T_1[2:0] ? uart_4 : _GEN_8; // @[playground/src/sim/sim_mmio.scala 101:{79,79}]
  wire [7:0] _GEN_10 = 3'h5 == _rdata_T_1[2:0] ? uart_5 : _GEN_9; // @[playground/src/sim/sim_mmio.scala 101:{79,79}]
  wire [7:0] _GEN_11 = 3'h6 == _rdata_T_1[2:0] ? uart_6 : _GEN_10; // @[playground/src/sim/sim_mmio.scala 101:{79,79}]
  wire [7:0] _GEN_12 = 3'h7 == _rdata_T_1[2:0] ? uart_7 : _GEN_11; // @[playground/src/sim/sim_mmio.scala 101:{79,79}]
  wire [134:0] _GEN_391 = {{127'd0}, _GEN_12}; // @[playground/src/sim/sim_mmio.scala 101:79]
  wire [134:0] _rdata_T_5 = _GEN_391 << _rdata_T_4; // @[playground/src/sim/sim_mmio.scala 101:79]
  wire  _T_9 = io_mmioAxi_ra_bits_addr == 32'h200bff8; // @[playground/src/sim/sim_mmio.scala 102:52]
  wire  _T_10 = io_mmioAxi_ra_bits_addr == 32'h2004000; // @[playground/src/sim/sim_mmio.scala 104:52]
  wire  _T_11 = io_mmioAxi_ra_bits_addr == 32'ha1000100; // @[playground/src/sim/sim_mmio.scala 106:52]
  wire  _T_12 = io_mmioAxi_ra_bits_addr == 32'ha1000048; // @[playground/src/sim/sim_mmio.scala 108:52]
  wire [63:0] _rdata_T_6 = mtime % 64'hf4240; // @[playground/src/sim/sim_mmio.scala 109:39]
  wire  _T_15 = io_mmioAxi_ra_bits_addr == 32'ha100004c; // @[playground/src/sim/sim_mmio.scala 110:52]
  wire [63:0] _rdata_T_8 = mtime / 64'hf4240; // @[playground/src/sim/sim_mmio.scala 111:43]
  wire [63:0] _rdata_T_11 = {_rdata_T_8[31:0],32'h0}; // @[playground/src/sim/sim_mmio.scala 111:35]
  wire  _T_16 = io_mmioAxi_ra_bits_addr == 32'ha1000060; // @[playground/src/sim/sim_mmio.scala 112:52]
  wire  _T_17 = io_mmioAxi_ra_bits_addr == 32'h2000000; // @[playground/src/sim/sim_mmio.scala 115:52]
  wire  _T_22 = io_mmioAxi_ra_bits_addr >= 32'hc000000 & io_mmioAxi_ra_bits_addr < 32'hc003000; // @[playground/src/sim/sim_mmio.scala 117:65]
  wire  _T_27 = io_mmioAxi_ra_bits_addr >= 32'h43000000 & io_mmioAxi_ra_bits_addr < 32'h43000080; // @[playground/src/sim/sim_mmio.scala 119:72]
  wire  _T_32 = io_mmioAxi_ra_bits_addr >= 32'h40000000 & io_mmioAxi_ra_bits_addr < 32'h44000000; // @[playground/src/sim/sim_mmio.scala 123:70]
  wire  _T_37 = io_mmioAxi_ra_bits_addr >= 32'h30000000 & io_mmioAxi_ra_bits_addr < 32'h40000000; // @[playground/src/sim/sim_mmio.scala 125:71]
  wire  _T_39 = ~reset; // @[playground/src/sim/sim_mmio.scala 129:27]
  wire [63:0] _GEN_13 = io_mmioAxi_ra_bits_addr >= 32'h30000000 & io_mmioAxi_ra_bits_addr < 32'h40000000 ? flash_rdata
     : 64'h0; // @[playground/src/sim/sim_mmio.scala 125:134 126:27 128:29]
  wire [63:0] _GEN_14 = io_mmioAxi_ra_bits_addr >= 32'h40000000 & io_mmioAxi_ra_bits_addr < 32'h44000000 ? disk_rdata :
    _GEN_13; // @[playground/src/sim/sim_mmio.scala 123:131 124:27]
  wire [6:0] _GEN_15 = io_mmioAxi_ra_bits_addr >= 32'h43000000 & io_mmioAxi_ra_bits_addr < 32'h43000080 ?
    io_mmioAxi_ra_bits_addr[6:0] : 7'h0; // @[playground/src/sim/sim_mmio.scala 119:129 120:37 47:20]
  wire [2:0] _GEN_17 = io_mmioAxi_ra_bits_addr >= 32'h43000000 & io_mmioAxi_ra_bits_addr < 32'h43000080 ? 3'h4 : 3'h3; // @[playground/src/sim/sim_mmio.scala 119:129 122:37 99:25]
  wire [63:0] _GEN_18 = io_mmioAxi_ra_bits_addr >= 32'h43000000 & io_mmioAxi_ra_bits_addr < 32'h43000080 ? rdata :
    _GEN_14; // @[playground/src/sim/sim_mmio.scala 119:129 67:26]
  wire [6:0] _GEN_19 = io_mmioAxi_ra_bits_addr >= 32'hc000000 & io_mmioAxi_ra_bits_addr < 32'hc003000 ? 7'h0 : _GEN_15; // @[playground/src/sim/sim_mmio.scala 117:117 47:20]
  wire  _GEN_20 = io_mmioAxi_ra_bits_addr >= 32'hc000000 & io_mmioAxi_ra_bits_addr < 32'hc003000 ? 1'h0 : _T_27; // @[playground/src/sim/sim_mmio.scala 117:117 47:68]
  wire [2:0] _GEN_21 = io_mmioAxi_ra_bits_addr >= 32'hc000000 & io_mmioAxi_ra_bits_addr < 32'hc003000 ? 3'h3 : _GEN_17; // @[playground/src/sim/sim_mmio.scala 117:117 99:25]
  wire [63:0] _GEN_22 = io_mmioAxi_ra_bits_addr >= 32'hc000000 & io_mmioAxi_ra_bits_addr < 32'hc003000 ? rdata : _GEN_18
    ; // @[playground/src/sim/sim_mmio.scala 117:117 67:26]
  wire [63:0] _GEN_23 = io_mmioAxi_ra_bits_addr == 32'h2000000 ? 64'h0 : _GEN_22; // @[playground/src/sim/sim_mmio.scala 115:67 116:27]
  wire [6:0] _GEN_24 = io_mmioAxi_ra_bits_addr == 32'h2000000 ? 7'h0 : _GEN_19; // @[playground/src/sim/sim_mmio.scala 115:67 47:20]
  wire  _GEN_25 = io_mmioAxi_ra_bits_addr == 32'h2000000 ? 1'h0 : _GEN_20; // @[playground/src/sim/sim_mmio.scala 115:67 47:68]
  wire [2:0] _GEN_26 = io_mmioAxi_ra_bits_addr == 32'h2000000 ? 3'h3 : _GEN_21; // @[playground/src/sim/sim_mmio.scala 115:67 99:25]
  wire [63:0] _GEN_27 = io_mmioAxi_ra_bits_addr == 32'ha1000060 ? 64'h0 : _GEN_23; // @[playground/src/sim/sim_mmio.scala 112:70 114:27]
  wire [6:0] _GEN_28 = io_mmioAxi_ra_bits_addr == 32'ha1000060 ? 7'h0 : _GEN_24; // @[playground/src/sim/sim_mmio.scala 112:70 47:20]
  wire  _GEN_29 = io_mmioAxi_ra_bits_addr == 32'ha1000060 ? 1'h0 : _GEN_25; // @[playground/src/sim/sim_mmio.scala 112:70 47:68]
  wire [2:0] _GEN_30 = io_mmioAxi_ra_bits_addr == 32'ha1000060 ? 3'h3 : _GEN_26; // @[playground/src/sim/sim_mmio.scala 112:70 99:25]
  wire [63:0] _GEN_31 = io_mmioAxi_ra_bits_addr == 32'ha100004c ? _rdata_T_11 : _GEN_27; // @[playground/src/sim/sim_mmio.scala 110:76 111:29]
  wire [6:0] _GEN_32 = io_mmioAxi_ra_bits_addr == 32'ha100004c ? 7'h0 : _GEN_28; // @[playground/src/sim/sim_mmio.scala 110:76 47:20]
  wire  _GEN_33 = io_mmioAxi_ra_bits_addr == 32'ha100004c ? 1'h0 : _GEN_29; // @[playground/src/sim/sim_mmio.scala 110:76 47:68]
  wire [2:0] _GEN_34 = io_mmioAxi_ra_bits_addr == 32'ha100004c ? 3'h3 : _GEN_30; // @[playground/src/sim/sim_mmio.scala 110:76 99:25]
  wire [63:0] _GEN_35 = io_mmioAxi_ra_bits_addr == 32'ha1000048 ? {{32'd0}, _rdata_T_6[31:0]} : _GEN_31; // @[playground/src/sim/sim_mmio.scala 108:70 109:29]
  wire [6:0] _GEN_36 = io_mmioAxi_ra_bits_addr == 32'ha1000048 ? 7'h0 : _GEN_32; // @[playground/src/sim/sim_mmio.scala 108:70 47:20]
  wire  _GEN_37 = io_mmioAxi_ra_bits_addr == 32'ha1000048 ? 1'h0 : _GEN_33; // @[playground/src/sim/sim_mmio.scala 108:70 47:68]
  wire [2:0] _GEN_38 = io_mmioAxi_ra_bits_addr == 32'ha1000048 ? 3'h3 : _GEN_34; // @[playground/src/sim/sim_mmio.scala 108:70 99:25]
  wire [63:0] _GEN_39 = io_mmioAxi_ra_bits_addr == 32'ha1000100 ? 64'h190012c : _GEN_35; // @[playground/src/sim/sim_mmio.scala 106:85 107:29]
  wire [6:0] _GEN_40 = io_mmioAxi_ra_bits_addr == 32'ha1000100 ? 7'h0 : _GEN_36; // @[playground/src/sim/sim_mmio.scala 106:85 47:20]
  wire  _GEN_41 = io_mmioAxi_ra_bits_addr == 32'ha1000100 ? 1'h0 : _GEN_37; // @[playground/src/sim/sim_mmio.scala 106:85 47:68]
  wire [2:0] _GEN_42 = io_mmioAxi_ra_bits_addr == 32'ha1000100 ? 3'h3 : _GEN_38; // @[playground/src/sim/sim_mmio.scala 106:85 99:25]
  wire [63:0] _GEN_43 = io_mmioAxi_ra_bits_addr == 32'h2004000 ? mtimecmp : _GEN_39; // @[playground/src/sim/sim_mmio.scala 104:76 105:29]
  wire [6:0] _GEN_44 = io_mmioAxi_ra_bits_addr == 32'h2004000 ? 7'h0 : _GEN_40; // @[playground/src/sim/sim_mmio.scala 104:76 47:20]
  wire  _GEN_45 = io_mmioAxi_ra_bits_addr == 32'h2004000 ? 1'h0 : _GEN_41; // @[playground/src/sim/sim_mmio.scala 104:76 47:68]
  wire [2:0] _GEN_46 = io_mmioAxi_ra_bits_addr == 32'h2004000 ? 3'h3 : _GEN_42; // @[playground/src/sim/sim_mmio.scala 104:76 99:25]
  wire [63:0] _GEN_47 = io_mmioAxi_ra_bits_addr == 32'h200bff8 ? mtime : _GEN_43; // @[playground/src/sim/sim_mmio.scala 102:73 103:29]
  wire [6:0] _GEN_48 = io_mmioAxi_ra_bits_addr == 32'h200bff8 ? 7'h0 : _GEN_44; // @[playground/src/sim/sim_mmio.scala 102:73 47:20]
  wire  _GEN_49 = io_mmioAxi_ra_bits_addr == 32'h200bff8 ? 1'h0 : _GEN_45; // @[playground/src/sim/sim_mmio.scala 102:73 47:68]
  wire [2:0] _GEN_50 = io_mmioAxi_ra_bits_addr == 32'h200bff8 ? 3'h3 : _GEN_46; // @[playground/src/sim/sim_mmio.scala 102:73 99:25]
  wire [134:0] _GEN_51 = io_mmioAxi_ra_bits_addr >= 32'h10000000 & io_mmioAxi_ra_bits_addr <= 32'h10000007 ? _rdata_T_5
     : {{71'd0}, _GEN_47}; // @[playground/src/sim/sim_mmio.scala 100:115 101:29]
  wire [6:0] _GEN_52 = io_mmioAxi_ra_bits_addr >= 32'h10000000 & io_mmioAxi_ra_bits_addr <= 32'h10000007 ? 7'h0 :
    _GEN_48; // @[playground/src/sim/sim_mmio.scala 100:115 47:20]
  wire  _GEN_53 = io_mmioAxi_ra_bits_addr >= 32'h10000000 & io_mmioAxi_ra_bits_addr <= 32'h10000007 ? 1'h0 : _GEN_49; // @[playground/src/sim/sim_mmio.scala 100:115 47:68]
  wire [134:0] _GEN_58 = io_mmioAxi_ra_valid & raready ? _GEN_51 : {{71'd0}, rdata}; // @[playground/src/sim/sim_mmio.scala 67:26 96:49]
  wire [6:0] _GEN_59 = io_mmioAxi_ra_valid & raready ? _GEN_52 : 7'h0; // @[playground/src/sim/sim_mmio.scala 47:20 96:49]
  wire  _GEN_60 = io_mmioAxi_ra_valid & raready & _GEN_53; // @[playground/src/sim/sim_mmio.scala 96:49 47:68]
  wire  _T_40 = 3'h1 == state; // @[playground/src/sim/sim_mmio.scala 85:18]
  wire  _T_45 = waddr >= 32'h10000000 & waddr <= 32'h10000007; // @[playground/src/sim/sim_mmio.scala 139:46]
  wire [2:0] offset_1 = waddr[2:0]; // @[playground/src/sim/sim_mmio.scala 140:39]
  wire [31:0] _T_47 = waddr - 32'h10000000; // @[playground/src/sim/sim_mmio.scala 141:32]
  wire [6:0] _uart_T = offset_1 * 4'h8; // @[playground/src/sim/sim_mmio.scala 141:72]
  wire [63:0] _uart_T_1 = inputwd >> _uart_T; // @[playground/src/sim/sim_mmio.scala 141:62]
  wire [7:0] _GEN_61 = 3'h0 == _T_47[2:0] ? _uart_T_1[7:0] : uart_0; // @[playground/src/sim/sim_mmio.scala 141:{50,50} 50:23]
  wire [7:0] _GEN_62 = 3'h1 == _T_47[2:0] ? _uart_T_1[7:0] : uart_1; // @[playground/src/sim/sim_mmio.scala 141:{50,50} 50:23]
  wire [7:0] _GEN_63 = 3'h2 == _T_47[2:0] ? _uart_T_1[7:0] : uart_2; // @[playground/src/sim/sim_mmio.scala 141:{50,50} 50:23]
  wire [7:0] _GEN_64 = 3'h3 == _T_47[2:0] ? _uart_T_1[7:0] : uart_3; // @[playground/src/sim/sim_mmio.scala 141:{50,50} 50:23]
  wire [7:0] _GEN_65 = 3'h4 == _T_47[2:0] ? _uart_T_1[7:0] : uart_4; // @[playground/src/sim/sim_mmio.scala 141:{50,50} 50:23]
  wire [7:0] _GEN_66 = 3'h5 == _T_47[2:0] ? _uart_T_1[7:0] : 8'h20; // @[playground/src/sim/sim_mmio.scala 141:{50,50} 84:13]
  wire [7:0] _GEN_67 = 3'h6 == _T_47[2:0] ? _uart_T_1[7:0] : uart_6; // @[playground/src/sim/sim_mmio.scala 141:{50,50} 50:23]
  wire [7:0] _GEN_68 = 3'h7 == _T_47[2:0] ? _uart_T_1[7:0] : uart_7; // @[playground/src/sim/sim_mmio.scala 141:{50,50} 50:23]
  wire [31:0] _T_49 = waddr & 32'h7; // @[playground/src/sim/sim_mmio.scala 142:33]
  wire  _T_50 = _T_49 == 32'h0; // @[playground/src/sim/sim_mmio.scala 142:42]
  wire  _T_54 = waddr == 32'h2004000; // @[playground/src/sim/sim_mmio.scala 145:34]
  wire  _T_55 = waddr == 32'ha10003f8; // @[playground/src/sim/sim_mmio.scala 148:32]
  wire  _T_63 = waddr >= 32'ha0000000 & waddr <= 32'ha0075300; // @[playground/src/sim/sim_mmio.scala 150:55]
  wire  _T_100 = waddr == 32'ha1000100; // @[playground/src/sim/sim_mmio.scala 154:38]
  wire  _T_101 = waddr == 32'ha1000104; // @[playground/src/sim/sim_mmio.scala 156:38]
  wire  _T_102 = waddr >= 32'hc000000; // @[playground/src/sim/sim_mmio.scala 158:38]
  wire  _T_104 = waddr >= 32'hc000000 & waddr <= 32'hc202000; // @[playground/src/sim/sim_mmio.scala 158:55]
  wire  _T_105 = waddr == 32'h2000000; // @[playground/src/sim/sim_mmio.scala 160:38]
  wire  _T_110 = _T_102 & waddr < 32'hc003000; // @[playground/src/sim/sim_mmio.scala 162:51]
  wire  _T_115 = waddr >= 32'h43000000 & waddr < 32'h43000080; // @[playground/src/sim/sim_mmio.scala 164:58]
  wire [5:0] _sdcard_io_wdata_T_1 = {offset_1,3'h0}; // @[playground/src/sim/sim_mmio.scala 166:58]
  wire [63:0] _sdcard_io_wdata_T_2 = inputwd >> _sdcard_io_wdata_T_1; // @[playground/src/sim/sim_mmio.scala 166:52]
  wire [32:0] _T_121 = {{1'd0}, waddr}; // @[playground/src/sim/sim_mmio.scala 170:40]
  wire [31:0] _T_126 = waddr + 32'h1; // @[playground/src/sim/sim_mmio.scala 170:40]
  wire [31:0] _T_130 = waddr + 32'h2; // @[playground/src/sim/sim_mmio.scala 170:40]
  wire [31:0] _T_134 = waddr + 32'h3; // @[playground/src/sim/sim_mmio.scala 170:40]
  wire [31:0] _T_138 = waddr + 32'h4; // @[playground/src/sim/sim_mmio.scala 170:40]
  wire [31:0] _T_142 = waddr + 32'h5; // @[playground/src/sim/sim_mmio.scala 170:40]
  wire [31:0] _T_146 = waddr + 32'h6; // @[playground/src/sim/sim_mmio.scala 170:40]
  wire [31:0] _T_150 = waddr + 32'h7; // @[playground/src/sim/sim_mmio.scala 170:40]
  wire [6:0] _GEN_88 = waddr >= 32'h43000000 & waddr < 32'h43000080 ? waddr[6:0] : 7'h0; // @[playground/src/sim/sim_mmio.scala 164:95 165:41 47:20]
  wire [63:0] _GEN_89 = waddr >= 32'h43000000 & waddr < 32'h43000080 ? _sdcard_io_wdata_T_2 : 64'h0; // @[playground/src/sim/sim_mmio.scala 164:95 166:41 47:96]
  wire  _GEN_93 = waddr >= 32'h43000000 & waddr < 32'h43000080 ? 1'h0 : _T_32; // @[playground/src/sim/sim_mmio.scala 164:95 55:19]
  wire [6:0] _GEN_110 = _T_102 & waddr < 32'hc003000 ? 7'h0 : _GEN_88; // @[playground/src/sim/sim_mmio.scala 162:85 47:20]
  wire [63:0] _GEN_111 = _T_102 & waddr < 32'hc003000 ? 64'h0 : _GEN_89; // @[playground/src/sim/sim_mmio.scala 162:85 47:96]
  wire  _GEN_112 = _T_102 & waddr < 32'hc003000 ? 1'h0 : _T_115; // @[playground/src/sim/sim_mmio.scala 162:85 47:42]
  wire  _GEN_115 = _T_102 & waddr < 32'hc003000 ? 1'h0 : _GEN_93; // @[playground/src/sim/sim_mmio.scala 162:85 55:19]
  wire [6:0] _GEN_132 = waddr == 32'h2000000 ? 7'h0 : _GEN_110; // @[playground/src/sim/sim_mmio.scala 160:53 47:20]
  wire [63:0] _GEN_133 = waddr == 32'h2000000 ? 64'h0 : _GEN_111; // @[playground/src/sim/sim_mmio.scala 160:53 47:96]
  wire  _GEN_134 = waddr == 32'h2000000 ? 1'h0 : _GEN_112; // @[playground/src/sim/sim_mmio.scala 160:53 47:42]
  wire  _GEN_137 = waddr == 32'h2000000 ? 1'h0 : _GEN_115; // @[playground/src/sim/sim_mmio.scala 160:53 55:19]
  wire [6:0] _GEN_154 = waddr >= 32'hc000000 & waddr <= 32'hc202000 ? 7'h0 : _GEN_132; // @[playground/src/sim/sim_mmio.scala 158:80 47:20]
  wire [63:0] _GEN_155 = waddr >= 32'hc000000 & waddr <= 32'hc202000 ? 64'h0 : _GEN_133; // @[playground/src/sim/sim_mmio.scala 158:80 47:96]
  wire  _GEN_156 = waddr >= 32'hc000000 & waddr <= 32'hc202000 ? 1'h0 : _GEN_134; // @[playground/src/sim/sim_mmio.scala 158:80 47:42]
  wire  _GEN_159 = waddr >= 32'hc000000 & waddr <= 32'hc202000 ? 1'h0 : _GEN_137; // @[playground/src/sim/sim_mmio.scala 158:80 55:19]
  wire [6:0] _GEN_177 = waddr == 32'ha1000104 ? 7'h0 : _GEN_154; // @[playground/src/sim/sim_mmio.scala 156:56 47:20]
  wire [63:0] _GEN_178 = waddr == 32'ha1000104 ? 64'h0 : _GEN_155; // @[playground/src/sim/sim_mmio.scala 156:56 47:96]
  wire  _GEN_179 = waddr == 32'ha1000104 ? 1'h0 : _GEN_156; // @[playground/src/sim/sim_mmio.scala 156:56 47:42]
  wire  _GEN_182 = waddr == 32'ha1000104 ? 1'h0 : _GEN_159; // @[playground/src/sim/sim_mmio.scala 156:56 55:19]
  wire [6:0] _GEN_201 = waddr == 32'ha1000100 ? 7'h0 : _GEN_177; // @[playground/src/sim/sim_mmio.scala 154:56 47:20]
  wire [63:0] _GEN_202 = waddr == 32'ha1000100 ? 64'h0 : _GEN_178; // @[playground/src/sim/sim_mmio.scala 154:56 47:96]
  wire  _GEN_203 = waddr == 32'ha1000100 ? 1'h0 : _GEN_179; // @[playground/src/sim/sim_mmio.scala 154:56 47:42]
  wire  _GEN_206 = waddr == 32'ha1000100 ? 1'h0 : _GEN_182; // @[playground/src/sim/sim_mmio.scala 154:56 55:19]
  wire [6:0] _GEN_236 = waddr >= 32'ha0000000 & waddr <= 32'ha0075300 ? 7'h0 : _GEN_201; // @[playground/src/sim/sim_mmio.scala 150:92 47:20]
  wire [63:0] _GEN_237 = waddr >= 32'ha0000000 & waddr <= 32'ha0075300 ? 64'h0 : _GEN_202; // @[playground/src/sim/sim_mmio.scala 150:92 47:96]
  wire  _GEN_238 = waddr >= 32'ha0000000 & waddr <= 32'ha0075300 ? 1'h0 : _GEN_203; // @[playground/src/sim/sim_mmio.scala 150:92 47:42]
  wire  _GEN_241 = waddr >= 32'ha0000000 & waddr <= 32'ha0075300 ? 1'h0 : _GEN_206; // @[playground/src/sim/sim_mmio.scala 150:92 55:19]
  wire [6:0] _GEN_271 = waddr == 32'ha10003f8 ? 7'h0 : _GEN_236; // @[playground/src/sim/sim_mmio.scala 148:50 47:20]
  wire [63:0] _GEN_272 = waddr == 32'ha10003f8 ? 64'h0 : _GEN_237; // @[playground/src/sim/sim_mmio.scala 148:50 47:96]
  wire  _GEN_273 = waddr == 32'ha10003f8 ? 1'h0 : _GEN_238; // @[playground/src/sim/sim_mmio.scala 148:50 47:42]
  wire  _GEN_276 = waddr == 32'ha10003f8 ? 1'h0 : _GEN_241; // @[playground/src/sim/sim_mmio.scala 148:50 55:19]
  wire [63:0] _GEN_293 = waddr == 32'h2004000 ? inputwd : mtimecmp; // @[playground/src/sim/sim_mmio.scala 145:58 146:30 52:27]
  wire [6:0] _GEN_307 = waddr == 32'h2004000 ? 7'h0 : _GEN_271; // @[playground/src/sim/sim_mmio.scala 145:58 47:20]
  wire [63:0] _GEN_308 = waddr == 32'h2004000 ? 64'h0 : _GEN_272; // @[playground/src/sim/sim_mmio.scala 145:58 47:96]
  wire  _GEN_309 = waddr == 32'h2004000 ? 1'h0 : _GEN_273; // @[playground/src/sim/sim_mmio.scala 145:58 47:42]
  wire  _GEN_312 = waddr == 32'h2004000 ? 1'h0 : _GEN_276; // @[playground/src/sim/sim_mmio.scala 145:58 55:19]
  wire [7:0] _GEN_329 = waddr >= 32'h10000000 & waddr <= 32'h10000007 ? _GEN_61 : uart_0; // @[playground/src/sim/sim_mmio.scala 139:79 50:23]
  wire [7:0] _GEN_330 = waddr >= 32'h10000000 & waddr <= 32'h10000007 ? _GEN_62 : uart_1; // @[playground/src/sim/sim_mmio.scala 139:79 50:23]
  wire [7:0] _GEN_331 = waddr >= 32'h10000000 & waddr <= 32'h10000007 ? _GEN_63 : uart_2; // @[playground/src/sim/sim_mmio.scala 139:79 50:23]
  wire [7:0] _GEN_332 = waddr >= 32'h10000000 & waddr <= 32'h10000007 ? _GEN_64 : uart_3; // @[playground/src/sim/sim_mmio.scala 139:79 50:23]
  wire [7:0] _GEN_333 = waddr >= 32'h10000000 & waddr <= 32'h10000007 ? _GEN_65 : uart_4; // @[playground/src/sim/sim_mmio.scala 139:79 50:23]
  wire [7:0] _GEN_334 = waddr >= 32'h10000000 & waddr <= 32'h10000007 ? _GEN_66 : 8'h20; // @[playground/src/sim/sim_mmio.scala 139:79 84:13]
  wire [7:0] _GEN_335 = waddr >= 32'h10000000 & waddr <= 32'h10000007 ? _GEN_67 : uart_6; // @[playground/src/sim/sim_mmio.scala 139:79 50:23]
  wire [7:0] _GEN_336 = waddr >= 32'h10000000 & waddr <= 32'h10000007 ? _GEN_68 : uart_7; // @[playground/src/sim/sim_mmio.scala 139:79 50:23]
  wire [63:0] _GEN_337 = waddr >= 32'h10000000 & waddr <= 32'h10000007 ? mtimecmp : _GEN_293; // @[playground/src/sim/sim_mmio.scala 139:79 52:27]
  wire [6:0] _GEN_351 = waddr >= 32'h10000000 & waddr <= 32'h10000007 ? 7'h0 : _GEN_307; // @[playground/src/sim/sim_mmio.scala 139:79 47:20]
  wire [63:0] _GEN_352 = waddr >= 32'h10000000 & waddr <= 32'h10000007 ? 64'h0 : _GEN_308; // @[playground/src/sim/sim_mmio.scala 139:79 47:96]
  wire  _GEN_353 = waddr >= 32'h10000000 & waddr <= 32'h10000007 ? 1'h0 : _GEN_309; // @[playground/src/sim/sim_mmio.scala 139:79 47:42]
  wire  _GEN_356 = waddr >= 32'h10000000 & waddr <= 32'h10000007 ? 1'h0 : _GEN_312; // @[playground/src/sim/sim_mmio.scala 139:79 55:19]
  wire [2:0] _GEN_373 = io_mmioAxi_wd_bits_last ? 3'h2 : state; // @[playground/src/sim/sim_mmio.scala 176:46 177:29 78:24]
  wire  _GEN_374 = io_mmioAxi_wd_bits_last ? 1'h0 : 1'h1; // @[playground/src/sim/sim_mmio.scala 135:21 176:46 178:29]
  wire [6:0] _GEN_398 = io_mmioAxi_wd_valid ? _GEN_351 : 7'h0; // @[playground/src/sim/sim_mmio.scala 136:38 47:20]
  wire [63:0] _GEN_399 = io_mmioAxi_wd_valid ? _GEN_352 : 64'h0; // @[playground/src/sim/sim_mmio.scala 136:38 47:96]
  wire  _GEN_400 = io_mmioAxi_wd_valid & _GEN_353; // @[playground/src/sim/sim_mmio.scala 136:38 47:42]
  wire  _GEN_403 = io_mmioAxi_wd_valid & _GEN_356; // @[playground/src/sim/sim_mmio.scala 136:38 55:19]
  wire [7:0] _offset_T_1 = offset + 8'h1; // @[playground/src/sim/sim_mmio.scala 191:35]
  wire  _GEN_422 = islast ? 1'h0 : 1'h1; // @[playground/src/sim/sim_mmio.scala 189:21 192:29 193:29]
  wire [2:0] _GEN_423 = islast ? 3'h0 : state; // @[playground/src/sim/sim_mmio.scala 192:29 194:29 78:24]
  wire [7:0] _GEN_424 = io_mmioAxi_rd_ready & rdvalid ? _offset_T_1 : offset; // @[playground/src/sim/sim_mmio.scala 190:49 191:25 69:26]
  wire  _GEN_425 = io_mmioAxi_rd_ready & rdvalid ? _GEN_422 : 1'h1; // @[playground/src/sim/sim_mmio.scala 189:21 190:49]
  wire [2:0] _GEN_426 = io_mmioAxi_rd_ready & rdvalid ? _GEN_423 : state; // @[playground/src/sim/sim_mmio.scala 190:49 78:24]
  wire [5:0] _rdata_T_13 = {io_mmioAxi_ra_bits_addr[2:0],3'h0}; // @[playground/src/sim/sim_mmio.scala 199:44]
  wire [126:0] _GEN_392 = {{63'd0}, sdcard_rdata}; // @[playground/src/sim/sim_mmio.scala 199:38]
  wire [126:0] _rdata_T_14 = _GEN_392 << _rdata_T_13; // @[playground/src/sim/sim_mmio.scala 199:38]
  wire [126:0] _GEN_427 = 3'h4 == state ? _rdata_T_14 : {{63'd0}, rdata}; // @[playground/src/sim/sim_mmio.scala 85:18 199:19 67:26]
  wire [2:0] _GEN_428 = 3'h4 == state ? 3'h3 : state; // @[playground/src/sim/sim_mmio.scala 85:18 200:19 78:24]
  wire  _GEN_429 = 3'h3 == state ? _GEN_425 : rdvalid; // @[playground/src/sim/sim_mmio.scala 85:18 65:26]
  wire [7:0] _GEN_430 = 3'h3 == state ? _GEN_424 : offset; // @[playground/src/sim/sim_mmio.scala 85:18 69:26]
  wire [2:0] _GEN_431 = 3'h3 == state ? _GEN_426 : _GEN_428; // @[playground/src/sim/sim_mmio.scala 85:18]
  wire [126:0] _GEN_432 = 3'h3 == state ? {{63'd0}, rdata} : _GEN_427; // @[playground/src/sim/sim_mmio.scala 85:18 67:26]
  wire [126:0] _GEN_436 = 3'h2 == state ? {{63'd0}, rdata} : _GEN_432; // @[playground/src/sim/sim_mmio.scala 85:18 67:26]
  wire [6:0] _GEN_461 = 3'h1 == state ? _GEN_398 : 7'h0; // @[playground/src/sim/sim_mmio.scala 85:18 47:20]
  wire [63:0] _GEN_462 = 3'h1 == state ? _GEN_399 : 64'h0; // @[playground/src/sim/sim_mmio.scala 85:18 47:96]
  wire  _GEN_466 = 3'h1 == state & _GEN_403; // @[playground/src/sim/sim_mmio.scala 85:18 55:19]
  wire [126:0] _GEN_486 = 3'h1 == state ? {{63'd0}, rdata} : _GEN_436; // @[playground/src/sim/sim_mmio.scala 85:18 67:26]
  wire [134:0] _GEN_494 = 3'h0 == state ? _GEN_58 : {{8'd0}, _GEN_486}; // @[playground/src/sim/sim_mmio.scala 85:18]
  wire [134:0] _GEN_2 = reset ? 135'h0 : _GEN_494; // @[playground/src/sim/sim_mmio.scala 67:{26,26}]
  wire  _GEN_262 = ~_T_32; // @[playground/src/sim/sim_mmio.scala 129:27]
  wire  _GEN_268 = ~_T_1 & _T_40 & io_mmioAxi_wd_valid; // @[playground/src/sim/sim_mmio.scala 143:31]
  wire  _GEN_300 = _GEN_268 & ~_T_45 & ~_T_54; // @[playground/src/sim/sim_mmio.scala 149:31]
  SdCard sdcard ( // @[playground/src/sim/sim_mmio.scala 46:24]
    .addr(sdcard_addr),
    .wen(sdcard_wen),
    .wdata(sdcard_wdata),
    .clock(sdcard_clock),
    .cen(sdcard_cen),
    .rdata(sdcard_rdata)
  );
  assign disk_disk_rdata_MPORT_en = 1'h1;
  assign disk_disk_rdata_MPORT_addr = _disk_rdata_T_2[25:0];
  assign disk_disk_rdata_MPORT_data = disk[disk_disk_rdata_MPORT_addr]; // @[playground/src/sim/sim_mmio.scala 55:19]
  assign disk_disk_rdata_MPORT_1_en = 1'h1;
  assign disk_disk_rdata_MPORT_1_addr = _disk_rdata_T_6[25:0];
  assign disk_disk_rdata_MPORT_1_data = disk[disk_disk_rdata_MPORT_1_addr]; // @[playground/src/sim/sim_mmio.scala 55:19]
  assign disk_disk_rdata_MPORT_2_en = 1'h1;
  assign disk_disk_rdata_MPORT_2_addr = _disk_rdata_T_10[25:0];
  assign disk_disk_rdata_MPORT_2_data = disk[disk_disk_rdata_MPORT_2_addr]; // @[playground/src/sim/sim_mmio.scala 55:19]
  assign disk_disk_rdata_MPORT_3_en = 1'h1;
  assign disk_disk_rdata_MPORT_3_addr = _disk_rdata_T_14[25:0];
  assign disk_disk_rdata_MPORT_3_data = disk[disk_disk_rdata_MPORT_3_addr]; // @[playground/src/sim/sim_mmio.scala 55:19]
  assign disk_disk_rdata_MPORT_4_en = 1'h1;
  assign disk_disk_rdata_MPORT_4_addr = _disk_rdata_T_18[25:0];
  assign disk_disk_rdata_MPORT_4_data = disk[disk_disk_rdata_MPORT_4_addr]; // @[playground/src/sim/sim_mmio.scala 55:19]
  assign disk_disk_rdata_MPORT_5_en = 1'h1;
  assign disk_disk_rdata_MPORT_5_addr = _disk_rdata_T_22[25:0];
  assign disk_disk_rdata_MPORT_5_data = disk[disk_disk_rdata_MPORT_5_addr]; // @[playground/src/sim/sim_mmio.scala 55:19]
  assign disk_disk_rdata_MPORT_6_en = 1'h1;
  assign disk_disk_rdata_MPORT_6_addr = _disk_rdata_T_26[25:0];
  assign disk_disk_rdata_MPORT_6_data = disk[disk_disk_rdata_MPORT_6_addr]; // @[playground/src/sim/sim_mmio.scala 55:19]
  assign disk_disk_rdata_MPORT_7_en = 1'h1;
  assign disk_disk_rdata_MPORT_7_addr = _disk_rdata_T_30[25:0];
  assign disk_disk_rdata_MPORT_7_data = disk[disk_disk_rdata_MPORT_7_addr]; // @[playground/src/sim/sim_mmio.scala 55:19]
  assign disk_MPORT_4_data = io_mmioAxi_wd_bits_data[7:0];
  assign disk_MPORT_4_addr = _T_121[25:0];
  assign disk_MPORT_4_mask = 1'h1;
  assign disk_MPORT_4_en = _T_1 ? 1'h0 : _GEN_466;
  assign disk_MPORT_5_data = io_mmioAxi_wd_bits_data[15:8];
  assign disk_MPORT_5_addr = _T_126[25:0];
  assign disk_MPORT_5_mask = 1'h1;
  assign disk_MPORT_5_en = _T_1 ? 1'h0 : _GEN_466;
  assign disk_MPORT_6_data = io_mmioAxi_wd_bits_data[23:16];
  assign disk_MPORT_6_addr = _T_130[25:0];
  assign disk_MPORT_6_mask = 1'h1;
  assign disk_MPORT_6_en = _T_1 ? 1'h0 : _GEN_466;
  assign disk_MPORT_7_data = io_mmioAxi_wd_bits_data[31:24];
  assign disk_MPORT_7_addr = _T_134[25:0];
  assign disk_MPORT_7_mask = 1'h1;
  assign disk_MPORT_7_en = _T_1 ? 1'h0 : _GEN_466;
  assign disk_MPORT_8_data = io_mmioAxi_wd_bits_data[39:32];
  assign disk_MPORT_8_addr = _T_138[25:0];
  assign disk_MPORT_8_mask = 1'h1;
  assign disk_MPORT_8_en = _T_1 ? 1'h0 : _GEN_466;
  assign disk_MPORT_9_data = io_mmioAxi_wd_bits_data[47:40];
  assign disk_MPORT_9_addr = _T_142[25:0];
  assign disk_MPORT_9_mask = 1'h1;
  assign disk_MPORT_9_en = _T_1 ? 1'h0 : _GEN_466;
  assign disk_MPORT_10_data = io_mmioAxi_wd_bits_data[55:48];
  assign disk_MPORT_10_addr = _T_146[25:0];
  assign disk_MPORT_10_mask = 1'h1;
  assign disk_MPORT_10_en = _T_1 ? 1'h0 : _GEN_466;
  assign disk_MPORT_11_data = io_mmioAxi_wd_bits_data[63:56];
  assign disk_MPORT_11_addr = _T_150[25:0];
  assign disk_MPORT_11_mask = 1'h1;
  assign disk_MPORT_11_en = _T_1 ? 1'h0 : _GEN_466;
  assign flash_flash_rdata_MPORT_en = 1'h1;
  assign flash_flash_rdata_MPORT_addr = _flash_rdata_T_2[27:0];
  assign flash_flash_rdata_MPORT_data = flash[flash_flash_rdata_MPORT_addr]; // @[playground/src/sim/sim_mmio.scala 56:20]
  assign flash_flash_rdata_MPORT_1_en = 1'h1;
  assign flash_flash_rdata_MPORT_1_addr = _flash_rdata_T_6[27:0];
  assign flash_flash_rdata_MPORT_1_data = flash[flash_flash_rdata_MPORT_1_addr]; // @[playground/src/sim/sim_mmio.scala 56:20]
  assign flash_flash_rdata_MPORT_2_en = 1'h1;
  assign flash_flash_rdata_MPORT_2_addr = _flash_rdata_T_10[27:0];
  assign flash_flash_rdata_MPORT_2_data = flash[flash_flash_rdata_MPORT_2_addr]; // @[playground/src/sim/sim_mmio.scala 56:20]
  assign flash_flash_rdata_MPORT_3_en = 1'h1;
  assign flash_flash_rdata_MPORT_3_addr = _flash_rdata_T_14[27:0];
  assign flash_flash_rdata_MPORT_3_data = flash[flash_flash_rdata_MPORT_3_addr]; // @[playground/src/sim/sim_mmio.scala 56:20]
  assign flash_flash_rdata_MPORT_4_en = 1'h1;
  assign flash_flash_rdata_MPORT_4_addr = _flash_rdata_T_18[27:0];
  assign flash_flash_rdata_MPORT_4_data = flash[flash_flash_rdata_MPORT_4_addr]; // @[playground/src/sim/sim_mmio.scala 56:20]
  assign flash_flash_rdata_MPORT_5_en = 1'h1;
  assign flash_flash_rdata_MPORT_5_addr = _flash_rdata_T_22[27:0];
  assign flash_flash_rdata_MPORT_5_data = flash[flash_flash_rdata_MPORT_5_addr]; // @[playground/src/sim/sim_mmio.scala 56:20]
  assign flash_flash_rdata_MPORT_6_en = 1'h1;
  assign flash_flash_rdata_MPORT_6_addr = _flash_rdata_T_26[27:0];
  assign flash_flash_rdata_MPORT_6_data = flash[flash_flash_rdata_MPORT_6_addr]; // @[playground/src/sim/sim_mmio.scala 56:20]
  assign flash_flash_rdata_MPORT_7_en = 1'h1;
  assign flash_flash_rdata_MPORT_7_addr = _flash_rdata_T_29[27:0];
  assign flash_flash_rdata_MPORT_7_data = flash[flash_flash_rdata_MPORT_7_addr]; // @[playground/src/sim/sim_mmio.scala 56:20]
  assign io_mmioAxi_wa_ready = waready; // @[playground/src/sim/sim_mmio.scala 207:25]
  assign io_mmioAxi_wd_ready = wdready; // @[playground/src/sim/sim_mmio.scala 208:25]
  assign io_mmioAxi_ra_ready = raready; // @[playground/src/sim/sim_mmio.scala 209:25]
  assign io_mmioAxi_rd_valid = rdvalid; // @[playground/src/sim/sim_mmio.scala 210:25]
  assign io_mmioAxi_rd_bits_data = rdata; // @[playground/src/sim/sim_mmio.scala 211:29]
  assign io_mmioAxi_rd_bits_last = offset == 8'h0; // @[playground/src/sim/sim_mmio.scala 79:27]
  assign sdcard_addr = 3'h0 == state ? _GEN_59 : _GEN_461; // @[playground/src/sim/sim_mmio.scala 85:18]
  assign sdcard_wen = 3'h0 == state ? 1'h0 : 3'h1 == state & _GEN_400; // @[playground/src/sim/sim_mmio.scala 85:18 47:42]
  assign sdcard_wdata = 3'h0 == state ? 64'h0 : _GEN_462; // @[playground/src/sim/sim_mmio.scala 85:18 47:96]
  assign sdcard_clock = clock; // @[playground/src/sim/sim_mmio.scala 48:21]
  assign sdcard_cen = 3'h0 == state & _GEN_60; // @[playground/src/sim/sim_mmio.scala 85:18 47:68]
  always @(posedge clock) begin
    if (disk_MPORT_4_en & disk_MPORT_4_mask) begin
      disk[disk_MPORT_4_addr] <= disk_MPORT_4_data; // @[playground/src/sim/sim_mmio.scala 55:19]
    end
    if (disk_MPORT_5_en & disk_MPORT_5_mask) begin
      disk[disk_MPORT_5_addr] <= disk_MPORT_5_data; // @[playground/src/sim/sim_mmio.scala 55:19]
    end
    if (disk_MPORT_6_en & disk_MPORT_6_mask) begin
      disk[disk_MPORT_6_addr] <= disk_MPORT_6_data; // @[playground/src/sim/sim_mmio.scala 55:19]
    end
    if (disk_MPORT_7_en & disk_MPORT_7_mask) begin
      disk[disk_MPORT_7_addr] <= disk_MPORT_7_data; // @[playground/src/sim/sim_mmio.scala 55:19]
    end
    if (disk_MPORT_8_en & disk_MPORT_8_mask) begin
      disk[disk_MPORT_8_addr] <= disk_MPORT_8_data; // @[playground/src/sim/sim_mmio.scala 55:19]
    end
    if (disk_MPORT_9_en & disk_MPORT_9_mask) begin
      disk[disk_MPORT_9_addr] <= disk_MPORT_9_data; // @[playground/src/sim/sim_mmio.scala 55:19]
    end
    if (disk_MPORT_10_en & disk_MPORT_10_mask) begin
      disk[disk_MPORT_10_addr] <= disk_MPORT_10_data; // @[playground/src/sim/sim_mmio.scala 55:19]
    end
    if (disk_MPORT_11_en & disk_MPORT_11_mask) begin
      disk[disk_MPORT_11_addr] <= disk_MPORT_11_data; // @[playground/src/sim/sim_mmio.scala 55:19]
    end
    if (reset) begin // @[playground/src/sim/sim_mmio.scala 50:23]
      uart_0 <= 8'h0; // @[playground/src/sim/sim_mmio.scala 50:23]
    end else if (!(3'h0 == state)) begin // @[playground/src/sim/sim_mmio.scala 85:18]
      if (3'h1 == state) begin // @[playground/src/sim/sim_mmio.scala 85:18]
        if (io_mmioAxi_wd_valid) begin // @[playground/src/sim/sim_mmio.scala 136:38]
          uart_0 <= _GEN_329;
        end
      end
    end
    if (reset) begin // @[playground/src/sim/sim_mmio.scala 50:23]
      uart_1 <= 8'h0; // @[playground/src/sim/sim_mmio.scala 50:23]
    end else if (!(3'h0 == state)) begin // @[playground/src/sim/sim_mmio.scala 85:18]
      if (3'h1 == state) begin // @[playground/src/sim/sim_mmio.scala 85:18]
        if (io_mmioAxi_wd_valid) begin // @[playground/src/sim/sim_mmio.scala 136:38]
          uart_1 <= _GEN_330;
        end
      end
    end
    if (reset) begin // @[playground/src/sim/sim_mmio.scala 50:23]
      uart_2 <= 8'h0; // @[playground/src/sim/sim_mmio.scala 50:23]
    end else if (!(3'h0 == state)) begin // @[playground/src/sim/sim_mmio.scala 85:18]
      if (3'h1 == state) begin // @[playground/src/sim/sim_mmio.scala 85:18]
        if (io_mmioAxi_wd_valid) begin // @[playground/src/sim/sim_mmio.scala 136:38]
          uart_2 <= _GEN_331;
        end
      end
    end
    if (reset) begin // @[playground/src/sim/sim_mmio.scala 50:23]
      uart_3 <= 8'h0; // @[playground/src/sim/sim_mmio.scala 50:23]
    end else if (!(3'h0 == state)) begin // @[playground/src/sim/sim_mmio.scala 85:18]
      if (3'h1 == state) begin // @[playground/src/sim/sim_mmio.scala 85:18]
        if (io_mmioAxi_wd_valid) begin // @[playground/src/sim/sim_mmio.scala 136:38]
          uart_3 <= _GEN_332;
        end
      end
    end
    if (reset) begin // @[playground/src/sim/sim_mmio.scala 50:23]
      uart_4 <= 8'h0; // @[playground/src/sim/sim_mmio.scala 50:23]
    end else if (!(3'h0 == state)) begin // @[playground/src/sim/sim_mmio.scala 85:18]
      if (3'h1 == state) begin // @[playground/src/sim/sim_mmio.scala 85:18]
        if (io_mmioAxi_wd_valid) begin // @[playground/src/sim/sim_mmio.scala 136:38]
          uart_4 <= _GEN_333;
        end
      end
    end
    if (reset) begin // @[playground/src/sim/sim_mmio.scala 50:23]
      uart_5 <= 8'h0; // @[playground/src/sim/sim_mmio.scala 50:23]
    end else if (3'h0 == state) begin // @[playground/src/sim/sim_mmio.scala 85:18]
      uart_5 <= 8'h20; // @[playground/src/sim/sim_mmio.scala 84:13]
    end else if (3'h1 == state) begin // @[playground/src/sim/sim_mmio.scala 85:18]
      if (io_mmioAxi_wd_valid) begin // @[playground/src/sim/sim_mmio.scala 136:38]
        uart_5 <= _GEN_334;
      end else begin
        uart_5 <= 8'h20; // @[playground/src/sim/sim_mmio.scala 84:13]
      end
    end else begin
      uart_5 <= 8'h20; // @[playground/src/sim/sim_mmio.scala 84:13]
    end
    if (reset) begin // @[playground/src/sim/sim_mmio.scala 50:23]
      uart_6 <= 8'h0; // @[playground/src/sim/sim_mmio.scala 50:23]
    end else if (!(3'h0 == state)) begin // @[playground/src/sim/sim_mmio.scala 85:18]
      if (3'h1 == state) begin // @[playground/src/sim/sim_mmio.scala 85:18]
        if (io_mmioAxi_wd_valid) begin // @[playground/src/sim/sim_mmio.scala 136:38]
          uart_6 <= _GEN_335;
        end
      end
    end
    if (reset) begin // @[playground/src/sim/sim_mmio.scala 50:23]
      uart_7 <= 8'h0; // @[playground/src/sim/sim_mmio.scala 50:23]
    end else if (!(3'h0 == state)) begin // @[playground/src/sim/sim_mmio.scala 85:18]
      if (3'h1 == state) begin // @[playground/src/sim/sim_mmio.scala 85:18]
        if (io_mmioAxi_wd_valid) begin // @[playground/src/sim/sim_mmio.scala 136:38]
          uart_7 <= _GEN_336;
        end
      end
    end
    if (reset) begin // @[playground/src/sim/sim_mmio.scala 51:24]
      mtime <= 64'h0; // @[playground/src/sim/sim_mmio.scala 51:24]
    end else begin
      mtime <= _mtime_T_1;
    end
    if (reset) begin // @[playground/src/sim/sim_mmio.scala 52:27]
      mtimecmp <= 64'h0; // @[playground/src/sim/sim_mmio.scala 52:27]
    end else if (!(3'h0 == state)) begin // @[playground/src/sim/sim_mmio.scala 85:18]
      if (3'h1 == state) begin // @[playground/src/sim/sim_mmio.scala 85:18]
        if (io_mmioAxi_wd_valid) begin // @[playground/src/sim/sim_mmio.scala 136:38]
          mtimecmp <= _GEN_337;
        end
      end
    end
    if (reset) begin // @[playground/src/sim/sim_mmio.scala 58:27]
      waready <= 1'h0; // @[playground/src/sim/sim_mmio.scala 58:27]
    end else if (3'h0 == state) begin // @[playground/src/sim/sim_mmio.scala 85:18]
      if (io_mmioAxi_wa_valid & waready) begin // @[playground/src/sim/sim_mmio.scala 90:49]
        waready <= 1'h0; // @[playground/src/sim/sim_mmio.scala 93:26]
      end else begin
        waready <= 1'h1; // @[playground/src/sim/sim_mmio.scala 87:21]
      end
    end
    if (reset) begin // @[playground/src/sim/sim_mmio.scala 59:27]
      wdready <= 1'h0; // @[playground/src/sim/sim_mmio.scala 59:27]
    end else if (!(3'h0 == state)) begin // @[playground/src/sim/sim_mmio.scala 85:18]
      if (3'h1 == state) begin // @[playground/src/sim/sim_mmio.scala 85:18]
        if (io_mmioAxi_wd_valid) begin // @[playground/src/sim/sim_mmio.scala 136:38]
          wdready <= _GEN_374;
        end else begin
          wdready <= 1'h1; // @[playground/src/sim/sim_mmio.scala 135:21]
        end
      end
    end
    if (reset) begin // @[playground/src/sim/sim_mmio.scala 60:26]
      waddr <= 32'h0; // @[playground/src/sim/sim_mmio.scala 60:26]
    end else if (3'h0 == state) begin // @[playground/src/sim/sim_mmio.scala 85:18]
      if (io_mmioAxi_wa_valid & waready) begin // @[playground/src/sim/sim_mmio.scala 90:49]
        waddr <= io_mmioAxi_wa_bits_addr; // @[playground/src/sim/sim_mmio.scala 91:25]
      end
    end
    if (reset) begin // @[playground/src/sim/sim_mmio.scala 64:26]
      raready <= 1'h0; // @[playground/src/sim/sim_mmio.scala 64:26]
    end else if (3'h0 == state) begin // @[playground/src/sim/sim_mmio.scala 85:18]
      if (io_mmioAxi_ra_valid & raready) begin // @[playground/src/sim/sim_mmio.scala 96:49]
        raready <= 1'h0; // @[playground/src/sim/sim_mmio.scala 98:25]
      end else begin
        raready <= 1'h1; // @[playground/src/sim/sim_mmio.scala 88:21]
      end
    end
    if (reset) begin // @[playground/src/sim/sim_mmio.scala 65:26]
      rdvalid <= 1'h0; // @[playground/src/sim/sim_mmio.scala 65:26]
    end else if (!(3'h0 == state)) begin // @[playground/src/sim/sim_mmio.scala 85:18]
      if (!(3'h1 == state)) begin // @[playground/src/sim/sim_mmio.scala 85:18]
        if (!(3'h2 == state)) begin // @[playground/src/sim/sim_mmio.scala 85:18]
          rdvalid <= _GEN_429;
        end
      end
    end
    rdata <= _GEN_2[63:0]; // @[playground/src/sim/sim_mmio.scala 67:{26,26}]
    if (reset) begin // @[playground/src/sim/sim_mmio.scala 69:26]
      offset <= 8'h0; // @[playground/src/sim/sim_mmio.scala 69:26]
    end else if (3'h0 == state) begin // @[playground/src/sim/sim_mmio.scala 85:18]
      offset <= 8'h0; // @[playground/src/sim/sim_mmio.scala 89:21]
    end else if (!(3'h1 == state)) begin // @[playground/src/sim/sim_mmio.scala 85:18]
      if (!(3'h2 == state)) begin // @[playground/src/sim/sim_mmio.scala 85:18]
        offset <= _GEN_430;
      end
    end
    if (reset) begin // @[playground/src/sim/sim_mmio.scala 78:24]
      state <= 3'h0; // @[playground/src/sim/sim_mmio.scala 78:24]
    end else if (3'h0 == state) begin // @[playground/src/sim/sim_mmio.scala 85:18]
      if (io_mmioAxi_ra_valid & raready) begin // @[playground/src/sim/sim_mmio.scala 96:49]
        if (io_mmioAxi_ra_bits_addr >= 32'h10000000 & io_mmioAxi_ra_bits_addr <= 32'h10000007) begin // @[playground/src/sim/sim_mmio.scala 100:115]
          state <= 3'h3; // @[playground/src/sim/sim_mmio.scala 99:25]
        end else begin
          state <= _GEN_50;
        end
      end else if (io_mmioAxi_wa_valid & waready) begin // @[playground/src/sim/sim_mmio.scala 90:49]
        state <= 3'h1; // @[playground/src/sim/sim_mmio.scala 94:25]
      end
    end else if (3'h1 == state) begin // @[playground/src/sim/sim_mmio.scala 85:18]
      if (io_mmioAxi_wd_valid) begin // @[playground/src/sim/sim_mmio.scala 136:38]
        state <= _GEN_373;
      end
    end else if (3'h2 == state) begin // @[playground/src/sim/sim_mmio.scala 85:18]
      state <= 3'h0; // @[playground/src/sim/sim_mmio.scala 185:19]
    end else begin
      state <= _GEN_431;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1 & _T_3 & ~_T_8 & ~_T_9 & ~_T_10 & ~_T_11 & ~_T_12 & ~_T_15 & ~_T_16 & ~_T_17 & ~_T_22 & ~_T_27 & ~_T_32
           & ~_T_37 & ~reset) begin
          $fwrite(32'h80000002,"mmio invalid raddr: %x\n",io_mmioAxi_ra_bits_addr); // @[playground/src/sim/sim_mmio.scala 129:27]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~_T_1 & _T_40 & io_mmioAxi_wd_valid & _T_45 & _T_50 & _T_39) begin
          $fwrite(32'h80000002,"%c",inputwd[7:0]); // @[playground/src/sim/sim_mmio.scala 143:31]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_268 & ~_T_45 & ~_T_54 & _T_55 & _T_39) begin
          $fwrite(32'h80000002,"%c",inputwd[7:0]); // @[playground/src/sim/sim_mmio.scala 149:31]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_300 & ~_T_55 & ~_T_63 & ~_T_100 & ~_T_101 & ~_T_104 & ~_T_105 & ~_T_110 & ~_T_115 & _GEN_262 & _T_39
          ) begin
          $fwrite(32'h80000002,"mmio invalid waddr: %x\n",io_mmioAxi_wa_bits_addr); // @[playground/src/sim/sim_mmio.scala 173:31]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 67108864; initvar = initvar+1)
    disk[initvar] = _RAND_0[7:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 268435456; initvar = initvar+1)
    flash[initvar] = _RAND_1[7:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  uart_0 = _RAND_2[7:0];
  _RAND_3 = {1{`RANDOM}};
  uart_1 = _RAND_3[7:0];
  _RAND_4 = {1{`RANDOM}};
  uart_2 = _RAND_4[7:0];
  _RAND_5 = {1{`RANDOM}};
  uart_3 = _RAND_5[7:0];
  _RAND_6 = {1{`RANDOM}};
  uart_4 = _RAND_6[7:0];
  _RAND_7 = {1{`RANDOM}};
  uart_5 = _RAND_7[7:0];
  _RAND_8 = {1{`RANDOM}};
  uart_6 = _RAND_8[7:0];
  _RAND_9 = {1{`RANDOM}};
  uart_7 = _RAND_9[7:0];
  _RAND_10 = {2{`RANDOM}};
  mtime = _RAND_10[63:0];
  _RAND_11 = {2{`RANDOM}};
  mtimecmp = _RAND_11[63:0];
  _RAND_12 = {1{`RANDOM}};
  waready = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  wdready = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  waddr = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  raready = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  rdvalid = _RAND_16[0:0];
  _RAND_17 = {2{`RANDOM}};
  rdata = _RAND_17[63:0];
  _RAND_18 = {1{`RANDOM}};
  offset = _RAND_18[7:0];
  _RAND_19 = {1{`RANDOM}};
  state = _RAND_19[2:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module SimDma(
  input        clock,
  input        reset,
  output [7:0] io_dmaAxi_wstrb // @[playground/src/sim/sim_dma.scala 13:16]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  reg [7:0] wstrb_r; // @[playground/src/sim/sim_dma.scala 39:30]
  wire [8:0] _GEN_33 = {{1'd0}, wstrb_r}; // @[playground/src/sim/sim_dma.scala 101:25 39:30 99:47]
  wire [8:0] _GEN_99 = reset ? 9'h0 : _GEN_33; // @[playground/src/sim/sim_dma.scala 39:{30,30}]
  assign io_dmaAxi_wstrb = wstrb_r; // @[playground/src/sim/sim_dma.scala 127:25]
  always @(posedge clock) begin
    wstrb_r <= _GEN_99[7:0]; // @[playground/src/sim/sim_dma.scala 39:{30,30}]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  wstrb_r = _RAND_0[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module SimCrossbar(
  input         clock,
  input         reset,
  output        io_inAxi_wa_ready, // @[playground/src/sim/sim_crossbar.scala 10:16]
  input         io_inAxi_wa_valid, // @[playground/src/sim/sim_crossbar.scala 10:16]
  input  [3:0]  io_inAxi_wa_bits_id, // @[playground/src/sim/sim_crossbar.scala 10:16]
  input  [31:0] io_inAxi_wa_bits_addr, // @[playground/src/sim/sim_crossbar.scala 10:16]
  input  [7:0]  io_inAxi_wa_bits_len, // @[playground/src/sim/sim_crossbar.scala 10:16]
  input  [2:0]  io_inAxi_wa_bits_size, // @[playground/src/sim/sim_crossbar.scala 10:16]
  input  [1:0]  io_inAxi_wa_bits_burst, // @[playground/src/sim/sim_crossbar.scala 10:16]
  output        io_inAxi_wd_ready, // @[playground/src/sim/sim_crossbar.scala 10:16]
  input         io_inAxi_wd_valid, // @[playground/src/sim/sim_crossbar.scala 10:16]
  input  [63:0] io_inAxi_wd_bits_data, // @[playground/src/sim/sim_crossbar.scala 10:16]
  input  [7:0]  io_inAxi_wd_bits_strb, // @[playground/src/sim/sim_crossbar.scala 10:16]
  input         io_inAxi_wd_bits_last, // @[playground/src/sim/sim_crossbar.scala 10:16]
  input         io_inAxi_wr_ready, // @[playground/src/sim/sim_crossbar.scala 10:16]
  output        io_inAxi_wr_valid, // @[playground/src/sim/sim_crossbar.scala 10:16]
  output [3:0]  io_inAxi_wr_bits_id, // @[playground/src/sim/sim_crossbar.scala 10:16]
  output [1:0]  io_inAxi_wr_bits_resp, // @[playground/src/sim/sim_crossbar.scala 10:16]
  output        io_inAxi_ra_ready, // @[playground/src/sim/sim_crossbar.scala 10:16]
  input         io_inAxi_ra_valid, // @[playground/src/sim/sim_crossbar.scala 10:16]
  input  [3:0]  io_inAxi_ra_bits_id, // @[playground/src/sim/sim_crossbar.scala 10:16]
  input  [31:0] io_inAxi_ra_bits_addr, // @[playground/src/sim/sim_crossbar.scala 10:16]
  input  [7:0]  io_inAxi_ra_bits_len, // @[playground/src/sim/sim_crossbar.scala 10:16]
  input  [2:0]  io_inAxi_ra_bits_size, // @[playground/src/sim/sim_crossbar.scala 10:16]
  input  [1:0]  io_inAxi_ra_bits_burst, // @[playground/src/sim/sim_crossbar.scala 10:16]
  input         io_inAxi_rd_ready, // @[playground/src/sim/sim_crossbar.scala 10:16]
  output        io_inAxi_rd_valid, // @[playground/src/sim/sim_crossbar.scala 10:16]
  output [3:0]  io_inAxi_rd_bits_id, // @[playground/src/sim/sim_crossbar.scala 10:16]
  output [63:0] io_inAxi_rd_bits_data, // @[playground/src/sim/sim_crossbar.scala 10:16]
  output [1:0]  io_inAxi_rd_bits_resp, // @[playground/src/sim/sim_crossbar.scala 10:16]
  output        io_inAxi_rd_bits_last, // @[playground/src/sim/sim_crossbar.scala 10:16]
  input         io_memAxi_wa_ready, // @[playground/src/sim/sim_crossbar.scala 10:16]
  output        io_memAxi_wa_valid, // @[playground/src/sim/sim_crossbar.scala 10:16]
  output [3:0]  io_memAxi_wa_bits_id, // @[playground/src/sim/sim_crossbar.scala 10:16]
  output [31:0] io_memAxi_wa_bits_addr, // @[playground/src/sim/sim_crossbar.scala 10:16]
  output [7:0]  io_memAxi_wa_bits_len, // @[playground/src/sim/sim_crossbar.scala 10:16]
  output [2:0]  io_memAxi_wa_bits_size, // @[playground/src/sim/sim_crossbar.scala 10:16]
  output [1:0]  io_memAxi_wa_bits_burst, // @[playground/src/sim/sim_crossbar.scala 10:16]
  input         io_memAxi_wd_ready, // @[playground/src/sim/sim_crossbar.scala 10:16]
  output        io_memAxi_wd_valid, // @[playground/src/sim/sim_crossbar.scala 10:16]
  output [63:0] io_memAxi_wd_bits_data, // @[playground/src/sim/sim_crossbar.scala 10:16]
  output [7:0]  io_memAxi_wd_bits_strb, // @[playground/src/sim/sim_crossbar.scala 10:16]
  output        io_memAxi_wd_bits_last, // @[playground/src/sim/sim_crossbar.scala 10:16]
  output        io_memAxi_wr_ready, // @[playground/src/sim/sim_crossbar.scala 10:16]
  input         io_memAxi_wr_valid, // @[playground/src/sim/sim_crossbar.scala 10:16]
  input  [3:0]  io_memAxi_wr_bits_id, // @[playground/src/sim/sim_crossbar.scala 10:16]
  input  [1:0]  io_memAxi_wr_bits_resp, // @[playground/src/sim/sim_crossbar.scala 10:16]
  input         io_memAxi_ra_ready, // @[playground/src/sim/sim_crossbar.scala 10:16]
  output        io_memAxi_ra_valid, // @[playground/src/sim/sim_crossbar.scala 10:16]
  output [3:0]  io_memAxi_ra_bits_id, // @[playground/src/sim/sim_crossbar.scala 10:16]
  output [31:0] io_memAxi_ra_bits_addr, // @[playground/src/sim/sim_crossbar.scala 10:16]
  output [7:0]  io_memAxi_ra_bits_len, // @[playground/src/sim/sim_crossbar.scala 10:16]
  output [2:0]  io_memAxi_ra_bits_size, // @[playground/src/sim/sim_crossbar.scala 10:16]
  output [1:0]  io_memAxi_ra_bits_burst, // @[playground/src/sim/sim_crossbar.scala 10:16]
  output        io_memAxi_rd_ready, // @[playground/src/sim/sim_crossbar.scala 10:16]
  input         io_memAxi_rd_valid, // @[playground/src/sim/sim_crossbar.scala 10:16]
  input  [3:0]  io_memAxi_rd_bits_id, // @[playground/src/sim/sim_crossbar.scala 10:16]
  input  [63:0] io_memAxi_rd_bits_data, // @[playground/src/sim/sim_crossbar.scala 10:16]
  input  [1:0]  io_memAxi_rd_bits_resp, // @[playground/src/sim/sim_crossbar.scala 10:16]
  input         io_memAxi_rd_bits_last, // @[playground/src/sim/sim_crossbar.scala 10:16]
  input         io_mmioAxi_wa_ready, // @[playground/src/sim/sim_crossbar.scala 10:16]
  output        io_mmioAxi_wa_valid, // @[playground/src/sim/sim_crossbar.scala 10:16]
  output [31:0] io_mmioAxi_wa_bits_addr, // @[playground/src/sim/sim_crossbar.scala 10:16]
  input         io_mmioAxi_wd_ready, // @[playground/src/sim/sim_crossbar.scala 10:16]
  output        io_mmioAxi_wd_valid, // @[playground/src/sim/sim_crossbar.scala 10:16]
  output [63:0] io_mmioAxi_wd_bits_data, // @[playground/src/sim/sim_crossbar.scala 10:16]
  output [7:0]  io_mmioAxi_wd_bits_strb, // @[playground/src/sim/sim_crossbar.scala 10:16]
  output        io_mmioAxi_wd_bits_last, // @[playground/src/sim/sim_crossbar.scala 10:16]
  input         io_mmioAxi_ra_ready, // @[playground/src/sim/sim_crossbar.scala 10:16]
  output        io_mmioAxi_ra_valid, // @[playground/src/sim/sim_crossbar.scala 10:16]
  output [31:0] io_mmioAxi_ra_bits_addr, // @[playground/src/sim/sim_crossbar.scala 10:16]
  output        io_mmioAxi_rd_ready, // @[playground/src/sim/sim_crossbar.scala 10:16]
  input         io_mmioAxi_rd_valid, // @[playground/src/sim/sim_crossbar.scala 10:16]
  input  [63:0] io_mmioAxi_rd_bits_data, // @[playground/src/sim/sim_crossbar.scala 10:16]
  input         io_mmioAxi_rd_bits_last // @[playground/src/sim/sim_crossbar.scala 10:16]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  reg [1:0] state; // @[playground/src/sim/sim_crossbar.scala 19:24]
  wire  _GEN_1 = (io_inAxi_ra_valid | io_inAxi_wa_valid) & io_inAxi_rd_ready; // @[playground/src/sim/sim_crossbar.scala 28:63 30:26 playground/src/axi/axi.scala 87:18]
  wire  _GEN_2 = (io_inAxi_ra_valid | io_inAxi_wa_valid) & io_memAxi_rd_valid; // @[playground/src/axi/axi.scala 105:18 playground/src/sim/sim_crossbar.scala 28:63 30:26]
  wire [3:0] _GEN_3 = io_inAxi_ra_valid | io_inAxi_wa_valid ? io_memAxi_rd_bits_id : 4'h0; // @[playground/src/sim/sim_crossbar.scala 28:63 30:26 playground/src/axi/axi.scala 68:23]
  wire [63:0] _GEN_4 = io_inAxi_ra_valid | io_inAxi_wa_valid ? io_memAxi_rd_bits_data : 64'h0; // @[playground/src/sim/sim_crossbar.scala 28:63 30:26 playground/src/axi/axi.scala 68:23]
  wire [1:0] _GEN_5 = io_inAxi_ra_valid | io_inAxi_wa_valid ? io_memAxi_rd_bits_resp : 2'h0; // @[playground/src/sim/sim_crossbar.scala 28:63 30:26 playground/src/axi/axi.scala 68:23]
  wire  _GEN_6 = (io_inAxi_ra_valid | io_inAxi_wa_valid) & io_memAxi_rd_bits_last; // @[playground/src/sim/sim_crossbar.scala 28:63 30:26 playground/src/axi/axi.scala 68:23]
  wire  _GEN_7 = io_inAxi_ra_valid | io_inAxi_wa_valid ? io_memAxi_ra_ready : 1'h1; // @[playground/src/sim/sim_crossbar.scala 28:63 30:26 22:31]
  wire  _GEN_8 = (io_inAxi_ra_valid | io_inAxi_wa_valid) & io_inAxi_ra_valid; // @[playground/src/sim/sim_crossbar.scala 28:63 30:26 playground/src/axi/axi.scala 86:18]
  wire [3:0] _GEN_9 = io_inAxi_ra_valid | io_inAxi_wa_valid ? io_inAxi_ra_bits_id : 4'h0; // @[playground/src/sim/sim_crossbar.scala 28:63 30:26 playground/src/axi/axi.scala 41:23]
  wire [31:0] _GEN_10 = io_inAxi_ra_valid | io_inAxi_wa_valid ? io_inAxi_ra_bits_addr : 32'h0; // @[playground/src/sim/sim_crossbar.scala 28:63 30:26 playground/src/axi/axi.scala 41:23]
  wire [7:0] _GEN_11 = io_inAxi_ra_valid | io_inAxi_wa_valid ? io_inAxi_ra_bits_len : 8'h0; // @[playground/src/sim/sim_crossbar.scala 28:63 30:26 playground/src/axi/axi.scala 41:23]
  wire [2:0] _GEN_12 = io_inAxi_ra_valid | io_inAxi_wa_valid ? io_inAxi_ra_bits_size : 3'h0; // @[playground/src/sim/sim_crossbar.scala 28:63 30:26 playground/src/axi/axi.scala 41:23]
  wire [1:0] _GEN_13 = io_inAxi_ra_valid | io_inAxi_wa_valid ? io_inAxi_ra_bits_burst : 2'h0; // @[playground/src/sim/sim_crossbar.scala 28:63 30:26 playground/src/axi/axi.scala 41:23]
  wire  _GEN_14 = (io_inAxi_ra_valid | io_inAxi_wa_valid) & io_inAxi_wr_ready; // @[playground/src/sim/sim_crossbar.scala 28:63 30:26 playground/src/axi/axi.scala 85:18]
  wire  _GEN_15 = io_inAxi_ra_valid | io_inAxi_wa_valid ? io_memAxi_wr_valid : 1'h1; // @[playground/src/sim/sim_crossbar.scala 28:63 30:26 24:31]
  wire [3:0] _GEN_16 = io_inAxi_ra_valid | io_inAxi_wa_valid ? io_memAxi_wr_bits_id : 4'h0; // @[playground/src/sim/sim_crossbar.scala 28:63 30:26 playground/src/axi/axi.scala 58:23]
  wire [1:0] _GEN_17 = io_inAxi_ra_valid | io_inAxi_wa_valid ? io_memAxi_wr_bits_resp : 2'h0; // @[playground/src/sim/sim_crossbar.scala 28:63 30:26 playground/src/axi/axi.scala 58:23]
  wire  _GEN_18 = (io_inAxi_ra_valid | io_inAxi_wa_valid) & io_memAxi_wd_ready; // @[playground/src/axi/axi.scala 102:18 playground/src/sim/sim_crossbar.scala 28:63 30:26]
  wire  _GEN_19 = (io_inAxi_ra_valid | io_inAxi_wa_valid) & io_inAxi_wd_valid; // @[playground/src/sim/sim_crossbar.scala 28:63 30:26 playground/src/axi/axi.scala 84:18]
  wire [63:0] _GEN_20 = io_inAxi_ra_valid | io_inAxi_wa_valid ? io_inAxi_wd_bits_data : 64'h0; // @[playground/src/sim/sim_crossbar.scala 28:63 30:26 playground/src/axi/axi.scala 50:23]
  wire [7:0] _GEN_21 = io_inAxi_ra_valid | io_inAxi_wa_valid ? io_inAxi_wd_bits_strb : 8'h0; // @[playground/src/sim/sim_crossbar.scala 28:63 30:26 playground/src/axi/axi.scala 50:23]
  wire  _GEN_22 = (io_inAxi_ra_valid | io_inAxi_wa_valid) & io_inAxi_wd_bits_last; // @[playground/src/sim/sim_crossbar.scala 28:63 30:26 playground/src/axi/axi.scala 50:23]
  wire  _GEN_23 = io_inAxi_ra_valid | io_inAxi_wa_valid ? io_memAxi_wa_ready : 1'h1; // @[playground/src/sim/sim_crossbar.scala 28:63 30:26 23:31]
  wire  _GEN_24 = (io_inAxi_ra_valid | io_inAxi_wa_valid) & io_inAxi_wa_valid; // @[playground/src/sim/sim_crossbar.scala 28:63 30:26 playground/src/axi/axi.scala 83:18]
  wire [3:0] _GEN_25 = io_inAxi_ra_valid | io_inAxi_wa_valid ? io_inAxi_wa_bits_id : 4'h0; // @[playground/src/sim/sim_crossbar.scala 28:63 30:26 playground/src/axi/axi.scala 41:23]
  wire [31:0] _GEN_26 = io_inAxi_ra_valid | io_inAxi_wa_valid ? io_inAxi_wa_bits_addr : 32'h0; // @[playground/src/sim/sim_crossbar.scala 28:63 30:26 playground/src/axi/axi.scala 41:23]
  wire [7:0] _GEN_27 = io_inAxi_ra_valid | io_inAxi_wa_valid ? io_inAxi_wa_bits_len : 8'h0; // @[playground/src/sim/sim_crossbar.scala 28:63 30:26 playground/src/axi/axi.scala 41:23]
  wire [2:0] _GEN_28 = io_inAxi_ra_valid | io_inAxi_wa_valid ? io_inAxi_wa_bits_size : 3'h0; // @[playground/src/sim/sim_crossbar.scala 28:63 30:26 playground/src/axi/axi.scala 41:23]
  wire [1:0] _GEN_29 = io_inAxi_ra_valid | io_inAxi_wa_valid ? io_inAxi_wa_bits_burst : 2'h0; // @[playground/src/sim/sim_crossbar.scala 28:63 30:26 playground/src/axi/axi.scala 41:23]
  wire  _GEN_31 = (io_inAxi_ra_valid & (io_inAxi_ra_bits_addr > 32'h90000000 | io_inAxi_ra_bits_addr < 32'h80000000) |
    io_inAxi_wa_valid & (io_inAxi_wa_bits_addr > 32'h90000000 | io_inAxi_wa_bits_addr < 32'h80000000)) &
    io_inAxi_rd_ready; // @[playground/src/sim/sim_crossbar.scala 25:289 27:26 playground/src/axi/axi.scala 87:18]
  wire  _GEN_32 = io_inAxi_ra_valid & (io_inAxi_ra_bits_addr > 32'h90000000 | io_inAxi_ra_bits_addr < 32'h80000000) |
    io_inAxi_wa_valid & (io_inAxi_wa_bits_addr > 32'h90000000 | io_inAxi_wa_bits_addr < 32'h80000000) ?
    io_mmioAxi_rd_valid : _GEN_2; // @[playground/src/sim/sim_crossbar.scala 25:289 27:26]
  wire [3:0] _GEN_33 = io_inAxi_ra_valid & (io_inAxi_ra_bits_addr > 32'h90000000 | io_inAxi_ra_bits_addr < 32'h80000000)
     | io_inAxi_wa_valid & (io_inAxi_wa_bits_addr > 32'h90000000 | io_inAxi_wa_bits_addr < 32'h80000000) ? 4'h0 : _GEN_3
    ; // @[playground/src/sim/sim_crossbar.scala 25:289 27:26]
  wire [63:0] _GEN_34 = io_inAxi_ra_valid & (io_inAxi_ra_bits_addr > 32'h90000000 | io_inAxi_ra_bits_addr < 32'h80000000
    ) | io_inAxi_wa_valid & (io_inAxi_wa_bits_addr > 32'h90000000 | io_inAxi_wa_bits_addr < 32'h80000000) ?
    io_mmioAxi_rd_bits_data : _GEN_4; // @[playground/src/sim/sim_crossbar.scala 25:289 27:26]
  wire [1:0] _GEN_35 = io_inAxi_ra_valid & (io_inAxi_ra_bits_addr > 32'h90000000 | io_inAxi_ra_bits_addr < 32'h80000000)
     | io_inAxi_wa_valid & (io_inAxi_wa_bits_addr > 32'h90000000 | io_inAxi_wa_bits_addr < 32'h80000000) ? 2'h0 : _GEN_5
    ; // @[playground/src/sim/sim_crossbar.scala 25:289 27:26]
  wire  _GEN_36 = io_inAxi_ra_valid & (io_inAxi_ra_bits_addr > 32'h90000000 | io_inAxi_ra_bits_addr < 32'h80000000) |
    io_inAxi_wa_valid & (io_inAxi_wa_bits_addr > 32'h90000000 | io_inAxi_wa_bits_addr < 32'h80000000) ?
    io_mmioAxi_rd_bits_last : _GEN_6; // @[playground/src/sim/sim_crossbar.scala 25:289 27:26]
  wire  _GEN_37 = io_inAxi_ra_valid & (io_inAxi_ra_bits_addr > 32'h90000000 | io_inAxi_ra_bits_addr < 32'h80000000) |
    io_inAxi_wa_valid & (io_inAxi_wa_bits_addr > 32'h90000000 | io_inAxi_wa_bits_addr < 32'h80000000) ?
    io_mmioAxi_ra_ready : _GEN_7; // @[playground/src/sim/sim_crossbar.scala 25:289 27:26]
  wire  _GEN_38 = (io_inAxi_ra_valid & (io_inAxi_ra_bits_addr > 32'h90000000 | io_inAxi_ra_bits_addr < 32'h80000000) |
    io_inAxi_wa_valid & (io_inAxi_wa_bits_addr > 32'h90000000 | io_inAxi_wa_bits_addr < 32'h80000000)) &
    io_inAxi_ra_valid; // @[playground/src/sim/sim_crossbar.scala 25:289 27:26 playground/src/axi/axi.scala 86:18]
  wire [31:0] _GEN_40 = io_inAxi_ra_valid & (io_inAxi_ra_bits_addr > 32'h90000000 | io_inAxi_ra_bits_addr < 32'h80000000
    ) | io_inAxi_wa_valid & (io_inAxi_wa_bits_addr > 32'h90000000 | io_inAxi_wa_bits_addr < 32'h80000000) ?
    io_inAxi_ra_bits_addr : 32'h0; // @[playground/src/sim/sim_crossbar.scala 25:289 27:26 playground/src/axi/axi.scala 41:23]
  wire  _GEN_45 = io_inAxi_ra_valid & (io_inAxi_ra_bits_addr > 32'h90000000 | io_inAxi_ra_bits_addr < 32'h80000000) |
    io_inAxi_wa_valid & (io_inAxi_wa_bits_addr > 32'h90000000 | io_inAxi_wa_bits_addr < 32'h80000000) | _GEN_15; // @[playground/src/sim/sim_crossbar.scala 25:289 27:26]
  wire [3:0] _GEN_46 = io_inAxi_ra_valid & (io_inAxi_ra_bits_addr > 32'h90000000 | io_inAxi_ra_bits_addr < 32'h80000000)
     | io_inAxi_wa_valid & (io_inAxi_wa_bits_addr > 32'h90000000 | io_inAxi_wa_bits_addr < 32'h80000000) ? 4'h0 :
    _GEN_16; // @[playground/src/sim/sim_crossbar.scala 25:289 27:26]
  wire [1:0] _GEN_47 = io_inAxi_ra_valid & (io_inAxi_ra_bits_addr > 32'h90000000 | io_inAxi_ra_bits_addr < 32'h80000000)
     | io_inAxi_wa_valid & (io_inAxi_wa_bits_addr > 32'h90000000 | io_inAxi_wa_bits_addr < 32'h80000000) ? 2'h0 :
    _GEN_17; // @[playground/src/sim/sim_crossbar.scala 25:289 27:26]
  wire  _GEN_48 = io_inAxi_ra_valid & (io_inAxi_ra_bits_addr > 32'h90000000 | io_inAxi_ra_bits_addr < 32'h80000000) |
    io_inAxi_wa_valid & (io_inAxi_wa_bits_addr > 32'h90000000 | io_inAxi_wa_bits_addr < 32'h80000000) ?
    io_mmioAxi_wd_ready : _GEN_18; // @[playground/src/sim/sim_crossbar.scala 25:289 27:26]
  wire  _GEN_49 = (io_inAxi_ra_valid & (io_inAxi_ra_bits_addr > 32'h90000000 | io_inAxi_ra_bits_addr < 32'h80000000) |
    io_inAxi_wa_valid & (io_inAxi_wa_bits_addr > 32'h90000000 | io_inAxi_wa_bits_addr < 32'h80000000)) &
    io_inAxi_wd_valid; // @[playground/src/sim/sim_crossbar.scala 25:289 27:26 playground/src/axi/axi.scala 84:18]
  wire [63:0] _GEN_50 = io_inAxi_ra_valid & (io_inAxi_ra_bits_addr > 32'h90000000 | io_inAxi_ra_bits_addr < 32'h80000000
    ) | io_inAxi_wa_valid & (io_inAxi_wa_bits_addr > 32'h90000000 | io_inAxi_wa_bits_addr < 32'h80000000) ?
    io_inAxi_wd_bits_data : 64'h0; // @[playground/src/sim/sim_crossbar.scala 25:289 27:26 playground/src/axi/axi.scala 50:23]
  wire [7:0] _GEN_51 = io_inAxi_ra_valid & (io_inAxi_ra_bits_addr > 32'h90000000 | io_inAxi_ra_bits_addr < 32'h80000000)
     | io_inAxi_wa_valid & (io_inAxi_wa_bits_addr > 32'h90000000 | io_inAxi_wa_bits_addr < 32'h80000000) ?
    io_inAxi_wd_bits_strb : 8'h0; // @[playground/src/sim/sim_crossbar.scala 25:289 27:26 playground/src/axi/axi.scala 50:23]
  wire  _GEN_52 = (io_inAxi_ra_valid & (io_inAxi_ra_bits_addr > 32'h90000000 | io_inAxi_ra_bits_addr < 32'h80000000) |
    io_inAxi_wa_valid & (io_inAxi_wa_bits_addr > 32'h90000000 | io_inAxi_wa_bits_addr < 32'h80000000)) &
    io_inAxi_wd_bits_last; // @[playground/src/sim/sim_crossbar.scala 25:289 27:26 playground/src/axi/axi.scala 50:23]
  wire  _GEN_53 = io_inAxi_ra_valid & (io_inAxi_ra_bits_addr > 32'h90000000 | io_inAxi_ra_bits_addr < 32'h80000000) |
    io_inAxi_wa_valid & (io_inAxi_wa_bits_addr > 32'h90000000 | io_inAxi_wa_bits_addr < 32'h80000000) ?
    io_mmioAxi_wa_ready : _GEN_23; // @[playground/src/sim/sim_crossbar.scala 25:289 27:26]
  wire  _GEN_54 = (io_inAxi_ra_valid & (io_inAxi_ra_bits_addr > 32'h90000000 | io_inAxi_ra_bits_addr < 32'h80000000) |
    io_inAxi_wa_valid & (io_inAxi_wa_bits_addr > 32'h90000000 | io_inAxi_wa_bits_addr < 32'h80000000)) &
    io_inAxi_wa_valid; // @[playground/src/sim/sim_crossbar.scala 25:289 27:26 playground/src/axi/axi.scala 83:18]
  wire [31:0] _GEN_56 = io_inAxi_ra_valid & (io_inAxi_ra_bits_addr > 32'h90000000 | io_inAxi_ra_bits_addr < 32'h80000000
    ) | io_inAxi_wa_valid & (io_inAxi_wa_bits_addr > 32'h90000000 | io_inAxi_wa_bits_addr < 32'h80000000) ?
    io_inAxi_wa_bits_addr : 32'h0; // @[playground/src/sim/sim_crossbar.scala 25:289 27:26 playground/src/axi/axi.scala 41:23]
  wire  _GEN_60 = io_inAxi_ra_valid & (io_inAxi_ra_bits_addr > 32'h90000000 | io_inAxi_ra_bits_addr < 32'h80000000) |
    io_inAxi_wa_valid & (io_inAxi_wa_bits_addr > 32'h90000000 | io_inAxi_wa_bits_addr < 32'h80000000) ? 1'h0 : _GEN_1; // @[playground/src/sim/sim_crossbar.scala 25:289 playground/src/axi/axi.scala 87:18]
  wire  _GEN_61 = io_inAxi_ra_valid & (io_inAxi_ra_bits_addr > 32'h90000000 | io_inAxi_ra_bits_addr < 32'h80000000) |
    io_inAxi_wa_valid & (io_inAxi_wa_bits_addr > 32'h90000000 | io_inAxi_wa_bits_addr < 32'h80000000) ? 1'h0 : _GEN_8; // @[playground/src/sim/sim_crossbar.scala 25:289 playground/src/axi/axi.scala 86:18]
  wire [3:0] _GEN_62 = io_inAxi_ra_valid & (io_inAxi_ra_bits_addr > 32'h90000000 | io_inAxi_ra_bits_addr < 32'h80000000)
     | io_inAxi_wa_valid & (io_inAxi_wa_bits_addr > 32'h90000000 | io_inAxi_wa_bits_addr < 32'h80000000) ? 4'h0 : _GEN_9
    ; // @[playground/src/sim/sim_crossbar.scala 25:289 playground/src/axi/axi.scala 41:23]
  wire [31:0] _GEN_63 = io_inAxi_ra_valid & (io_inAxi_ra_bits_addr > 32'h90000000 | io_inAxi_ra_bits_addr < 32'h80000000
    ) | io_inAxi_wa_valid & (io_inAxi_wa_bits_addr > 32'h90000000 | io_inAxi_wa_bits_addr < 32'h80000000) ? 32'h0 :
    _GEN_10; // @[playground/src/sim/sim_crossbar.scala 25:289 playground/src/axi/axi.scala 41:23]
  wire [7:0] _GEN_64 = io_inAxi_ra_valid & (io_inAxi_ra_bits_addr > 32'h90000000 | io_inAxi_ra_bits_addr < 32'h80000000)
     | io_inAxi_wa_valid & (io_inAxi_wa_bits_addr > 32'h90000000 | io_inAxi_wa_bits_addr < 32'h80000000) ? 8'h0 :
    _GEN_11; // @[playground/src/sim/sim_crossbar.scala 25:289 playground/src/axi/axi.scala 41:23]
  wire [2:0] _GEN_65 = io_inAxi_ra_valid & (io_inAxi_ra_bits_addr > 32'h90000000 | io_inAxi_ra_bits_addr < 32'h80000000)
     | io_inAxi_wa_valid & (io_inAxi_wa_bits_addr > 32'h90000000 | io_inAxi_wa_bits_addr < 32'h80000000) ? 3'h0 :
    _GEN_12; // @[playground/src/sim/sim_crossbar.scala 25:289 playground/src/axi/axi.scala 41:23]
  wire [1:0] _GEN_66 = io_inAxi_ra_valid & (io_inAxi_ra_bits_addr > 32'h90000000 | io_inAxi_ra_bits_addr < 32'h80000000)
     | io_inAxi_wa_valid & (io_inAxi_wa_bits_addr > 32'h90000000 | io_inAxi_wa_bits_addr < 32'h80000000) ? 2'h0 :
    _GEN_13; // @[playground/src/sim/sim_crossbar.scala 25:289 playground/src/axi/axi.scala 41:23]
  wire  _GEN_67 = io_inAxi_ra_valid & (io_inAxi_ra_bits_addr > 32'h90000000 | io_inAxi_ra_bits_addr < 32'h80000000) |
    io_inAxi_wa_valid & (io_inAxi_wa_bits_addr > 32'h90000000 | io_inAxi_wa_bits_addr < 32'h80000000) ? 1'h0 : _GEN_14; // @[playground/src/sim/sim_crossbar.scala 25:289 playground/src/axi/axi.scala 85:18]
  wire  _GEN_68 = io_inAxi_ra_valid & (io_inAxi_ra_bits_addr > 32'h90000000 | io_inAxi_ra_bits_addr < 32'h80000000) |
    io_inAxi_wa_valid & (io_inAxi_wa_bits_addr > 32'h90000000 | io_inAxi_wa_bits_addr < 32'h80000000) ? 1'h0 : _GEN_19; // @[playground/src/sim/sim_crossbar.scala 25:289 playground/src/axi/axi.scala 84:18]
  wire [63:0] _GEN_69 = io_inAxi_ra_valid & (io_inAxi_ra_bits_addr > 32'h90000000 | io_inAxi_ra_bits_addr < 32'h80000000
    ) | io_inAxi_wa_valid & (io_inAxi_wa_bits_addr > 32'h90000000 | io_inAxi_wa_bits_addr < 32'h80000000) ? 64'h0 :
    _GEN_20; // @[playground/src/sim/sim_crossbar.scala 25:289 playground/src/axi/axi.scala 50:23]
  wire [7:0] _GEN_70 = io_inAxi_ra_valid & (io_inAxi_ra_bits_addr > 32'h90000000 | io_inAxi_ra_bits_addr < 32'h80000000)
     | io_inAxi_wa_valid & (io_inAxi_wa_bits_addr > 32'h90000000 | io_inAxi_wa_bits_addr < 32'h80000000) ? 8'h0 :
    _GEN_21; // @[playground/src/sim/sim_crossbar.scala 25:289 playground/src/axi/axi.scala 50:23]
  wire  _GEN_71 = io_inAxi_ra_valid & (io_inAxi_ra_bits_addr > 32'h90000000 | io_inAxi_ra_bits_addr < 32'h80000000) |
    io_inAxi_wa_valid & (io_inAxi_wa_bits_addr > 32'h90000000 | io_inAxi_wa_bits_addr < 32'h80000000) ? 1'h0 : _GEN_22; // @[playground/src/sim/sim_crossbar.scala 25:289 playground/src/axi/axi.scala 50:23]
  wire  _GEN_72 = io_inAxi_ra_valid & (io_inAxi_ra_bits_addr > 32'h90000000 | io_inAxi_ra_bits_addr < 32'h80000000) |
    io_inAxi_wa_valid & (io_inAxi_wa_bits_addr > 32'h90000000 | io_inAxi_wa_bits_addr < 32'h80000000) ? 1'h0 : _GEN_24; // @[playground/src/sim/sim_crossbar.scala 25:289 playground/src/axi/axi.scala 83:18]
  wire [3:0] _GEN_73 = io_inAxi_ra_valid & (io_inAxi_ra_bits_addr > 32'h90000000 | io_inAxi_ra_bits_addr < 32'h80000000)
     | io_inAxi_wa_valid & (io_inAxi_wa_bits_addr > 32'h90000000 | io_inAxi_wa_bits_addr < 32'h80000000) ? 4'h0 :
    _GEN_25; // @[playground/src/sim/sim_crossbar.scala 25:289 playground/src/axi/axi.scala 41:23]
  wire [31:0] _GEN_74 = io_inAxi_ra_valid & (io_inAxi_ra_bits_addr > 32'h90000000 | io_inAxi_ra_bits_addr < 32'h80000000
    ) | io_inAxi_wa_valid & (io_inAxi_wa_bits_addr > 32'h90000000 | io_inAxi_wa_bits_addr < 32'h80000000) ? 32'h0 :
    _GEN_26; // @[playground/src/sim/sim_crossbar.scala 25:289 playground/src/axi/axi.scala 41:23]
  wire [7:0] _GEN_75 = io_inAxi_ra_valid & (io_inAxi_ra_bits_addr > 32'h90000000 | io_inAxi_ra_bits_addr < 32'h80000000)
     | io_inAxi_wa_valid & (io_inAxi_wa_bits_addr > 32'h90000000 | io_inAxi_wa_bits_addr < 32'h80000000) ? 8'h0 :
    _GEN_27; // @[playground/src/sim/sim_crossbar.scala 25:289 playground/src/axi/axi.scala 41:23]
  wire [2:0] _GEN_76 = io_inAxi_ra_valid & (io_inAxi_ra_bits_addr > 32'h90000000 | io_inAxi_ra_bits_addr < 32'h80000000)
     | io_inAxi_wa_valid & (io_inAxi_wa_bits_addr > 32'h90000000 | io_inAxi_wa_bits_addr < 32'h80000000) ? 3'h0 :
    _GEN_28; // @[playground/src/sim/sim_crossbar.scala 25:289 playground/src/axi/axi.scala 41:23]
  wire [1:0] _GEN_77 = io_inAxi_ra_valid & (io_inAxi_ra_bits_addr > 32'h90000000 | io_inAxi_ra_bits_addr < 32'h80000000)
     | io_inAxi_wa_valid & (io_inAxi_wa_bits_addr > 32'h90000000 | io_inAxi_wa_bits_addr < 32'h80000000) ? 2'h0 :
    _GEN_29; // @[playground/src/sim/sim_crossbar.scala 25:289 playground/src/axi/axi.scala 41:23]
  wire [1:0] _GEN_79 = io_mmioAxi_rd_valid & io_mmioAxi_rd_bits_last | io_mmioAxi_wd_valid & io_mmioAxi_wd_bits_last ? 2'h0
     : state; // @[playground/src/sim/sim_crossbar.scala 41:119 42:23 19:24]
  wire  _GEN_80 = 2'h2 == state & io_inAxi_rd_ready; // @[playground/src/sim/sim_crossbar.scala 20:18 40:22 playground/src/axi/axi.scala 87:18]
  wire  _GEN_81 = 2'h2 == state & io_mmioAxi_rd_valid; // @[playground/src/axi/axi.scala 105:18 playground/src/sim/sim_crossbar.scala 20:18 40:22]
  wire [63:0] _GEN_83 = 2'h2 == state ? io_mmioAxi_rd_bits_data : 64'h0; // @[playground/src/sim/sim_crossbar.scala 20:18 40:22 playground/src/axi/axi.scala 68:23]
  wire  _GEN_85 = 2'h2 == state & io_mmioAxi_rd_bits_last; // @[playground/src/sim/sim_crossbar.scala 20:18 40:22 playground/src/axi/axi.scala 68:23]
  wire  _GEN_86 = 2'h2 == state & io_mmioAxi_ra_ready; // @[playground/src/axi/axi.scala 104:18 playground/src/sim/sim_crossbar.scala 20:18 40:22]
  wire  _GEN_87 = 2'h2 == state & io_inAxi_ra_valid; // @[playground/src/sim/sim_crossbar.scala 20:18 40:22 playground/src/axi/axi.scala 86:18]
  wire [31:0] _GEN_89 = 2'h2 == state ? io_inAxi_ra_bits_addr : 32'h0; // @[playground/src/sim/sim_crossbar.scala 20:18 40:22 playground/src/axi/axi.scala 41:23]
  wire  _GEN_97 = 2'h2 == state & io_mmioAxi_wd_ready; // @[playground/src/axi/axi.scala 102:18 playground/src/sim/sim_crossbar.scala 20:18 40:22]
  wire  _GEN_98 = 2'h2 == state & io_inAxi_wd_valid; // @[playground/src/sim/sim_crossbar.scala 20:18 40:22 playground/src/axi/axi.scala 84:18]
  wire [63:0] _GEN_99 = 2'h2 == state ? io_inAxi_wd_bits_data : 64'h0; // @[playground/src/sim/sim_crossbar.scala 20:18 40:22 playground/src/axi/axi.scala 50:23]
  wire [7:0] _GEN_100 = 2'h2 == state ? io_inAxi_wd_bits_strb : 8'h0; // @[playground/src/sim/sim_crossbar.scala 20:18 40:22 playground/src/axi/axi.scala 50:23]
  wire  _GEN_101 = 2'h2 == state & io_inAxi_wd_bits_last; // @[playground/src/sim/sim_crossbar.scala 20:18 40:22 playground/src/axi/axi.scala 50:23]
  wire  _GEN_102 = 2'h2 == state & io_mmioAxi_wa_ready; // @[playground/src/axi/axi.scala 101:18 playground/src/sim/sim_crossbar.scala 20:18 40:22]
  wire  _GEN_103 = 2'h2 == state & io_inAxi_wa_valid; // @[playground/src/sim/sim_crossbar.scala 20:18 40:22 playground/src/axi/axi.scala 83:18]
  wire [31:0] _GEN_105 = 2'h2 == state ? io_inAxi_wa_bits_addr : 32'h0; // @[playground/src/sim/sim_crossbar.scala 20:18 40:22 playground/src/axi/axi.scala 41:23]
  wire  _GEN_110 = 2'h1 == state & io_inAxi_rd_ready; // @[playground/src/sim/sim_crossbar.scala 20:18 34:22 playground/src/axi/axi.scala 87:18]
  wire  _GEN_111 = 2'h1 == state ? io_memAxi_rd_valid : _GEN_81; // @[playground/src/sim/sim_crossbar.scala 20:18 34:22]
  wire [3:0] _GEN_112 = 2'h1 == state ? io_memAxi_rd_bits_id : 4'h0; // @[playground/src/sim/sim_crossbar.scala 20:18 34:22]
  wire [63:0] _GEN_113 = 2'h1 == state ? io_memAxi_rd_bits_data : _GEN_83; // @[playground/src/sim/sim_crossbar.scala 20:18 34:22]
  wire [1:0] _GEN_114 = 2'h1 == state ? io_memAxi_rd_bits_resp : 2'h0; // @[playground/src/sim/sim_crossbar.scala 20:18 34:22]
  wire  _GEN_115 = 2'h1 == state ? io_memAxi_rd_bits_last : _GEN_85; // @[playground/src/sim/sim_crossbar.scala 20:18 34:22]
  wire  _GEN_116 = 2'h1 == state ? io_memAxi_ra_ready : _GEN_86; // @[playground/src/sim/sim_crossbar.scala 20:18 34:22]
  wire  _GEN_117 = 2'h1 == state & io_inAxi_ra_valid; // @[playground/src/sim/sim_crossbar.scala 20:18 34:22 playground/src/axi/axi.scala 86:18]
  wire [3:0] _GEN_118 = 2'h1 == state ? io_inAxi_ra_bits_id : 4'h0; // @[playground/src/sim/sim_crossbar.scala 20:18 34:22 playground/src/axi/axi.scala 41:23]
  wire [31:0] _GEN_119 = 2'h1 == state ? io_inAxi_ra_bits_addr : 32'h0; // @[playground/src/sim/sim_crossbar.scala 20:18 34:22 playground/src/axi/axi.scala 41:23]
  wire [7:0] _GEN_120 = 2'h1 == state ? io_inAxi_ra_bits_len : 8'h0; // @[playground/src/sim/sim_crossbar.scala 20:18 34:22 playground/src/axi/axi.scala 41:23]
  wire [2:0] _GEN_121 = 2'h1 == state ? io_inAxi_ra_bits_size : 3'h0; // @[playground/src/sim/sim_crossbar.scala 20:18 34:22 playground/src/axi/axi.scala 41:23]
  wire [1:0] _GEN_122 = 2'h1 == state ? io_inAxi_ra_bits_burst : 2'h0; // @[playground/src/sim/sim_crossbar.scala 20:18 34:22 playground/src/axi/axi.scala 41:23]
  wire  _GEN_123 = 2'h1 == state & io_inAxi_wr_ready; // @[playground/src/sim/sim_crossbar.scala 20:18 34:22 playground/src/axi/axi.scala 85:18]
  wire  _GEN_124 = 2'h1 == state ? io_memAxi_wr_valid : 2'h2 == state; // @[playground/src/sim/sim_crossbar.scala 20:18 34:22]
  wire [3:0] _GEN_125 = 2'h1 == state ? io_memAxi_wr_bits_id : 4'h0; // @[playground/src/sim/sim_crossbar.scala 20:18 34:22]
  wire [1:0] _GEN_126 = 2'h1 == state ? io_memAxi_wr_bits_resp : 2'h0; // @[playground/src/sim/sim_crossbar.scala 20:18 34:22]
  wire  _GEN_127 = 2'h1 == state ? io_memAxi_wd_ready : _GEN_97; // @[playground/src/sim/sim_crossbar.scala 20:18 34:22]
  wire  _GEN_128 = 2'h1 == state & io_inAxi_wd_valid; // @[playground/src/sim/sim_crossbar.scala 20:18 34:22 playground/src/axi/axi.scala 84:18]
  wire [63:0] _GEN_129 = 2'h1 == state ? io_inAxi_wd_bits_data : 64'h0; // @[playground/src/sim/sim_crossbar.scala 20:18 34:22 playground/src/axi/axi.scala 50:23]
  wire [7:0] _GEN_130 = 2'h1 == state ? io_inAxi_wd_bits_strb : 8'h0; // @[playground/src/sim/sim_crossbar.scala 20:18 34:22 playground/src/axi/axi.scala 50:23]
  wire  _GEN_131 = 2'h1 == state & io_inAxi_wd_bits_last; // @[playground/src/sim/sim_crossbar.scala 20:18 34:22 playground/src/axi/axi.scala 50:23]
  wire  _GEN_132 = 2'h1 == state ? io_memAxi_wa_ready : _GEN_102; // @[playground/src/sim/sim_crossbar.scala 20:18 34:22]
  wire  _GEN_133 = 2'h1 == state & io_inAxi_wa_valid; // @[playground/src/sim/sim_crossbar.scala 20:18 34:22 playground/src/axi/axi.scala 83:18]
  wire [3:0] _GEN_134 = 2'h1 == state ? io_inAxi_wa_bits_id : 4'h0; // @[playground/src/sim/sim_crossbar.scala 20:18 34:22 playground/src/axi/axi.scala 41:23]
  wire [31:0] _GEN_135 = 2'h1 == state ? io_inAxi_wa_bits_addr : 32'h0; // @[playground/src/sim/sim_crossbar.scala 20:18 34:22 playground/src/axi/axi.scala 41:23]
  wire [7:0] _GEN_136 = 2'h1 == state ? io_inAxi_wa_bits_len : 8'h0; // @[playground/src/sim/sim_crossbar.scala 20:18 34:22 playground/src/axi/axi.scala 41:23]
  wire [2:0] _GEN_137 = 2'h1 == state ? io_inAxi_wa_bits_size : 3'h0; // @[playground/src/sim/sim_crossbar.scala 20:18 34:22 playground/src/axi/axi.scala 41:23]
  wire [1:0] _GEN_138 = 2'h1 == state ? io_inAxi_wa_bits_burst : 2'h0; // @[playground/src/sim/sim_crossbar.scala 20:18 34:22 playground/src/axi/axi.scala 41:23]
  wire  _GEN_140 = 2'h1 == state ? 1'h0 : _GEN_80; // @[playground/src/sim/sim_crossbar.scala 20:18 playground/src/axi/axi.scala 87:18]
  wire  _GEN_141 = 2'h1 == state ? 1'h0 : _GEN_87; // @[playground/src/sim/sim_crossbar.scala 20:18 playground/src/axi/axi.scala 86:18]
  wire [31:0] _GEN_143 = 2'h1 == state ? 32'h0 : _GEN_89; // @[playground/src/sim/sim_crossbar.scala 20:18 playground/src/axi/axi.scala 41:23]
  wire  _GEN_148 = 2'h1 == state ? 1'h0 : _GEN_98; // @[playground/src/sim/sim_crossbar.scala 20:18 playground/src/axi/axi.scala 84:18]
  wire [63:0] _GEN_149 = 2'h1 == state ? 64'h0 : _GEN_99; // @[playground/src/sim/sim_crossbar.scala 20:18 playground/src/axi/axi.scala 50:23]
  wire [7:0] _GEN_150 = 2'h1 == state ? 8'h0 : _GEN_100; // @[playground/src/sim/sim_crossbar.scala 20:18 playground/src/axi/axi.scala 50:23]
  wire  _GEN_151 = 2'h1 == state ? 1'h0 : _GEN_101; // @[playground/src/sim/sim_crossbar.scala 20:18 playground/src/axi/axi.scala 50:23]
  wire  _GEN_152 = 2'h1 == state ? 1'h0 : _GEN_103; // @[playground/src/sim/sim_crossbar.scala 20:18 playground/src/axi/axi.scala 83:18]
  wire [31:0] _GEN_154 = 2'h1 == state ? 32'h0 : _GEN_105; // @[playground/src/sim/sim_crossbar.scala 20:18 playground/src/axi/axi.scala 41:23]
  assign io_inAxi_wa_ready = 2'h0 == state ? _GEN_53 : _GEN_132; // @[playground/src/sim/sim_crossbar.scala 20:18]
  assign io_inAxi_wd_ready = 2'h0 == state ? _GEN_48 : _GEN_127; // @[playground/src/sim/sim_crossbar.scala 20:18]
  assign io_inAxi_wr_valid = 2'h0 == state ? _GEN_45 : _GEN_124; // @[playground/src/sim/sim_crossbar.scala 20:18]
  assign io_inAxi_wr_bits_id = 2'h0 == state ? _GEN_46 : _GEN_125; // @[playground/src/sim/sim_crossbar.scala 20:18]
  assign io_inAxi_wr_bits_resp = 2'h0 == state ? _GEN_47 : _GEN_126; // @[playground/src/sim/sim_crossbar.scala 20:18]
  assign io_inAxi_ra_ready = 2'h0 == state ? _GEN_37 : _GEN_116; // @[playground/src/sim/sim_crossbar.scala 20:18]
  assign io_inAxi_rd_valid = 2'h0 == state ? _GEN_32 : _GEN_111; // @[playground/src/sim/sim_crossbar.scala 20:18]
  assign io_inAxi_rd_bits_id = 2'h0 == state ? _GEN_33 : _GEN_112; // @[playground/src/sim/sim_crossbar.scala 20:18]
  assign io_inAxi_rd_bits_data = 2'h0 == state ? _GEN_34 : _GEN_113; // @[playground/src/sim/sim_crossbar.scala 20:18]
  assign io_inAxi_rd_bits_resp = 2'h0 == state ? _GEN_35 : _GEN_114; // @[playground/src/sim/sim_crossbar.scala 20:18]
  assign io_inAxi_rd_bits_last = 2'h0 == state ? _GEN_36 : _GEN_115; // @[playground/src/sim/sim_crossbar.scala 20:18]
  assign io_memAxi_wa_valid = 2'h0 == state ? _GEN_72 : _GEN_133; // @[playground/src/sim/sim_crossbar.scala 20:18]
  assign io_memAxi_wa_bits_id = 2'h0 == state ? _GEN_73 : _GEN_134; // @[playground/src/sim/sim_crossbar.scala 20:18]
  assign io_memAxi_wa_bits_addr = 2'h0 == state ? _GEN_74 : _GEN_135; // @[playground/src/sim/sim_crossbar.scala 20:18]
  assign io_memAxi_wa_bits_len = 2'h0 == state ? _GEN_75 : _GEN_136; // @[playground/src/sim/sim_crossbar.scala 20:18]
  assign io_memAxi_wa_bits_size = 2'h0 == state ? _GEN_76 : _GEN_137; // @[playground/src/sim/sim_crossbar.scala 20:18]
  assign io_memAxi_wa_bits_burst = 2'h0 == state ? _GEN_77 : _GEN_138; // @[playground/src/sim/sim_crossbar.scala 20:18]
  assign io_memAxi_wd_valid = 2'h0 == state ? _GEN_68 : _GEN_128; // @[playground/src/sim/sim_crossbar.scala 20:18]
  assign io_memAxi_wd_bits_data = 2'h0 == state ? _GEN_69 : _GEN_129; // @[playground/src/sim/sim_crossbar.scala 20:18]
  assign io_memAxi_wd_bits_strb = 2'h0 == state ? _GEN_70 : _GEN_130; // @[playground/src/sim/sim_crossbar.scala 20:18]
  assign io_memAxi_wd_bits_last = 2'h0 == state ? _GEN_71 : _GEN_131; // @[playground/src/sim/sim_crossbar.scala 20:18]
  assign io_memAxi_wr_ready = 2'h0 == state ? _GEN_67 : _GEN_123; // @[playground/src/sim/sim_crossbar.scala 20:18]
  assign io_memAxi_ra_valid = 2'h0 == state ? _GEN_61 : _GEN_117; // @[playground/src/sim/sim_crossbar.scala 20:18]
  assign io_memAxi_ra_bits_id = 2'h0 == state ? _GEN_62 : _GEN_118; // @[playground/src/sim/sim_crossbar.scala 20:18]
  assign io_memAxi_ra_bits_addr = 2'h0 == state ? _GEN_63 : _GEN_119; // @[playground/src/sim/sim_crossbar.scala 20:18]
  assign io_memAxi_ra_bits_len = 2'h0 == state ? _GEN_64 : _GEN_120; // @[playground/src/sim/sim_crossbar.scala 20:18]
  assign io_memAxi_ra_bits_size = 2'h0 == state ? _GEN_65 : _GEN_121; // @[playground/src/sim/sim_crossbar.scala 20:18]
  assign io_memAxi_ra_bits_burst = 2'h0 == state ? _GEN_66 : _GEN_122; // @[playground/src/sim/sim_crossbar.scala 20:18]
  assign io_memAxi_rd_ready = 2'h0 == state ? _GEN_60 : _GEN_110; // @[playground/src/sim/sim_crossbar.scala 20:18]
  assign io_mmioAxi_wa_valid = 2'h0 == state ? _GEN_54 : _GEN_152; // @[playground/src/sim/sim_crossbar.scala 20:18]
  assign io_mmioAxi_wa_bits_addr = 2'h0 == state ? _GEN_56 : _GEN_154; // @[playground/src/sim/sim_crossbar.scala 20:18]
  assign io_mmioAxi_wd_valid = 2'h0 == state ? _GEN_49 : _GEN_148; // @[playground/src/sim/sim_crossbar.scala 20:18]
  assign io_mmioAxi_wd_bits_data = 2'h0 == state ? _GEN_50 : _GEN_149; // @[playground/src/sim/sim_crossbar.scala 20:18]
  assign io_mmioAxi_wd_bits_strb = 2'h0 == state ? _GEN_51 : _GEN_150; // @[playground/src/sim/sim_crossbar.scala 20:18]
  assign io_mmioAxi_wd_bits_last = 2'h0 == state ? _GEN_52 : _GEN_151; // @[playground/src/sim/sim_crossbar.scala 20:18]
  assign io_mmioAxi_ra_valid = 2'h0 == state ? _GEN_38 : _GEN_141; // @[playground/src/sim/sim_crossbar.scala 20:18]
  assign io_mmioAxi_ra_bits_addr = 2'h0 == state ? _GEN_40 : _GEN_143; // @[playground/src/sim/sim_crossbar.scala 20:18]
  assign io_mmioAxi_rd_ready = 2'h0 == state ? _GEN_31 : _GEN_140; // @[playground/src/sim/sim_crossbar.scala 20:18]
  always @(posedge clock) begin
    if (reset) begin // @[playground/src/sim/sim_crossbar.scala 19:24]
      state <= 2'h0; // @[playground/src/sim/sim_crossbar.scala 19:24]
    end else if (2'h0 == state) begin // @[playground/src/sim/sim_crossbar.scala 20:18]
      if (io_inAxi_ra_valid & (io_inAxi_ra_bits_addr > 32'h90000000 | io_inAxi_ra_bits_addr < 32'h80000000) |
        io_inAxi_wa_valid & (io_inAxi_wa_bits_addr > 32'h90000000 | io_inAxi_wa_bits_addr < 32'h80000000)) begin // @[playground/src/sim/sim_crossbar.scala 25:289]
        state <= 2'h2; // @[playground/src/sim/sim_crossbar.scala 26:23]
      end else if (io_inAxi_ra_valid | io_inAxi_wa_valid) begin // @[playground/src/sim/sim_crossbar.scala 28:63]
        state <= 2'h1; // @[playground/src/sim/sim_crossbar.scala 29:23]
      end
    end else if (2'h1 == state) begin // @[playground/src/sim/sim_crossbar.scala 20:18]
      if (io_memAxi_rd_valid & io_memAxi_rd_bits_last | io_memAxi_wd_valid & io_memAxi_wd_bits_last) begin // @[playground/src/sim/sim_crossbar.scala 35:115]
        state <= 2'h0; // @[playground/src/sim/sim_crossbar.scala 36:23]
      end
    end else if (2'h2 == state) begin // @[playground/src/sim/sim_crossbar.scala 20:18]
      state <= _GEN_79;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TransAXI(
  output        io_raw_axi_awready, // @[playground/src/sim/bus.scala 10:16]
  input         io_raw_axi_awvalid, // @[playground/src/sim/bus.scala 10:16]
  input  [31:0] io_raw_axi_awaddr, // @[playground/src/sim/bus.scala 10:16]
  input  [3:0]  io_raw_axi_awid, // @[playground/src/sim/bus.scala 10:16]
  input  [7:0]  io_raw_axi_awlen, // @[playground/src/sim/bus.scala 10:16]
  input  [2:0]  io_raw_axi_awsize, // @[playground/src/sim/bus.scala 10:16]
  input  [1:0]  io_raw_axi_awburst, // @[playground/src/sim/bus.scala 10:16]
  output        io_raw_axi_wready, // @[playground/src/sim/bus.scala 10:16]
  input         io_raw_axi_wvalid, // @[playground/src/sim/bus.scala 10:16]
  input  [63:0] io_raw_axi_wdata, // @[playground/src/sim/bus.scala 10:16]
  input  [7:0]  io_raw_axi_wstrb, // @[playground/src/sim/bus.scala 10:16]
  input         io_raw_axi_wlast, // @[playground/src/sim/bus.scala 10:16]
  input         io_raw_axi_bready, // @[playground/src/sim/bus.scala 10:16]
  output        io_raw_axi_bvalid, // @[playground/src/sim/bus.scala 10:16]
  output [1:0]  io_raw_axi_bresp, // @[playground/src/sim/bus.scala 10:16]
  output [3:0]  io_raw_axi_bid, // @[playground/src/sim/bus.scala 10:16]
  output        io_raw_axi_arready, // @[playground/src/sim/bus.scala 10:16]
  input         io_raw_axi_arvalid, // @[playground/src/sim/bus.scala 10:16]
  input  [31:0] io_raw_axi_araddr, // @[playground/src/sim/bus.scala 10:16]
  input  [3:0]  io_raw_axi_arid, // @[playground/src/sim/bus.scala 10:16]
  input  [7:0]  io_raw_axi_arlen, // @[playground/src/sim/bus.scala 10:16]
  input  [2:0]  io_raw_axi_arsize, // @[playground/src/sim/bus.scala 10:16]
  input  [1:0]  io_raw_axi_arburst, // @[playground/src/sim/bus.scala 10:16]
  input         io_raw_axi_rready, // @[playground/src/sim/bus.scala 10:16]
  output        io_raw_axi_rvalid, // @[playground/src/sim/bus.scala 10:16]
  output [1:0]  io_raw_axi_rresp, // @[playground/src/sim/bus.scala 10:16]
  output [63:0] io_raw_axi_rdata, // @[playground/src/sim/bus.scala 10:16]
  output        io_raw_axi_rlast, // @[playground/src/sim/bus.scala 10:16]
  output [3:0]  io_raw_axi_rid, // @[playground/src/sim/bus.scala 10:16]
  input         io_bun_axi_wa_ready, // @[playground/src/sim/bus.scala 10:16]
  output        io_bun_axi_wa_valid, // @[playground/src/sim/bus.scala 10:16]
  output [3:0]  io_bun_axi_wa_bits_id, // @[playground/src/sim/bus.scala 10:16]
  output [31:0] io_bun_axi_wa_bits_addr, // @[playground/src/sim/bus.scala 10:16]
  output [7:0]  io_bun_axi_wa_bits_len, // @[playground/src/sim/bus.scala 10:16]
  output [2:0]  io_bun_axi_wa_bits_size, // @[playground/src/sim/bus.scala 10:16]
  output [1:0]  io_bun_axi_wa_bits_burst, // @[playground/src/sim/bus.scala 10:16]
  input         io_bun_axi_wd_ready, // @[playground/src/sim/bus.scala 10:16]
  output        io_bun_axi_wd_valid, // @[playground/src/sim/bus.scala 10:16]
  output [63:0] io_bun_axi_wd_bits_data, // @[playground/src/sim/bus.scala 10:16]
  output [7:0]  io_bun_axi_wd_bits_strb, // @[playground/src/sim/bus.scala 10:16]
  output        io_bun_axi_wd_bits_last, // @[playground/src/sim/bus.scala 10:16]
  output        io_bun_axi_wr_ready, // @[playground/src/sim/bus.scala 10:16]
  input         io_bun_axi_wr_valid, // @[playground/src/sim/bus.scala 10:16]
  input  [3:0]  io_bun_axi_wr_bits_id, // @[playground/src/sim/bus.scala 10:16]
  input  [1:0]  io_bun_axi_wr_bits_resp, // @[playground/src/sim/bus.scala 10:16]
  input         io_bun_axi_ra_ready, // @[playground/src/sim/bus.scala 10:16]
  output        io_bun_axi_ra_valid, // @[playground/src/sim/bus.scala 10:16]
  output [3:0]  io_bun_axi_ra_bits_id, // @[playground/src/sim/bus.scala 10:16]
  output [31:0] io_bun_axi_ra_bits_addr, // @[playground/src/sim/bus.scala 10:16]
  output [7:0]  io_bun_axi_ra_bits_len, // @[playground/src/sim/bus.scala 10:16]
  output [2:0]  io_bun_axi_ra_bits_size, // @[playground/src/sim/bus.scala 10:16]
  output [1:0]  io_bun_axi_ra_bits_burst, // @[playground/src/sim/bus.scala 10:16]
  output        io_bun_axi_rd_ready, // @[playground/src/sim/bus.scala 10:16]
  input         io_bun_axi_rd_valid, // @[playground/src/sim/bus.scala 10:16]
  input  [3:0]  io_bun_axi_rd_bits_id, // @[playground/src/sim/bus.scala 10:16]
  input  [63:0] io_bun_axi_rd_bits_data, // @[playground/src/sim/bus.scala 10:16]
  input  [1:0]  io_bun_axi_rd_bits_resp, // @[playground/src/sim/bus.scala 10:16]
  input         io_bun_axi_rd_bits_last // @[playground/src/sim/bus.scala 10:16]
);
  assign io_raw_axi_awready = io_bun_axi_wa_ready; // @[playground/src/sim/bus.scala 16:30]
  assign io_raw_axi_wready = io_bun_axi_wd_ready; // @[playground/src/sim/bus.scala 24:30]
  assign io_raw_axi_bvalid = io_bun_axi_wr_valid; // @[playground/src/sim/bus.scala 31:30]
  assign io_raw_axi_bresp = io_bun_axi_wr_bits_resp; // @[playground/src/sim/bus.scala 32:30]
  assign io_raw_axi_bid = io_bun_axi_wr_bits_id; // @[playground/src/sim/bus.scala 33:30]
  assign io_raw_axi_arready = io_bun_axi_ra_ready; // @[playground/src/sim/bus.scala 35:30]
  assign io_raw_axi_rvalid = io_bun_axi_rd_valid; // @[playground/src/sim/bus.scala 44:30]
  assign io_raw_axi_rresp = io_bun_axi_rd_bits_resp; // @[playground/src/sim/bus.scala 45:30]
  assign io_raw_axi_rdata = io_bun_axi_rd_bits_data; // @[playground/src/sim/bus.scala 46:30]
  assign io_raw_axi_rlast = io_bun_axi_rd_bits_last; // @[playground/src/sim/bus.scala 47:30]
  assign io_raw_axi_rid = io_bun_axi_rd_bits_id; // @[playground/src/sim/bus.scala 48:30]
  assign io_bun_axi_wa_valid = io_raw_axi_awvalid; // @[playground/src/sim/bus.scala 17:30]
  assign io_bun_axi_wa_bits_id = io_raw_axi_awid; // @[playground/src/sim/bus.scala 19:30]
  assign io_bun_axi_wa_bits_addr = io_raw_axi_awaddr; // @[playground/src/sim/bus.scala 18:30]
  assign io_bun_axi_wa_bits_len = io_raw_axi_awlen; // @[playground/src/sim/bus.scala 20:30]
  assign io_bun_axi_wa_bits_size = io_raw_axi_awsize; // @[playground/src/sim/bus.scala 21:30]
  assign io_bun_axi_wa_bits_burst = io_raw_axi_awburst; // @[playground/src/sim/bus.scala 22:30]
  assign io_bun_axi_wd_valid = io_raw_axi_wvalid; // @[playground/src/sim/bus.scala 25:30]
  assign io_bun_axi_wd_bits_data = io_raw_axi_wdata; // @[playground/src/sim/bus.scala 26:30]
  assign io_bun_axi_wd_bits_strb = io_raw_axi_wstrb; // @[playground/src/sim/bus.scala 27:30]
  assign io_bun_axi_wd_bits_last = io_raw_axi_wlast; // @[playground/src/sim/bus.scala 28:30]
  assign io_bun_axi_wr_ready = io_raw_axi_bready; // @[playground/src/sim/bus.scala 30:30]
  assign io_bun_axi_ra_valid = io_raw_axi_arvalid; // @[playground/src/sim/bus.scala 36:30]
  assign io_bun_axi_ra_bits_id = io_raw_axi_arid; // @[playground/src/sim/bus.scala 38:30]
  assign io_bun_axi_ra_bits_addr = io_raw_axi_araddr; // @[playground/src/sim/bus.scala 37:30]
  assign io_bun_axi_ra_bits_len = io_raw_axi_arlen; // @[playground/src/sim/bus.scala 39:30]
  assign io_bun_axi_ra_bits_size = io_raw_axi_arsize; // @[playground/src/sim/bus.scala 40:30]
  assign io_bun_axi_ra_bits_burst = io_raw_axi_arburst; // @[playground/src/sim/bus.scala 41:30]
  assign io_bun_axi_rd_ready = io_raw_axi_rready; // @[playground/src/sim/bus.scala 43:30]
endmodule
module newtop(
  input   clock,
  input   reset
);
  wire  cpu_clock; // @[playground/src/sim/sim_core.scala 17:21]
  wire  cpu_reset; // @[playground/src/sim/sim_core.scala 17:21]
  wire  cpu_io_master_awready; // @[playground/src/sim/sim_core.scala 17:21]
  wire  cpu_io_master_awvalid; // @[playground/src/sim/sim_core.scala 17:21]
  wire [31:0] cpu_io_master_awaddr; // @[playground/src/sim/sim_core.scala 17:21]
  wire [3:0] cpu_io_master_awid; // @[playground/src/sim/sim_core.scala 17:21]
  wire [7:0] cpu_io_master_awlen; // @[playground/src/sim/sim_core.scala 17:21]
  wire [2:0] cpu_io_master_awsize; // @[playground/src/sim/sim_core.scala 17:21]
  wire [1:0] cpu_io_master_awburst; // @[playground/src/sim/sim_core.scala 17:21]
  wire  cpu_io_master_wready; // @[playground/src/sim/sim_core.scala 17:21]
  wire  cpu_io_master_wvalid; // @[playground/src/sim/sim_core.scala 17:21]
  wire [63:0] cpu_io_master_wdata; // @[playground/src/sim/sim_core.scala 17:21]
  wire [7:0] cpu_io_master_wstrb; // @[playground/src/sim/sim_core.scala 17:21]
  wire  cpu_io_master_wlast; // @[playground/src/sim/sim_core.scala 17:21]
  wire  cpu_io_master_bready; // @[playground/src/sim/sim_core.scala 17:21]
  wire  cpu_io_master_bvalid; // @[playground/src/sim/sim_core.scala 17:21]
  wire [1:0] cpu_io_master_bresp; // @[playground/src/sim/sim_core.scala 17:21]
  wire [3:0] cpu_io_master_bid; // @[playground/src/sim/sim_core.scala 17:21]
  wire  cpu_io_master_arready; // @[playground/src/sim/sim_core.scala 17:21]
  wire  cpu_io_master_arvalid; // @[playground/src/sim/sim_core.scala 17:21]
  wire [31:0] cpu_io_master_araddr; // @[playground/src/sim/sim_core.scala 17:21]
  wire [3:0] cpu_io_master_arid; // @[playground/src/sim/sim_core.scala 17:21]
  wire [7:0] cpu_io_master_arlen; // @[playground/src/sim/sim_core.scala 17:21]
  wire [2:0] cpu_io_master_arsize; // @[playground/src/sim/sim_core.scala 17:21]
  wire [1:0] cpu_io_master_arburst; // @[playground/src/sim/sim_core.scala 17:21]
  wire  cpu_io_master_rready; // @[playground/src/sim/sim_core.scala 17:21]
  wire  cpu_io_master_rvalid; // @[playground/src/sim/sim_core.scala 17:21]
  wire [1:0] cpu_io_master_rresp; // @[playground/src/sim/sim_core.scala 17:21]
  wire [63:0] cpu_io_master_rdata; // @[playground/src/sim/sim_core.scala 17:21]
  wire  cpu_io_master_rlast; // @[playground/src/sim/sim_core.scala 17:21]
  wire [3:0] cpu_io_master_rid; // @[playground/src/sim/sim_core.scala 17:21]
  wire  cpu_io_slave_awready; // @[playground/src/sim/sim_core.scala 17:21]
  wire  cpu_io_slave_awvalid; // @[playground/src/sim/sim_core.scala 17:21]
  wire [31:0] cpu_io_slave_awaddr; // @[playground/src/sim/sim_core.scala 17:21]
  wire [3:0] cpu_io_slave_awid; // @[playground/src/sim/sim_core.scala 17:21]
  wire [7:0] cpu_io_slave_awlen; // @[playground/src/sim/sim_core.scala 17:21]
  wire [2:0] cpu_io_slave_awsize; // @[playground/src/sim/sim_core.scala 17:21]
  wire [1:0] cpu_io_slave_awburst; // @[playground/src/sim/sim_core.scala 17:21]
  wire  cpu_io_slave_wready; // @[playground/src/sim/sim_core.scala 17:21]
  wire  cpu_io_slave_wvalid; // @[playground/src/sim/sim_core.scala 17:21]
  wire [63:0] cpu_io_slave_wdata; // @[playground/src/sim/sim_core.scala 17:21]
  wire [7:0] cpu_io_slave_wstrb; // @[playground/src/sim/sim_core.scala 17:21]
  wire  cpu_io_slave_wlast; // @[playground/src/sim/sim_core.scala 17:21]
  wire  cpu_io_slave_bready; // @[playground/src/sim/sim_core.scala 17:21]
  wire  cpu_io_slave_bvalid; // @[playground/src/sim/sim_core.scala 17:21]
  wire [1:0] cpu_io_slave_bresp; // @[playground/src/sim/sim_core.scala 17:21]
  wire [3:0] cpu_io_slave_bid; // @[playground/src/sim/sim_core.scala 17:21]
  wire  cpu_io_slave_arready; // @[playground/src/sim/sim_core.scala 17:21]
  wire  cpu_io_slave_arvalid; // @[playground/src/sim/sim_core.scala 17:21]
  wire [31:0] cpu_io_slave_araddr; // @[playground/src/sim/sim_core.scala 17:21]
  wire [3:0] cpu_io_slave_arid; // @[playground/src/sim/sim_core.scala 17:21]
  wire [7:0] cpu_io_slave_arlen; // @[playground/src/sim/sim_core.scala 17:21]
  wire [2:0] cpu_io_slave_arsize; // @[playground/src/sim/sim_core.scala 17:21]
  wire [1:0] cpu_io_slave_arburst; // @[playground/src/sim/sim_core.scala 17:21]
  wire  cpu_io_slave_rready; // @[playground/src/sim/sim_core.scala 17:21]
  wire  cpu_io_slave_rvalid; // @[playground/src/sim/sim_core.scala 17:21]
  wire [1:0] cpu_io_slave_rresp; // @[playground/src/sim/sim_core.scala 17:21]
  wire [63:0] cpu_io_slave_rdata; // @[playground/src/sim/sim_core.scala 17:21]
  wire  cpu_io_slave_rlast; // @[playground/src/sim/sim_core.scala 17:21]
  wire [3:0] cpu_io_slave_rid; // @[playground/src/sim/sim_core.scala 17:21]
  wire  cpu_io_interrupt; // @[playground/src/sim/sim_core.scala 17:21]
  wire  mem_clock; // @[playground/src/sim/sim_core.scala 18:21]
  wire  mem_reset; // @[playground/src/sim/sim_core.scala 18:21]
  wire  mem_io_memAxi_wa_ready; // @[playground/src/sim/sim_core.scala 18:21]
  wire  mem_io_memAxi_wa_valid; // @[playground/src/sim/sim_core.scala 18:21]
  wire [3:0] mem_io_memAxi_wa_bits_id; // @[playground/src/sim/sim_core.scala 18:21]
  wire [31:0] mem_io_memAxi_wa_bits_addr; // @[playground/src/sim/sim_core.scala 18:21]
  wire [7:0] mem_io_memAxi_wa_bits_len; // @[playground/src/sim/sim_core.scala 18:21]
  wire [2:0] mem_io_memAxi_wa_bits_size; // @[playground/src/sim/sim_core.scala 18:21]
  wire [1:0] mem_io_memAxi_wa_bits_burst; // @[playground/src/sim/sim_core.scala 18:21]
  wire  mem_io_memAxi_wd_ready; // @[playground/src/sim/sim_core.scala 18:21]
  wire  mem_io_memAxi_wd_valid; // @[playground/src/sim/sim_core.scala 18:21]
  wire [63:0] mem_io_memAxi_wd_bits_data; // @[playground/src/sim/sim_core.scala 18:21]
  wire [7:0] mem_io_memAxi_wd_bits_strb; // @[playground/src/sim/sim_core.scala 18:21]
  wire  mem_io_memAxi_wd_bits_last; // @[playground/src/sim/sim_core.scala 18:21]
  wire  mem_io_memAxi_wr_ready; // @[playground/src/sim/sim_core.scala 18:21]
  wire  mem_io_memAxi_wr_valid; // @[playground/src/sim/sim_core.scala 18:21]
  wire [3:0] mem_io_memAxi_wr_bits_id; // @[playground/src/sim/sim_core.scala 18:21]
  wire [1:0] mem_io_memAxi_wr_bits_resp; // @[playground/src/sim/sim_core.scala 18:21]
  wire  mem_io_memAxi_ra_ready; // @[playground/src/sim/sim_core.scala 18:21]
  wire  mem_io_memAxi_ra_valid; // @[playground/src/sim/sim_core.scala 18:21]
  wire [3:0] mem_io_memAxi_ra_bits_id; // @[playground/src/sim/sim_core.scala 18:21]
  wire [31:0] mem_io_memAxi_ra_bits_addr; // @[playground/src/sim/sim_core.scala 18:21]
  wire [7:0] mem_io_memAxi_ra_bits_len; // @[playground/src/sim/sim_core.scala 18:21]
  wire [2:0] mem_io_memAxi_ra_bits_size; // @[playground/src/sim/sim_core.scala 18:21]
  wire [1:0] mem_io_memAxi_ra_bits_burst; // @[playground/src/sim/sim_core.scala 18:21]
  wire  mem_io_memAxi_rd_ready; // @[playground/src/sim/sim_core.scala 18:21]
  wire  mem_io_memAxi_rd_valid; // @[playground/src/sim/sim_core.scala 18:21]
  wire [3:0] mem_io_memAxi_rd_bits_id; // @[playground/src/sim/sim_core.scala 18:21]
  wire [63:0] mem_io_memAxi_rd_bits_data; // @[playground/src/sim/sim_core.scala 18:21]
  wire [1:0] mem_io_memAxi_rd_bits_resp; // @[playground/src/sim/sim_core.scala 18:21]
  wire  mem_io_memAxi_rd_bits_last; // @[playground/src/sim/sim_core.scala 18:21]
  wire  mmio_clock; // @[playground/src/sim/sim_core.scala 19:22]
  wire  mmio_reset; // @[playground/src/sim/sim_core.scala 19:22]
  wire  mmio_io_mmioAxi_wa_ready; // @[playground/src/sim/sim_core.scala 19:22]
  wire  mmio_io_mmioAxi_wa_valid; // @[playground/src/sim/sim_core.scala 19:22]
  wire [31:0] mmio_io_mmioAxi_wa_bits_addr; // @[playground/src/sim/sim_core.scala 19:22]
  wire  mmio_io_mmioAxi_wd_ready; // @[playground/src/sim/sim_core.scala 19:22]
  wire  mmio_io_mmioAxi_wd_valid; // @[playground/src/sim/sim_core.scala 19:22]
  wire [63:0] mmio_io_mmioAxi_wd_bits_data; // @[playground/src/sim/sim_core.scala 19:22]
  wire [7:0] mmio_io_mmioAxi_wd_bits_strb; // @[playground/src/sim/sim_core.scala 19:22]
  wire  mmio_io_mmioAxi_wd_bits_last; // @[playground/src/sim/sim_core.scala 19:22]
  wire  mmio_io_mmioAxi_ra_ready; // @[playground/src/sim/sim_core.scala 19:22]
  wire  mmio_io_mmioAxi_ra_valid; // @[playground/src/sim/sim_core.scala 19:22]
  wire [31:0] mmio_io_mmioAxi_ra_bits_addr; // @[playground/src/sim/sim_core.scala 19:22]
  wire  mmio_io_mmioAxi_rd_ready; // @[playground/src/sim/sim_core.scala 19:22]
  wire  mmio_io_mmioAxi_rd_valid; // @[playground/src/sim/sim_core.scala 19:22]
  wire [63:0] mmio_io_mmioAxi_rd_bits_data; // @[playground/src/sim/sim_core.scala 19:22]
  wire  mmio_io_mmioAxi_rd_bits_last; // @[playground/src/sim/sim_core.scala 19:22]
  wire  dma_clock; // @[playground/src/sim/sim_core.scala 20:21]
  wire  dma_reset; // @[playground/src/sim/sim_core.scala 20:21]
  wire [7:0] dma_io_dmaAxi_wstrb; // @[playground/src/sim/sim_core.scala 20:21]
  wire  crossBar_clock; // @[playground/src/sim/sim_core.scala 21:26]
  wire  crossBar_reset; // @[playground/src/sim/sim_core.scala 21:26]
  wire  crossBar_io_inAxi_wa_ready; // @[playground/src/sim/sim_core.scala 21:26]
  wire  crossBar_io_inAxi_wa_valid; // @[playground/src/sim/sim_core.scala 21:26]
  wire [3:0] crossBar_io_inAxi_wa_bits_id; // @[playground/src/sim/sim_core.scala 21:26]
  wire [31:0] crossBar_io_inAxi_wa_bits_addr; // @[playground/src/sim/sim_core.scala 21:26]
  wire [7:0] crossBar_io_inAxi_wa_bits_len; // @[playground/src/sim/sim_core.scala 21:26]
  wire [2:0] crossBar_io_inAxi_wa_bits_size; // @[playground/src/sim/sim_core.scala 21:26]
  wire [1:0] crossBar_io_inAxi_wa_bits_burst; // @[playground/src/sim/sim_core.scala 21:26]
  wire  crossBar_io_inAxi_wd_ready; // @[playground/src/sim/sim_core.scala 21:26]
  wire  crossBar_io_inAxi_wd_valid; // @[playground/src/sim/sim_core.scala 21:26]
  wire [63:0] crossBar_io_inAxi_wd_bits_data; // @[playground/src/sim/sim_core.scala 21:26]
  wire [7:0] crossBar_io_inAxi_wd_bits_strb; // @[playground/src/sim/sim_core.scala 21:26]
  wire  crossBar_io_inAxi_wd_bits_last; // @[playground/src/sim/sim_core.scala 21:26]
  wire  crossBar_io_inAxi_wr_ready; // @[playground/src/sim/sim_core.scala 21:26]
  wire  crossBar_io_inAxi_wr_valid; // @[playground/src/sim/sim_core.scala 21:26]
  wire [3:0] crossBar_io_inAxi_wr_bits_id; // @[playground/src/sim/sim_core.scala 21:26]
  wire [1:0] crossBar_io_inAxi_wr_bits_resp; // @[playground/src/sim/sim_core.scala 21:26]
  wire  crossBar_io_inAxi_ra_ready; // @[playground/src/sim/sim_core.scala 21:26]
  wire  crossBar_io_inAxi_ra_valid; // @[playground/src/sim/sim_core.scala 21:26]
  wire [3:0] crossBar_io_inAxi_ra_bits_id; // @[playground/src/sim/sim_core.scala 21:26]
  wire [31:0] crossBar_io_inAxi_ra_bits_addr; // @[playground/src/sim/sim_core.scala 21:26]
  wire [7:0] crossBar_io_inAxi_ra_bits_len; // @[playground/src/sim/sim_core.scala 21:26]
  wire [2:0] crossBar_io_inAxi_ra_bits_size; // @[playground/src/sim/sim_core.scala 21:26]
  wire [1:0] crossBar_io_inAxi_ra_bits_burst; // @[playground/src/sim/sim_core.scala 21:26]
  wire  crossBar_io_inAxi_rd_ready; // @[playground/src/sim/sim_core.scala 21:26]
  wire  crossBar_io_inAxi_rd_valid; // @[playground/src/sim/sim_core.scala 21:26]
  wire [3:0] crossBar_io_inAxi_rd_bits_id; // @[playground/src/sim/sim_core.scala 21:26]
  wire [63:0] crossBar_io_inAxi_rd_bits_data; // @[playground/src/sim/sim_core.scala 21:26]
  wire [1:0] crossBar_io_inAxi_rd_bits_resp; // @[playground/src/sim/sim_core.scala 21:26]
  wire  crossBar_io_inAxi_rd_bits_last; // @[playground/src/sim/sim_core.scala 21:26]
  wire  crossBar_io_memAxi_wa_ready; // @[playground/src/sim/sim_core.scala 21:26]
  wire  crossBar_io_memAxi_wa_valid; // @[playground/src/sim/sim_core.scala 21:26]
  wire [3:0] crossBar_io_memAxi_wa_bits_id; // @[playground/src/sim/sim_core.scala 21:26]
  wire [31:0] crossBar_io_memAxi_wa_bits_addr; // @[playground/src/sim/sim_core.scala 21:26]
  wire [7:0] crossBar_io_memAxi_wa_bits_len; // @[playground/src/sim/sim_core.scala 21:26]
  wire [2:0] crossBar_io_memAxi_wa_bits_size; // @[playground/src/sim/sim_core.scala 21:26]
  wire [1:0] crossBar_io_memAxi_wa_bits_burst; // @[playground/src/sim/sim_core.scala 21:26]
  wire  crossBar_io_memAxi_wd_ready; // @[playground/src/sim/sim_core.scala 21:26]
  wire  crossBar_io_memAxi_wd_valid; // @[playground/src/sim/sim_core.scala 21:26]
  wire [63:0] crossBar_io_memAxi_wd_bits_data; // @[playground/src/sim/sim_core.scala 21:26]
  wire [7:0] crossBar_io_memAxi_wd_bits_strb; // @[playground/src/sim/sim_core.scala 21:26]
  wire  crossBar_io_memAxi_wd_bits_last; // @[playground/src/sim/sim_core.scala 21:26]
  wire  crossBar_io_memAxi_wr_ready; // @[playground/src/sim/sim_core.scala 21:26]
  wire  crossBar_io_memAxi_wr_valid; // @[playground/src/sim/sim_core.scala 21:26]
  wire [3:0] crossBar_io_memAxi_wr_bits_id; // @[playground/src/sim/sim_core.scala 21:26]
  wire [1:0] crossBar_io_memAxi_wr_bits_resp; // @[playground/src/sim/sim_core.scala 21:26]
  wire  crossBar_io_memAxi_ra_ready; // @[playground/src/sim/sim_core.scala 21:26]
  wire  crossBar_io_memAxi_ra_valid; // @[playground/src/sim/sim_core.scala 21:26]
  wire [3:0] crossBar_io_memAxi_ra_bits_id; // @[playground/src/sim/sim_core.scala 21:26]
  wire [31:0] crossBar_io_memAxi_ra_bits_addr; // @[playground/src/sim/sim_core.scala 21:26]
  wire [7:0] crossBar_io_memAxi_ra_bits_len; // @[playground/src/sim/sim_core.scala 21:26]
  wire [2:0] crossBar_io_memAxi_ra_bits_size; // @[playground/src/sim/sim_core.scala 21:26]
  wire [1:0] crossBar_io_memAxi_ra_bits_burst; // @[playground/src/sim/sim_core.scala 21:26]
  wire  crossBar_io_memAxi_rd_ready; // @[playground/src/sim/sim_core.scala 21:26]
  wire  crossBar_io_memAxi_rd_valid; // @[playground/src/sim/sim_core.scala 21:26]
  wire [3:0] crossBar_io_memAxi_rd_bits_id; // @[playground/src/sim/sim_core.scala 21:26]
  wire [63:0] crossBar_io_memAxi_rd_bits_data; // @[playground/src/sim/sim_core.scala 21:26]
  wire [1:0] crossBar_io_memAxi_rd_bits_resp; // @[playground/src/sim/sim_core.scala 21:26]
  wire  crossBar_io_memAxi_rd_bits_last; // @[playground/src/sim/sim_core.scala 21:26]
  wire  crossBar_io_mmioAxi_wa_ready; // @[playground/src/sim/sim_core.scala 21:26]
  wire  crossBar_io_mmioAxi_wa_valid; // @[playground/src/sim/sim_core.scala 21:26]
  wire [31:0] crossBar_io_mmioAxi_wa_bits_addr; // @[playground/src/sim/sim_core.scala 21:26]
  wire  crossBar_io_mmioAxi_wd_ready; // @[playground/src/sim/sim_core.scala 21:26]
  wire  crossBar_io_mmioAxi_wd_valid; // @[playground/src/sim/sim_core.scala 21:26]
  wire [63:0] crossBar_io_mmioAxi_wd_bits_data; // @[playground/src/sim/sim_core.scala 21:26]
  wire [7:0] crossBar_io_mmioAxi_wd_bits_strb; // @[playground/src/sim/sim_core.scala 21:26]
  wire  crossBar_io_mmioAxi_wd_bits_last; // @[playground/src/sim/sim_core.scala 21:26]
  wire  crossBar_io_mmioAxi_ra_ready; // @[playground/src/sim/sim_core.scala 21:26]
  wire  crossBar_io_mmioAxi_ra_valid; // @[playground/src/sim/sim_core.scala 21:26]
  wire [31:0] crossBar_io_mmioAxi_ra_bits_addr; // @[playground/src/sim/sim_core.scala 21:26]
  wire  crossBar_io_mmioAxi_rd_ready; // @[playground/src/sim/sim_core.scala 21:26]
  wire  crossBar_io_mmioAxi_rd_valid; // @[playground/src/sim/sim_core.scala 21:26]
  wire [63:0] crossBar_io_mmioAxi_rd_bits_data; // @[playground/src/sim/sim_core.scala 21:26]
  wire  crossBar_io_mmioAxi_rd_bits_last; // @[playground/src/sim/sim_core.scala 21:26]
  wire  transAxi_io_raw_axi_awready; // @[playground/src/sim/sim_core.scala 22:26]
  wire  transAxi_io_raw_axi_awvalid; // @[playground/src/sim/sim_core.scala 22:26]
  wire [31:0] transAxi_io_raw_axi_awaddr; // @[playground/src/sim/sim_core.scala 22:26]
  wire [3:0] transAxi_io_raw_axi_awid; // @[playground/src/sim/sim_core.scala 22:26]
  wire [7:0] transAxi_io_raw_axi_awlen; // @[playground/src/sim/sim_core.scala 22:26]
  wire [2:0] transAxi_io_raw_axi_awsize; // @[playground/src/sim/sim_core.scala 22:26]
  wire [1:0] transAxi_io_raw_axi_awburst; // @[playground/src/sim/sim_core.scala 22:26]
  wire  transAxi_io_raw_axi_wready; // @[playground/src/sim/sim_core.scala 22:26]
  wire  transAxi_io_raw_axi_wvalid; // @[playground/src/sim/sim_core.scala 22:26]
  wire [63:0] transAxi_io_raw_axi_wdata; // @[playground/src/sim/sim_core.scala 22:26]
  wire [7:0] transAxi_io_raw_axi_wstrb; // @[playground/src/sim/sim_core.scala 22:26]
  wire  transAxi_io_raw_axi_wlast; // @[playground/src/sim/sim_core.scala 22:26]
  wire  transAxi_io_raw_axi_bready; // @[playground/src/sim/sim_core.scala 22:26]
  wire  transAxi_io_raw_axi_bvalid; // @[playground/src/sim/sim_core.scala 22:26]
  wire [1:0] transAxi_io_raw_axi_bresp; // @[playground/src/sim/sim_core.scala 22:26]
  wire [3:0] transAxi_io_raw_axi_bid; // @[playground/src/sim/sim_core.scala 22:26]
  wire  transAxi_io_raw_axi_arready; // @[playground/src/sim/sim_core.scala 22:26]
  wire  transAxi_io_raw_axi_arvalid; // @[playground/src/sim/sim_core.scala 22:26]
  wire [31:0] transAxi_io_raw_axi_araddr; // @[playground/src/sim/sim_core.scala 22:26]
  wire [3:0] transAxi_io_raw_axi_arid; // @[playground/src/sim/sim_core.scala 22:26]
  wire [7:0] transAxi_io_raw_axi_arlen; // @[playground/src/sim/sim_core.scala 22:26]
  wire [2:0] transAxi_io_raw_axi_arsize; // @[playground/src/sim/sim_core.scala 22:26]
  wire [1:0] transAxi_io_raw_axi_arburst; // @[playground/src/sim/sim_core.scala 22:26]
  wire  transAxi_io_raw_axi_rready; // @[playground/src/sim/sim_core.scala 22:26]
  wire  transAxi_io_raw_axi_rvalid; // @[playground/src/sim/sim_core.scala 22:26]
  wire [1:0] transAxi_io_raw_axi_rresp; // @[playground/src/sim/sim_core.scala 22:26]
  wire [63:0] transAxi_io_raw_axi_rdata; // @[playground/src/sim/sim_core.scala 22:26]
  wire  transAxi_io_raw_axi_rlast; // @[playground/src/sim/sim_core.scala 22:26]
  wire [3:0] transAxi_io_raw_axi_rid; // @[playground/src/sim/sim_core.scala 22:26]
  wire  transAxi_io_bun_axi_wa_ready; // @[playground/src/sim/sim_core.scala 22:26]
  wire  transAxi_io_bun_axi_wa_valid; // @[playground/src/sim/sim_core.scala 22:26]
  wire [3:0] transAxi_io_bun_axi_wa_bits_id; // @[playground/src/sim/sim_core.scala 22:26]
  wire [31:0] transAxi_io_bun_axi_wa_bits_addr; // @[playground/src/sim/sim_core.scala 22:26]
  wire [7:0] transAxi_io_bun_axi_wa_bits_len; // @[playground/src/sim/sim_core.scala 22:26]
  wire [2:0] transAxi_io_bun_axi_wa_bits_size; // @[playground/src/sim/sim_core.scala 22:26]
  wire [1:0] transAxi_io_bun_axi_wa_bits_burst; // @[playground/src/sim/sim_core.scala 22:26]
  wire  transAxi_io_bun_axi_wd_ready; // @[playground/src/sim/sim_core.scala 22:26]
  wire  transAxi_io_bun_axi_wd_valid; // @[playground/src/sim/sim_core.scala 22:26]
  wire [63:0] transAxi_io_bun_axi_wd_bits_data; // @[playground/src/sim/sim_core.scala 22:26]
  wire [7:0] transAxi_io_bun_axi_wd_bits_strb; // @[playground/src/sim/sim_core.scala 22:26]
  wire  transAxi_io_bun_axi_wd_bits_last; // @[playground/src/sim/sim_core.scala 22:26]
  wire  transAxi_io_bun_axi_wr_ready; // @[playground/src/sim/sim_core.scala 22:26]
  wire  transAxi_io_bun_axi_wr_valid; // @[playground/src/sim/sim_core.scala 22:26]
  wire [3:0] transAxi_io_bun_axi_wr_bits_id; // @[playground/src/sim/sim_core.scala 22:26]
  wire [1:0] transAxi_io_bun_axi_wr_bits_resp; // @[playground/src/sim/sim_core.scala 22:26]
  wire  transAxi_io_bun_axi_ra_ready; // @[playground/src/sim/sim_core.scala 22:26]
  wire  transAxi_io_bun_axi_ra_valid; // @[playground/src/sim/sim_core.scala 22:26]
  wire [3:0] transAxi_io_bun_axi_ra_bits_id; // @[playground/src/sim/sim_core.scala 22:26]
  wire [31:0] transAxi_io_bun_axi_ra_bits_addr; // @[playground/src/sim/sim_core.scala 22:26]
  wire [7:0] transAxi_io_bun_axi_ra_bits_len; // @[playground/src/sim/sim_core.scala 22:26]
  wire [2:0] transAxi_io_bun_axi_ra_bits_size; // @[playground/src/sim/sim_core.scala 22:26]
  wire [1:0] transAxi_io_bun_axi_ra_bits_burst; // @[playground/src/sim/sim_core.scala 22:26]
  wire  transAxi_io_bun_axi_rd_ready; // @[playground/src/sim/sim_core.scala 22:26]
  wire  transAxi_io_bun_axi_rd_valid; // @[playground/src/sim/sim_core.scala 22:26]
  wire [3:0] transAxi_io_bun_axi_rd_bits_id; // @[playground/src/sim/sim_core.scala 22:26]
  wire [63:0] transAxi_io_bun_axi_rd_bits_data; // @[playground/src/sim/sim_core.scala 22:26]
  wire [1:0] transAxi_io_bun_axi_rd_bits_resp; // @[playground/src/sim/sim_core.scala 22:26]
  wire  transAxi_io_bun_axi_rd_bits_last; // @[playground/src/sim/sim_core.scala 22:26]
  CPU cpu ( // @[playground/src/sim/sim_core.scala 17:21]
    .clock(cpu_clock),
    .reset(cpu_reset),
    .io_master_awready(cpu_io_master_awready),
    .io_master_awvalid(cpu_io_master_awvalid),
    .io_master_awaddr(cpu_io_master_awaddr),
    .io_master_awid(cpu_io_master_awid),
    .io_master_awlen(cpu_io_master_awlen),
    .io_master_awsize(cpu_io_master_awsize),
    .io_master_awburst(cpu_io_master_awburst),
    .io_master_wready(cpu_io_master_wready),
    .io_master_wvalid(cpu_io_master_wvalid),
    .io_master_wdata(cpu_io_master_wdata),
    .io_master_wstrb(cpu_io_master_wstrb),
    .io_master_wlast(cpu_io_master_wlast),
    .io_master_bready(cpu_io_master_bready),
    .io_master_bvalid(cpu_io_master_bvalid),
    .io_master_bresp(cpu_io_master_bresp),
    .io_master_bid(cpu_io_master_bid),
    .io_master_arready(cpu_io_master_arready),
    .io_master_arvalid(cpu_io_master_arvalid),
    .io_master_araddr(cpu_io_master_araddr),
    .io_master_arid(cpu_io_master_arid),
    .io_master_arlen(cpu_io_master_arlen),
    .io_master_arsize(cpu_io_master_arsize),
    .io_master_arburst(cpu_io_master_arburst),
    .io_master_rready(cpu_io_master_rready),
    .io_master_rvalid(cpu_io_master_rvalid),
    .io_master_rresp(cpu_io_master_rresp),
    .io_master_rdata(cpu_io_master_rdata),
    .io_master_rlast(cpu_io_master_rlast),
    .io_master_rid(cpu_io_master_rid),
    .io_slave_awready(cpu_io_slave_awready),
    .io_slave_awvalid(cpu_io_slave_awvalid),
    .io_slave_awaddr(cpu_io_slave_awaddr),
    .io_slave_awid(cpu_io_slave_awid),
    .io_slave_awlen(cpu_io_slave_awlen),
    .io_slave_awsize(cpu_io_slave_awsize),
    .io_slave_awburst(cpu_io_slave_awburst),
    .io_slave_wready(cpu_io_slave_wready),
    .io_slave_wvalid(cpu_io_slave_wvalid),
    .io_slave_wdata(cpu_io_slave_wdata),
    .io_slave_wstrb(cpu_io_slave_wstrb),
    .io_slave_wlast(cpu_io_slave_wlast),
    .io_slave_bready(cpu_io_slave_bready),
    .io_slave_bvalid(cpu_io_slave_bvalid),
    .io_slave_bresp(cpu_io_slave_bresp),
    .io_slave_bid(cpu_io_slave_bid),
    .io_slave_arready(cpu_io_slave_arready),
    .io_slave_arvalid(cpu_io_slave_arvalid),
    .io_slave_araddr(cpu_io_slave_araddr),
    .io_slave_arid(cpu_io_slave_arid),
    .io_slave_arlen(cpu_io_slave_arlen),
    .io_slave_arsize(cpu_io_slave_arsize),
    .io_slave_arburst(cpu_io_slave_arburst),
    .io_slave_rready(cpu_io_slave_rready),
    .io_slave_rvalid(cpu_io_slave_rvalid),
    .io_slave_rresp(cpu_io_slave_rresp),
    .io_slave_rdata(cpu_io_slave_rdata),
    .io_slave_rlast(cpu_io_slave_rlast),
    .io_slave_rid(cpu_io_slave_rid),
    .io_interrupt(cpu_io_interrupt)
  );
  SimMEM mem ( // @[playground/src/sim/sim_core.scala 18:21]
    .clock(mem_clock),
    .reset(mem_reset),
    .io_memAxi_wa_ready(mem_io_memAxi_wa_ready),
    .io_memAxi_wa_valid(mem_io_memAxi_wa_valid),
    .io_memAxi_wa_bits_id(mem_io_memAxi_wa_bits_id),
    .io_memAxi_wa_bits_addr(mem_io_memAxi_wa_bits_addr),
    .io_memAxi_wa_bits_len(mem_io_memAxi_wa_bits_len),
    .io_memAxi_wa_bits_size(mem_io_memAxi_wa_bits_size),
    .io_memAxi_wa_bits_burst(mem_io_memAxi_wa_bits_burst),
    .io_memAxi_wd_ready(mem_io_memAxi_wd_ready),
    .io_memAxi_wd_valid(mem_io_memAxi_wd_valid),
    .io_memAxi_wd_bits_data(mem_io_memAxi_wd_bits_data),
    .io_memAxi_wd_bits_strb(mem_io_memAxi_wd_bits_strb),
    .io_memAxi_wd_bits_last(mem_io_memAxi_wd_bits_last),
    .io_memAxi_wr_ready(mem_io_memAxi_wr_ready),
    .io_memAxi_wr_valid(mem_io_memAxi_wr_valid),
    .io_memAxi_wr_bits_id(mem_io_memAxi_wr_bits_id),
    .io_memAxi_wr_bits_resp(mem_io_memAxi_wr_bits_resp),
    .io_memAxi_ra_ready(mem_io_memAxi_ra_ready),
    .io_memAxi_ra_valid(mem_io_memAxi_ra_valid),
    .io_memAxi_ra_bits_id(mem_io_memAxi_ra_bits_id),
    .io_memAxi_ra_bits_addr(mem_io_memAxi_ra_bits_addr),
    .io_memAxi_ra_bits_len(mem_io_memAxi_ra_bits_len),
    .io_memAxi_ra_bits_size(mem_io_memAxi_ra_bits_size),
    .io_memAxi_ra_bits_burst(mem_io_memAxi_ra_bits_burst),
    .io_memAxi_rd_ready(mem_io_memAxi_rd_ready),
    .io_memAxi_rd_valid(mem_io_memAxi_rd_valid),
    .io_memAxi_rd_bits_id(mem_io_memAxi_rd_bits_id),
    .io_memAxi_rd_bits_data(mem_io_memAxi_rd_bits_data),
    .io_memAxi_rd_bits_resp(mem_io_memAxi_rd_bits_resp),
    .io_memAxi_rd_bits_last(mem_io_memAxi_rd_bits_last)
  );
  SimMMIO mmio ( // @[playground/src/sim/sim_core.scala 19:22]
    .clock(mmio_clock),
    .reset(mmio_reset),
    .io_mmioAxi_wa_ready(mmio_io_mmioAxi_wa_ready),
    .io_mmioAxi_wa_valid(mmio_io_mmioAxi_wa_valid),
    .io_mmioAxi_wa_bits_addr(mmio_io_mmioAxi_wa_bits_addr),
    .io_mmioAxi_wd_ready(mmio_io_mmioAxi_wd_ready),
    .io_mmioAxi_wd_valid(mmio_io_mmioAxi_wd_valid),
    .io_mmioAxi_wd_bits_data(mmio_io_mmioAxi_wd_bits_data),
    .io_mmioAxi_wd_bits_strb(mmio_io_mmioAxi_wd_bits_strb),
    .io_mmioAxi_wd_bits_last(mmio_io_mmioAxi_wd_bits_last),
    .io_mmioAxi_ra_ready(mmio_io_mmioAxi_ra_ready),
    .io_mmioAxi_ra_valid(mmio_io_mmioAxi_ra_valid),
    .io_mmioAxi_ra_bits_addr(mmio_io_mmioAxi_ra_bits_addr),
    .io_mmioAxi_rd_ready(mmio_io_mmioAxi_rd_ready),
    .io_mmioAxi_rd_valid(mmio_io_mmioAxi_rd_valid),
    .io_mmioAxi_rd_bits_data(mmio_io_mmioAxi_rd_bits_data),
    .io_mmioAxi_rd_bits_last(mmio_io_mmioAxi_rd_bits_last)
  );
  SimDma dma ( // @[playground/src/sim/sim_core.scala 20:21]
    .clock(dma_clock),
    .reset(dma_reset),
    .io_dmaAxi_wstrb(dma_io_dmaAxi_wstrb)
  );
  SimCrossbar crossBar ( // @[playground/src/sim/sim_core.scala 21:26]
    .clock(crossBar_clock),
    .reset(crossBar_reset),
    .io_inAxi_wa_ready(crossBar_io_inAxi_wa_ready),
    .io_inAxi_wa_valid(crossBar_io_inAxi_wa_valid),
    .io_inAxi_wa_bits_id(crossBar_io_inAxi_wa_bits_id),
    .io_inAxi_wa_bits_addr(crossBar_io_inAxi_wa_bits_addr),
    .io_inAxi_wa_bits_len(crossBar_io_inAxi_wa_bits_len),
    .io_inAxi_wa_bits_size(crossBar_io_inAxi_wa_bits_size),
    .io_inAxi_wa_bits_burst(crossBar_io_inAxi_wa_bits_burst),
    .io_inAxi_wd_ready(crossBar_io_inAxi_wd_ready),
    .io_inAxi_wd_valid(crossBar_io_inAxi_wd_valid),
    .io_inAxi_wd_bits_data(crossBar_io_inAxi_wd_bits_data),
    .io_inAxi_wd_bits_strb(crossBar_io_inAxi_wd_bits_strb),
    .io_inAxi_wd_bits_last(crossBar_io_inAxi_wd_bits_last),
    .io_inAxi_wr_ready(crossBar_io_inAxi_wr_ready),
    .io_inAxi_wr_valid(crossBar_io_inAxi_wr_valid),
    .io_inAxi_wr_bits_id(crossBar_io_inAxi_wr_bits_id),
    .io_inAxi_wr_bits_resp(crossBar_io_inAxi_wr_bits_resp),
    .io_inAxi_ra_ready(crossBar_io_inAxi_ra_ready),
    .io_inAxi_ra_valid(crossBar_io_inAxi_ra_valid),
    .io_inAxi_ra_bits_id(crossBar_io_inAxi_ra_bits_id),
    .io_inAxi_ra_bits_addr(crossBar_io_inAxi_ra_bits_addr),
    .io_inAxi_ra_bits_len(crossBar_io_inAxi_ra_bits_len),
    .io_inAxi_ra_bits_size(crossBar_io_inAxi_ra_bits_size),
    .io_inAxi_ra_bits_burst(crossBar_io_inAxi_ra_bits_burst),
    .io_inAxi_rd_ready(crossBar_io_inAxi_rd_ready),
    .io_inAxi_rd_valid(crossBar_io_inAxi_rd_valid),
    .io_inAxi_rd_bits_id(crossBar_io_inAxi_rd_bits_id),
    .io_inAxi_rd_bits_data(crossBar_io_inAxi_rd_bits_data),
    .io_inAxi_rd_bits_resp(crossBar_io_inAxi_rd_bits_resp),
    .io_inAxi_rd_bits_last(crossBar_io_inAxi_rd_bits_last),
    .io_memAxi_wa_ready(crossBar_io_memAxi_wa_ready),
    .io_memAxi_wa_valid(crossBar_io_memAxi_wa_valid),
    .io_memAxi_wa_bits_id(crossBar_io_memAxi_wa_bits_id),
    .io_memAxi_wa_bits_addr(crossBar_io_memAxi_wa_bits_addr),
    .io_memAxi_wa_bits_len(crossBar_io_memAxi_wa_bits_len),
    .io_memAxi_wa_bits_size(crossBar_io_memAxi_wa_bits_size),
    .io_memAxi_wa_bits_burst(crossBar_io_memAxi_wa_bits_burst),
    .io_memAxi_wd_ready(crossBar_io_memAxi_wd_ready),
    .io_memAxi_wd_valid(crossBar_io_memAxi_wd_valid),
    .io_memAxi_wd_bits_data(crossBar_io_memAxi_wd_bits_data),
    .io_memAxi_wd_bits_strb(crossBar_io_memAxi_wd_bits_strb),
    .io_memAxi_wd_bits_last(crossBar_io_memAxi_wd_bits_last),
    .io_memAxi_wr_ready(crossBar_io_memAxi_wr_ready),
    .io_memAxi_wr_valid(crossBar_io_memAxi_wr_valid),
    .io_memAxi_wr_bits_id(crossBar_io_memAxi_wr_bits_id),
    .io_memAxi_wr_bits_resp(crossBar_io_memAxi_wr_bits_resp),
    .io_memAxi_ra_ready(crossBar_io_memAxi_ra_ready),
    .io_memAxi_ra_valid(crossBar_io_memAxi_ra_valid),
    .io_memAxi_ra_bits_id(crossBar_io_memAxi_ra_bits_id),
    .io_memAxi_ra_bits_addr(crossBar_io_memAxi_ra_bits_addr),
    .io_memAxi_ra_bits_len(crossBar_io_memAxi_ra_bits_len),
    .io_memAxi_ra_bits_size(crossBar_io_memAxi_ra_bits_size),
    .io_memAxi_ra_bits_burst(crossBar_io_memAxi_ra_bits_burst),
    .io_memAxi_rd_ready(crossBar_io_memAxi_rd_ready),
    .io_memAxi_rd_valid(crossBar_io_memAxi_rd_valid),
    .io_memAxi_rd_bits_id(crossBar_io_memAxi_rd_bits_id),
    .io_memAxi_rd_bits_data(crossBar_io_memAxi_rd_bits_data),
    .io_memAxi_rd_bits_resp(crossBar_io_memAxi_rd_bits_resp),
    .io_memAxi_rd_bits_last(crossBar_io_memAxi_rd_bits_last),
    .io_mmioAxi_wa_ready(crossBar_io_mmioAxi_wa_ready),
    .io_mmioAxi_wa_valid(crossBar_io_mmioAxi_wa_valid),
    .io_mmioAxi_wa_bits_addr(crossBar_io_mmioAxi_wa_bits_addr),
    .io_mmioAxi_wd_ready(crossBar_io_mmioAxi_wd_ready),
    .io_mmioAxi_wd_valid(crossBar_io_mmioAxi_wd_valid),
    .io_mmioAxi_wd_bits_data(crossBar_io_mmioAxi_wd_bits_data),
    .io_mmioAxi_wd_bits_strb(crossBar_io_mmioAxi_wd_bits_strb),
    .io_mmioAxi_wd_bits_last(crossBar_io_mmioAxi_wd_bits_last),
    .io_mmioAxi_ra_ready(crossBar_io_mmioAxi_ra_ready),
    .io_mmioAxi_ra_valid(crossBar_io_mmioAxi_ra_valid),
    .io_mmioAxi_ra_bits_addr(crossBar_io_mmioAxi_ra_bits_addr),
    .io_mmioAxi_rd_ready(crossBar_io_mmioAxi_rd_ready),
    .io_mmioAxi_rd_valid(crossBar_io_mmioAxi_rd_valid),
    .io_mmioAxi_rd_bits_data(crossBar_io_mmioAxi_rd_bits_data),
    .io_mmioAxi_rd_bits_last(crossBar_io_mmioAxi_rd_bits_last)
  );
  TransAXI transAxi ( // @[playground/src/sim/sim_core.scala 22:26]
    .io_raw_axi_awready(transAxi_io_raw_axi_awready),
    .io_raw_axi_awvalid(transAxi_io_raw_axi_awvalid),
    .io_raw_axi_awaddr(transAxi_io_raw_axi_awaddr),
    .io_raw_axi_awid(transAxi_io_raw_axi_awid),
    .io_raw_axi_awlen(transAxi_io_raw_axi_awlen),
    .io_raw_axi_awsize(transAxi_io_raw_axi_awsize),
    .io_raw_axi_awburst(transAxi_io_raw_axi_awburst),
    .io_raw_axi_wready(transAxi_io_raw_axi_wready),
    .io_raw_axi_wvalid(transAxi_io_raw_axi_wvalid),
    .io_raw_axi_wdata(transAxi_io_raw_axi_wdata),
    .io_raw_axi_wstrb(transAxi_io_raw_axi_wstrb),
    .io_raw_axi_wlast(transAxi_io_raw_axi_wlast),
    .io_raw_axi_bready(transAxi_io_raw_axi_bready),
    .io_raw_axi_bvalid(transAxi_io_raw_axi_bvalid),
    .io_raw_axi_bresp(transAxi_io_raw_axi_bresp),
    .io_raw_axi_bid(transAxi_io_raw_axi_bid),
    .io_raw_axi_arready(transAxi_io_raw_axi_arready),
    .io_raw_axi_arvalid(transAxi_io_raw_axi_arvalid),
    .io_raw_axi_araddr(transAxi_io_raw_axi_araddr),
    .io_raw_axi_arid(transAxi_io_raw_axi_arid),
    .io_raw_axi_arlen(transAxi_io_raw_axi_arlen),
    .io_raw_axi_arsize(transAxi_io_raw_axi_arsize),
    .io_raw_axi_arburst(transAxi_io_raw_axi_arburst),
    .io_raw_axi_rready(transAxi_io_raw_axi_rready),
    .io_raw_axi_rvalid(transAxi_io_raw_axi_rvalid),
    .io_raw_axi_rresp(transAxi_io_raw_axi_rresp),
    .io_raw_axi_rdata(transAxi_io_raw_axi_rdata),
    .io_raw_axi_rlast(transAxi_io_raw_axi_rlast),
    .io_raw_axi_rid(transAxi_io_raw_axi_rid),
    .io_bun_axi_wa_ready(transAxi_io_bun_axi_wa_ready),
    .io_bun_axi_wa_valid(transAxi_io_bun_axi_wa_valid),
    .io_bun_axi_wa_bits_id(transAxi_io_bun_axi_wa_bits_id),
    .io_bun_axi_wa_bits_addr(transAxi_io_bun_axi_wa_bits_addr),
    .io_bun_axi_wa_bits_len(transAxi_io_bun_axi_wa_bits_len),
    .io_bun_axi_wa_bits_size(transAxi_io_bun_axi_wa_bits_size),
    .io_bun_axi_wa_bits_burst(transAxi_io_bun_axi_wa_bits_burst),
    .io_bun_axi_wd_ready(transAxi_io_bun_axi_wd_ready),
    .io_bun_axi_wd_valid(transAxi_io_bun_axi_wd_valid),
    .io_bun_axi_wd_bits_data(transAxi_io_bun_axi_wd_bits_data),
    .io_bun_axi_wd_bits_strb(transAxi_io_bun_axi_wd_bits_strb),
    .io_bun_axi_wd_bits_last(transAxi_io_bun_axi_wd_bits_last),
    .io_bun_axi_wr_ready(transAxi_io_bun_axi_wr_ready),
    .io_bun_axi_wr_valid(transAxi_io_bun_axi_wr_valid),
    .io_bun_axi_wr_bits_id(transAxi_io_bun_axi_wr_bits_id),
    .io_bun_axi_wr_bits_resp(transAxi_io_bun_axi_wr_bits_resp),
    .io_bun_axi_ra_ready(transAxi_io_bun_axi_ra_ready),
    .io_bun_axi_ra_valid(transAxi_io_bun_axi_ra_valid),
    .io_bun_axi_ra_bits_id(transAxi_io_bun_axi_ra_bits_id),
    .io_bun_axi_ra_bits_addr(transAxi_io_bun_axi_ra_bits_addr),
    .io_bun_axi_ra_bits_len(transAxi_io_bun_axi_ra_bits_len),
    .io_bun_axi_ra_bits_size(transAxi_io_bun_axi_ra_bits_size),
    .io_bun_axi_ra_bits_burst(transAxi_io_bun_axi_ra_bits_burst),
    .io_bun_axi_rd_ready(transAxi_io_bun_axi_rd_ready),
    .io_bun_axi_rd_valid(transAxi_io_bun_axi_rd_valid),
    .io_bun_axi_rd_bits_id(transAxi_io_bun_axi_rd_bits_id),
    .io_bun_axi_rd_bits_data(transAxi_io_bun_axi_rd_bits_data),
    .io_bun_axi_rd_bits_resp(transAxi_io_bun_axi_rd_bits_resp),
    .io_bun_axi_rd_bits_last(transAxi_io_bun_axi_rd_bits_last)
  );
  assign cpu_clock = clock;
  assign cpu_reset = reset;
  assign cpu_io_master_awready = transAxi_io_raw_axi_awready; // @[playground/src/sim/sim_core.scala 23:19]
  assign cpu_io_master_wready = transAxi_io_raw_axi_wready; // @[playground/src/sim/sim_core.scala 23:19]
  assign cpu_io_master_bvalid = transAxi_io_raw_axi_bvalid; // @[playground/src/sim/sim_core.scala 23:19]
  assign cpu_io_master_bresp = transAxi_io_raw_axi_bresp; // @[playground/src/sim/sim_core.scala 23:19]
  assign cpu_io_master_bid = transAxi_io_raw_axi_bid; // @[playground/src/sim/sim_core.scala 23:19]
  assign cpu_io_master_arready = transAxi_io_raw_axi_arready; // @[playground/src/sim/sim_core.scala 23:19]
  assign cpu_io_master_rvalid = transAxi_io_raw_axi_rvalid; // @[playground/src/sim/sim_core.scala 23:19]
  assign cpu_io_master_rresp = transAxi_io_raw_axi_rresp; // @[playground/src/sim/sim_core.scala 23:19]
  assign cpu_io_master_rdata = transAxi_io_raw_axi_rdata; // @[playground/src/sim/sim_core.scala 23:19]
  assign cpu_io_master_rlast = transAxi_io_raw_axi_rlast; // @[playground/src/sim/sim_core.scala 23:19]
  assign cpu_io_master_rid = transAxi_io_raw_axi_rid; // @[playground/src/sim/sim_core.scala 23:19]
  assign cpu_io_slave_awvalid = 1'h0; // @[playground/src/sim/sim_core.scala 27:19]
  assign cpu_io_slave_awaddr = 32'h0; // @[playground/src/sim/sim_core.scala 27:19]
  assign cpu_io_slave_awid = 4'h0; // @[playground/src/sim/sim_core.scala 27:19]
  assign cpu_io_slave_awlen = 8'h0; // @[playground/src/sim/sim_core.scala 27:19]
  assign cpu_io_slave_awsize = 3'h0; // @[playground/src/sim/sim_core.scala 27:19]
  assign cpu_io_slave_awburst = 2'h0; // @[playground/src/sim/sim_core.scala 27:19]
  assign cpu_io_slave_wvalid = 1'h0; // @[playground/src/sim/sim_core.scala 27:19]
  assign cpu_io_slave_wdata = 64'h0; // @[playground/src/sim/sim_core.scala 27:19]
  assign cpu_io_slave_wstrb = dma_io_dmaAxi_wstrb; // @[playground/src/sim/sim_core.scala 27:19]
  assign cpu_io_slave_wlast = 1'h0; // @[playground/src/sim/sim_core.scala 27:19]
  assign cpu_io_slave_bready = 1'h0; // @[playground/src/sim/sim_core.scala 27:19]
  assign cpu_io_slave_arvalid = 1'h0; // @[playground/src/sim/sim_core.scala 27:19]
  assign cpu_io_slave_araddr = 32'h0; // @[playground/src/sim/sim_core.scala 27:19]
  assign cpu_io_slave_arid = 4'h0; // @[playground/src/sim/sim_core.scala 27:19]
  assign cpu_io_slave_arlen = 8'h0; // @[playground/src/sim/sim_core.scala 27:19]
  assign cpu_io_slave_arsize = 3'h0; // @[playground/src/sim/sim_core.scala 27:19]
  assign cpu_io_slave_arburst = 2'h0; // @[playground/src/sim/sim_core.scala 27:19]
  assign cpu_io_slave_rready = 1'h0; // @[playground/src/sim/sim_core.scala 27:19]
  assign cpu_io_interrupt = 1'h0; // @[playground/src/sim/sim_core.scala 31:36]
  assign mem_clock = clock;
  assign mem_reset = reset;
  assign mem_io_memAxi_wa_valid = crossBar_io_memAxi_wa_valid; // @[playground/src/sim/sim_core.scala 26:24]
  assign mem_io_memAxi_wa_bits_id = crossBar_io_memAxi_wa_bits_id; // @[playground/src/sim/sim_core.scala 26:24]
  assign mem_io_memAxi_wa_bits_addr = crossBar_io_memAxi_wa_bits_addr; // @[playground/src/sim/sim_core.scala 26:24]
  assign mem_io_memAxi_wa_bits_len = crossBar_io_memAxi_wa_bits_len; // @[playground/src/sim/sim_core.scala 26:24]
  assign mem_io_memAxi_wa_bits_size = crossBar_io_memAxi_wa_bits_size; // @[playground/src/sim/sim_core.scala 26:24]
  assign mem_io_memAxi_wa_bits_burst = crossBar_io_memAxi_wa_bits_burst; // @[playground/src/sim/sim_core.scala 26:24]
  assign mem_io_memAxi_wd_valid = crossBar_io_memAxi_wd_valid; // @[playground/src/sim/sim_core.scala 26:24]
  assign mem_io_memAxi_wd_bits_data = crossBar_io_memAxi_wd_bits_data; // @[playground/src/sim/sim_core.scala 26:24]
  assign mem_io_memAxi_wd_bits_strb = crossBar_io_memAxi_wd_bits_strb; // @[playground/src/sim/sim_core.scala 26:24]
  assign mem_io_memAxi_wd_bits_last = crossBar_io_memAxi_wd_bits_last; // @[playground/src/sim/sim_core.scala 26:24]
  assign mem_io_memAxi_wr_ready = crossBar_io_memAxi_wr_ready; // @[playground/src/sim/sim_core.scala 26:24]
  assign mem_io_memAxi_ra_valid = crossBar_io_memAxi_ra_valid; // @[playground/src/sim/sim_core.scala 26:24]
  assign mem_io_memAxi_ra_bits_id = crossBar_io_memAxi_ra_bits_id; // @[playground/src/sim/sim_core.scala 26:24]
  assign mem_io_memAxi_ra_bits_addr = crossBar_io_memAxi_ra_bits_addr; // @[playground/src/sim/sim_core.scala 26:24]
  assign mem_io_memAxi_ra_bits_len = crossBar_io_memAxi_ra_bits_len; // @[playground/src/sim/sim_core.scala 26:24]
  assign mem_io_memAxi_ra_bits_size = crossBar_io_memAxi_ra_bits_size; // @[playground/src/sim/sim_core.scala 26:24]
  assign mem_io_memAxi_ra_bits_burst = crossBar_io_memAxi_ra_bits_burst; // @[playground/src/sim/sim_core.scala 26:24]
  assign mem_io_memAxi_rd_ready = crossBar_io_memAxi_rd_ready; // @[playground/src/sim/sim_core.scala 26:24]
  assign mmio_clock = clock;
  assign mmio_reset = reset;
  assign mmio_io_mmioAxi_wa_valid = crossBar_io_mmioAxi_wa_valid; // @[playground/src/sim/sim_core.scala 25:25]
  assign mmio_io_mmioAxi_wa_bits_addr = crossBar_io_mmioAxi_wa_bits_addr; // @[playground/src/sim/sim_core.scala 25:25]
  assign mmio_io_mmioAxi_wd_valid = crossBar_io_mmioAxi_wd_valid; // @[playground/src/sim/sim_core.scala 25:25]
  assign mmio_io_mmioAxi_wd_bits_data = crossBar_io_mmioAxi_wd_bits_data; // @[playground/src/sim/sim_core.scala 25:25]
  assign mmio_io_mmioAxi_wd_bits_strb = crossBar_io_mmioAxi_wd_bits_strb; // @[playground/src/sim/sim_core.scala 25:25]
  assign mmio_io_mmioAxi_wd_bits_last = crossBar_io_mmioAxi_wd_bits_last; // @[playground/src/sim/sim_core.scala 25:25]
  assign mmio_io_mmioAxi_ra_valid = crossBar_io_mmioAxi_ra_valid; // @[playground/src/sim/sim_core.scala 25:25]
  assign mmio_io_mmioAxi_ra_bits_addr = crossBar_io_mmioAxi_ra_bits_addr; // @[playground/src/sim/sim_core.scala 25:25]
  assign mmio_io_mmioAxi_rd_ready = crossBar_io_mmioAxi_rd_ready; // @[playground/src/sim/sim_core.scala 25:25]
  assign dma_clock = clock;
  assign dma_reset = reset;
  assign crossBar_clock = clock;
  assign crossBar_reset = reset;
  assign crossBar_io_inAxi_wa_valid = transAxi_io_bun_axi_wa_valid; // @[playground/src/sim/sim_core.scala 24:25]
  assign crossBar_io_inAxi_wa_bits_id = transAxi_io_bun_axi_wa_bits_id; // @[playground/src/sim/sim_core.scala 24:25]
  assign crossBar_io_inAxi_wa_bits_addr = transAxi_io_bun_axi_wa_bits_addr; // @[playground/src/sim/sim_core.scala 24:25]
  assign crossBar_io_inAxi_wa_bits_len = transAxi_io_bun_axi_wa_bits_len; // @[playground/src/sim/sim_core.scala 24:25]
  assign crossBar_io_inAxi_wa_bits_size = transAxi_io_bun_axi_wa_bits_size; // @[playground/src/sim/sim_core.scala 24:25]
  assign crossBar_io_inAxi_wa_bits_burst = transAxi_io_bun_axi_wa_bits_burst; // @[playground/src/sim/sim_core.scala 24:25]
  assign crossBar_io_inAxi_wd_valid = transAxi_io_bun_axi_wd_valid; // @[playground/src/sim/sim_core.scala 24:25]
  assign crossBar_io_inAxi_wd_bits_data = transAxi_io_bun_axi_wd_bits_data; // @[playground/src/sim/sim_core.scala 24:25]
  assign crossBar_io_inAxi_wd_bits_strb = transAxi_io_bun_axi_wd_bits_strb; // @[playground/src/sim/sim_core.scala 24:25]
  assign crossBar_io_inAxi_wd_bits_last = transAxi_io_bun_axi_wd_bits_last; // @[playground/src/sim/sim_core.scala 24:25]
  assign crossBar_io_inAxi_wr_ready = transAxi_io_bun_axi_wr_ready; // @[playground/src/sim/sim_core.scala 24:25]
  assign crossBar_io_inAxi_ra_valid = transAxi_io_bun_axi_ra_valid; // @[playground/src/sim/sim_core.scala 24:25]
  assign crossBar_io_inAxi_ra_bits_id = transAxi_io_bun_axi_ra_bits_id; // @[playground/src/sim/sim_core.scala 24:25]
  assign crossBar_io_inAxi_ra_bits_addr = transAxi_io_bun_axi_ra_bits_addr; // @[playground/src/sim/sim_core.scala 24:25]
  assign crossBar_io_inAxi_ra_bits_len = transAxi_io_bun_axi_ra_bits_len; // @[playground/src/sim/sim_core.scala 24:25]
  assign crossBar_io_inAxi_ra_bits_size = transAxi_io_bun_axi_ra_bits_size; // @[playground/src/sim/sim_core.scala 24:25]
  assign crossBar_io_inAxi_ra_bits_burst = transAxi_io_bun_axi_ra_bits_burst; // @[playground/src/sim/sim_core.scala 24:25]
  assign crossBar_io_inAxi_rd_ready = transAxi_io_bun_axi_rd_ready; // @[playground/src/sim/sim_core.scala 24:25]
  assign crossBar_io_memAxi_wa_ready = mem_io_memAxi_wa_ready; // @[playground/src/sim/sim_core.scala 26:24]
  assign crossBar_io_memAxi_wd_ready = mem_io_memAxi_wd_ready; // @[playground/src/sim/sim_core.scala 26:24]
  assign crossBar_io_memAxi_wr_valid = mem_io_memAxi_wr_valid; // @[playground/src/sim/sim_core.scala 26:24]
  assign crossBar_io_memAxi_wr_bits_id = mem_io_memAxi_wr_bits_id; // @[playground/src/sim/sim_core.scala 26:24]
  assign crossBar_io_memAxi_wr_bits_resp = mem_io_memAxi_wr_bits_resp; // @[playground/src/sim/sim_core.scala 26:24]
  assign crossBar_io_memAxi_ra_ready = mem_io_memAxi_ra_ready; // @[playground/src/sim/sim_core.scala 26:24]
  assign crossBar_io_memAxi_rd_valid = mem_io_memAxi_rd_valid; // @[playground/src/sim/sim_core.scala 26:24]
  assign crossBar_io_memAxi_rd_bits_id = mem_io_memAxi_rd_bits_id; // @[playground/src/sim/sim_core.scala 26:24]
  assign crossBar_io_memAxi_rd_bits_data = mem_io_memAxi_rd_bits_data; // @[playground/src/sim/sim_core.scala 26:24]
  assign crossBar_io_memAxi_rd_bits_resp = mem_io_memAxi_rd_bits_resp; // @[playground/src/sim/sim_core.scala 26:24]
  assign crossBar_io_memAxi_rd_bits_last = mem_io_memAxi_rd_bits_last; // @[playground/src/sim/sim_core.scala 26:24]
  assign crossBar_io_mmioAxi_wa_ready = mmio_io_mmioAxi_wa_ready; // @[playground/src/sim/sim_core.scala 25:25]
  assign crossBar_io_mmioAxi_wd_ready = mmio_io_mmioAxi_wd_ready; // @[playground/src/sim/sim_core.scala 25:25]
  assign crossBar_io_mmioAxi_ra_ready = mmio_io_mmioAxi_ra_ready; // @[playground/src/sim/sim_core.scala 25:25]
  assign crossBar_io_mmioAxi_rd_valid = mmio_io_mmioAxi_rd_valid; // @[playground/src/sim/sim_core.scala 25:25]
  assign crossBar_io_mmioAxi_rd_bits_data = mmio_io_mmioAxi_rd_bits_data; // @[playground/src/sim/sim_core.scala 25:25]
  assign crossBar_io_mmioAxi_rd_bits_last = mmio_io_mmioAxi_rd_bits_last; // @[playground/src/sim/sim_core.scala 25:25]
  assign transAxi_io_raw_axi_awvalid = cpu_io_master_awvalid; // @[playground/src/sim/sim_core.scala 23:19]
  assign transAxi_io_raw_axi_awaddr = cpu_io_master_awaddr; // @[playground/src/sim/sim_core.scala 23:19]
  assign transAxi_io_raw_axi_awid = cpu_io_master_awid; // @[playground/src/sim/sim_core.scala 23:19]
  assign transAxi_io_raw_axi_awlen = cpu_io_master_awlen; // @[playground/src/sim/sim_core.scala 23:19]
  assign transAxi_io_raw_axi_awsize = cpu_io_master_awsize; // @[playground/src/sim/sim_core.scala 23:19]
  assign transAxi_io_raw_axi_awburst = cpu_io_master_awburst; // @[playground/src/sim/sim_core.scala 23:19]
  assign transAxi_io_raw_axi_wvalid = cpu_io_master_wvalid; // @[playground/src/sim/sim_core.scala 23:19]
  assign transAxi_io_raw_axi_wdata = cpu_io_master_wdata; // @[playground/src/sim/sim_core.scala 23:19]
  assign transAxi_io_raw_axi_wstrb = cpu_io_master_wstrb; // @[playground/src/sim/sim_core.scala 23:19]
  assign transAxi_io_raw_axi_wlast = cpu_io_master_wlast; // @[playground/src/sim/sim_core.scala 23:19]
  assign transAxi_io_raw_axi_bready = cpu_io_master_bready; // @[playground/src/sim/sim_core.scala 23:19]
  assign transAxi_io_raw_axi_arvalid = cpu_io_master_arvalid; // @[playground/src/sim/sim_core.scala 23:19]
  assign transAxi_io_raw_axi_araddr = cpu_io_master_araddr; // @[playground/src/sim/sim_core.scala 23:19]
  assign transAxi_io_raw_axi_arid = cpu_io_master_arid; // @[playground/src/sim/sim_core.scala 23:19]
  assign transAxi_io_raw_axi_arlen = cpu_io_master_arlen; // @[playground/src/sim/sim_core.scala 23:19]
  assign transAxi_io_raw_axi_arsize = cpu_io_master_arsize; // @[playground/src/sim/sim_core.scala 23:19]
  assign transAxi_io_raw_axi_arburst = cpu_io_master_arburst; // @[playground/src/sim/sim_core.scala 23:19]
  assign transAxi_io_raw_axi_rready = cpu_io_master_rready; // @[playground/src/sim/sim_core.scala 23:19]
  assign transAxi_io_bun_axi_wa_ready = crossBar_io_inAxi_wa_ready; // @[playground/src/sim/sim_core.scala 24:25]
  assign transAxi_io_bun_axi_wd_ready = crossBar_io_inAxi_wd_ready; // @[playground/src/sim/sim_core.scala 24:25]
  assign transAxi_io_bun_axi_wr_valid = crossBar_io_inAxi_wr_valid; // @[playground/src/sim/sim_core.scala 24:25]
  assign transAxi_io_bun_axi_wr_bits_id = crossBar_io_inAxi_wr_bits_id; // @[playground/src/sim/sim_core.scala 24:25]
  assign transAxi_io_bun_axi_wr_bits_resp = crossBar_io_inAxi_wr_bits_resp; // @[playground/src/sim/sim_core.scala 24:25]
  assign transAxi_io_bun_axi_ra_ready = crossBar_io_inAxi_ra_ready; // @[playground/src/sim/sim_core.scala 24:25]
  assign transAxi_io_bun_axi_rd_valid = crossBar_io_inAxi_rd_valid; // @[playground/src/sim/sim_core.scala 24:25]
  assign transAxi_io_bun_axi_rd_bits_id = crossBar_io_inAxi_rd_bits_id; // @[playground/src/sim/sim_core.scala 24:25]
  assign transAxi_io_bun_axi_rd_bits_data = crossBar_io_inAxi_rd_bits_data; // @[playground/src/sim/sim_core.scala 24:25]
  assign transAxi_io_bun_axi_rd_bits_resp = crossBar_io_inAxi_rd_bits_resp; // @[playground/src/sim/sim_core.scala 24:25]
  assign transAxi_io_bun_axi_rd_bits_last = crossBar_io_inAxi_rd_bits_last; // @[playground/src/sim/sim_core.scala 24:25]
endmodule
