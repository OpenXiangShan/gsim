module UpdateRegs (
    input  [2047:0]     regs_data,
    input clock
);


endmodule